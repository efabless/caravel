*SPICE netlist created from verilog structural netlist module mgmt_protect by vlog2Spice (qflow)
*This file may contain array delimiters, not for use in simulation.

** Start of included library ./pdk/sky130_ef_io.spice
* Power pads library (sky130 power pads + overlays) sky130_ef_io
* Includes corner and fill cell subcircuits

*----------------------------------------------------------
* sky130_ef_io__vccd_hvc_pad
* Power pad connects pad to VCCD with unconnected HV clamp
*----------------------------------------------------------

.SUBCKT sky130_ef_io__vccd_hvc_pad AMUXBUS_A AMUXBUS_B DRN_HVC SRC_BDY_HVC VCCD_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying power pad (connects P_PAD to VCCD)
Xsky130_fd_io__top_power_hvc_base_q0 AMUXBUS_A AMUXBUS_B DRN_HVC VDDIO VCCD VCCD_PAD SRC_BDY_HVC VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_power_hvc_wpadv2

.ENDS

*----------------------------------------------------------
* sky130_ef_io__vccd_lvc_pad
* Power pad connects pad to VCCD with unconnected LV clamp
*----------------------------------------------------------

.SUBCKT sky130_ef_io__vccd_lvc_pad AMUXBUS_A AMUXBUS_B DRN_LVC1 DRN_LVC2 SRC_BDY_LVC1 SRC_BDY_LVC2 BDY2_B2B VCCD_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying power pad (connects P_PAD to VCCD)
Xsky130_fd_io__top_power_lvc_base_q0 AMUXBUS_A AMUXBUS_B BDY2_B2B DRN_LVC1 DRN_LVC2 VDDIO VCCD VCCD_PAD SRC_BDY_LVC1 SRC_BDY_LVC2 VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_power_lvc_wpad

.ENDS

*----------------------------------------------------------
* sky130_ef_io__vdda_lvc_pad
* Power pad connects pad to VDDA with unconnected LV clamp
*----------------------------------------------------------

.SUBCKT sky130_ef_io__vdda_lvc_pad AMUXBUS_A AMUXBUS_B DRN_LVC1 DRN_LVC2 SRC_BDY_LVC1 SRC_BDY_LVC2 BDY2_B2B VDDA_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying power pad (connects P_PAD to VDDA)
Xsky130_fd_io__top_power_lvc_base_q0 AMUXBUS_A AMUXBUS_B BDY2_B2B DRN_LVC1 DRN_LVC2 VDDIO VDDA VDDA_PAD SRC_BDY_LVC1 SRC_BDY_LVC2 VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_power_lvc_wpad

.ENDS

*----------------------------------------------------------
* sky130_ef_io__vdda_lvc_pad
* Power pad connects pad to VDDA with unconnected HV clamp
*----------------------------------------------------------

.SUBCKT sky130_ef_io__vdda_hvc_pad AMUXBUS_A AMUXBUS_B DRN_HVC SRC_BDY_HVC VDDA_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying power pad (connects P_PAD to VDDA)
Xsky130_fd_io__top_power_hvc_base_q0 AMUXBUS_A AMUXBUS_B DRN_HVC VDDIO VDDA VDDA_PAD SRC_BDY_HVC VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_power_hvc_wpadv2

.ENDS

*----------------------------------------------------------
* sky130_ef_io__vddio_lvc_pad
* Power pad connects pad to VDDIO with unconnected LV clamp
*----------------------------------------------------------

.SUBCKT sky130_ef_io__vddio_lvc_pad AMUXBUS_A AMUXBUS_B DRN_LVC1 DRN_LVC2 SRC_BDY_LVC1 SRC_BDY_LVC2 BDY2_B2B VDDIO_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying power pad (connects P_PAD and VDDIO_Q to VDDIO)
Xsky130_fd_io__top_power_lvc_base_q0 AMUXBUS_A AMUXBUS_B BDY2_B2B DRN_LVC1 DRN_LVC2 VDDIO VDDIO VDDIO_PAD SRC_BDY_LVC1 SRC_BDY_LVC2 VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_power_lvc_wpad

.ENDS

*----------------------------------------------------------
* sky130_ef_io__vddio_hvc_pad
* Power pad connects pad to VDDIO with unconnected HV clamp
*----------------------------------------------------------

.SUBCKT sky130_ef_io__vddio_hvc_pad AMUXBUS_A AMUXBUS_B DRN_HVC SRC_BDY_HVC VDDIO_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying power pad (connects P_PAD and VDDIO_Q to VDDIO)
Xsky130_fd_io__top_power_hvc_base_q0 AMUXBUS_A AMUXBUS_B DRN_HVC VDDIO VDDIO VDDIO_PAD SRC_BDY_HVC VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_power_hvc_wpadv2

.ENDS

*----------------------------------------------------------
* sky130_ef_io__vssd_lvc_pad
* Ground pad connects pad to VSSD with unconnected LV clamp
*----------------------------------------------------------

.SUBCKT sky130_ef_io__vssd_lvc_pad AMUXBUS_A AMUXBUS_B DRN_LVC1 DRN_LVC2 SRC_BDY_LVC1 SRC_BDY_LVC2 BDY2_B2B VSSD_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying ground pad (connects G_PAD to VSSD)
Xsky130_fd_io__top_ground_lvc_base_q0 AMUXBUS_A AMUXBUS_B BDY2_B2B DRN_LVC1 DRN_LVC2 VSSD VSSD_PAD VDDIO SRC_BDY_LVC1 SRC_BDY_LVC2 VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_ground_lvc_wpad

.ENDS

*----------------------------------------------------------
* sky130_ef_io__vssd_hvc_pad
* Ground pad connects pad to VSSD with unconnected HV clamp
*----------------------------------------------------------

.SUBCKT sky130_ef_io__vssd_hvc_pad AMUXBUS_A AMUXBUS_B DRN_HVC SRC_BDY_HVC VSSD_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying ground pad (connects G_PAD to VSSD)
Xsky130_fd_io__top_ground_hvc_base_q0 AMUXBUS_A AMUXBUS_B DRN_HVC VSSD VSSD_PAD VDDIO SRC_BDY_HVC VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_ground_hvc_wpad

.ENDS

*----------------------------------------------------------
* sky130_ef_io__vssio_lvc_pad
* Ground pad connects pad to VSSIO with unconnected LV clamp
*----------------------------------------------------------

.SUBCKT sky130_ef_io__vssio_lvc_pad AMUXBUS_A AMUXBUS_B DRN_LVC1 DRN_LVC2 SRC_BDY_LVC1 SRC_BDY_LVC2 BDY2_B2B VSSIO_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying ground pad (connects G_PAD and VSSIO_Q to VSSIO)
Xsky130_fd_io__top_ground_lvc_base_q0 AMUXBUS_A AMUXBUS_B BDY2_B2B DRN_LVC1 DRN_LVC2 VSSIO VSSIO_PAD VDDIO SRC_BDY_LVC1 SRC_BDY_LVC2 VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_ground_lvc_wpad

.ENDS

*----------------------------------------------------------
* sky130_ef_io__vssio_hvc_pad
* Ground pad connects pad to VSSIO with unconnected HV clamp
*----------------------------------------------------------

.SUBCKT sky130_ef_io__vssio_hvc_pad AMUXBUS_A AMUXBUS_B DRN_HVC SRC_BDY_HVC VSSIO_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying ground pad (connects G_PAD and VSSIO_Q to VSSIO)
Xsky130_fd_io__top_ground_hvc_base_q0 AMUXBUS_A AMUXBUS_B DRN_HVC VSSIO VSSIO_PAD VDDIO SRC_BDY_HVC VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_ground_hvc_wpad

.ENDS

*----------------------------------------------------------
* sky130_ef_io__vssa_lvc_pad
* Ground pad connects pad to VSSA with unconnected LV clamp
*----------------------------------------------------------

.SUBCKT sky130_ef_io__vssa_lvc_pad AMUXBUS_A AMUXBUS_B DRN_LVC1 DRN_LVC2 SRC_BDY_LVC1 SRC_BDY_LVC2 BDY2_B2B VSSA_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying ground pad (connects G_PAD to VSSA)
Xsky130_fd_io__top_ground_lvc_base_q0 AMUXBUS_A AMUXBUS_B BDY2_B2B DRN_LVC1 DRN_LVC2 VSSA VSSA_PAD VDDIO SRC_BDY_LVC1 SRC_BDY_LVC2 VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_ground_lvc_wpad

.ENDS

*----------------------------------------------------------
* sky130_ef_io__vssa_lvc_pad
* Ground pad connects pad to VSSA with unconnected HV clamp
*----------------------------------------------------------

.SUBCKT sky130_ef_io__vssa_hvc_pad AMUXBUS_A AMUXBUS_B DRN_HVC SRC_BDY_HVC VSSA_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying ground pad (connects G_PAD to VSSA)
Xsky130_fd_io__top_ground_hvc_base_q0 AMUXBUS_A AMUXBUS_B DRN_HVC VSSA VSSA_PAD VDDIO SRC_BDY_HVC VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_ground_hvc_wpad
.ENDS

*----------------------------------------------------------
* sky130_ef_io__corner_pad
* Plain corner pad
*----------------------------------------------------------

.SUBCKT sky130_ef_io__corner_pad AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
* Corner pad has no active circuitry
.ENDS

*----------------------------------------------------------
* sky130_fd_io__com_bus_slice
* SkyWater padframe filler
*----------------------------------------------------------

.SUBCKT sky130_fd_io__com_bus_slice AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
* Bus filler has no active circuitry
.ENDS

*----------------------------------------------------------
* sky130_ef_io__com_bus_slice_1um
* 1um wide padframe filler
*----------------------------------------------------------

.SUBCKT sky130_ef_io__com_bus_slice_1um AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
* Bus filler has no active circuitry
.ENDS

*----------------------------------------------------------
* sky130_ef_io__com_bus_slice_5um
* 5um wide padframe filler
*----------------------------------------------------------

.SUBCKT sky130_ef_io__com_bus_slice_5um AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
* Bus filler has no active circuitry
.ENDS

*----------------------------------------------------------
* sky130_ef_io__com_bus_slice_10um
* 10um wide padframe filler
*----------------------------------------------------------

.SUBCKT sky130_ef_io__com_bus_slice_10um AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
* Bus filler has no active circuitry
.ENDS

*----------------------------------------------------------
* sky130_ef_io__com_bus_slice_20um
* 20um wide padframe filler
*----------------------------------------------------------

.SUBCKT sky130_ef_io__com_bus_slice_20um AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
* Bus filler has no active circuitry
.ENDS

*----------------------------------------------------------
* sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
* A 20um-wide padframe filler that connects VCCHIB and VCCD as well as
* VSWITCH and VDDIO
*----------------------------------------------------------

.SUBCKT sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um AMUXBUS_A AMUXBUS_B VSSA VDDA VDDIO_Q VDDIO VCCD VSSIO VSSD VSSIO_Q
* Bus filler has no active circuitry
.ENDS

*----------------------------------------------------------
* sky130_ef_io__disconnect_vdda_slice_5um
* A 5um-wide padframe filler that doesn't connect VDDA
* through it
*----------------------------------------------------------

.SUBCKT sky130_ef_io__disconnect_vdda_slice_5um AMUXBUS_A AMUXBUS_B VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
* Bus filler has no active circuitry
.ENDS

*----------------------------------------------------------
* sky130_ef_io__disconnect_vccd_slice_5um
* A 5um-wide padframe filler that doesn't connect VCCD
* through it
*----------------------------------------------------------

.SUBCKT sky130_ef_io__disconnect_vccd_slice_5um AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VSSIO VSSIO_Q
* Bus filler has no active circuitry
.ENDS

*----------------------------------------------------------
* sky130_ef_io__gpiov2_pad
* Wrapper around SkyWater gpiov2 pad
*----------------------------------------------------------

.SUBCKT sky130_ef_io__gpiov2_pad IN_H PAD_A_NOESD_H PAD_A_ESD_0_H PAD_A_ESD_1_H PAD DM[2] DM[1] DM[0] HLD_H_N IN INP_DIS IB_MODE_SEL ENABLE_H ENABLE_VDDA_H ENABLE_INP_H OE_N TIE_HI_ESD TIE_LO_ESD SLOW VTRIP_SEL HLD_OVR ANALOG_EN ANALOG_SEL ENABLE_VDDIO ENABLE_VSWITCH_H ANALOG_POL OUT AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate original version with metal4-only power bus
Xgpiov2_base_q0 AMUXBUS_A AMUXBUS_B ANALOG_EN ANALOG_POL ANALOG_SEL DM[2] DM[1] DM[0] ENABLE_H ENABLE_INP_H ENABLE_VDDA_H ENABLE_VDDIO ENABLE_VSWITCH_H HLD_H_N HLD_OVR IB_MODE_SEL IN IN_H INP_DIS OE_N OUT PAD PAD_A_ESD_0_H PAD_A_ESD_1_H PAD_A_NOESD_H SLOW TIE_HI_ESD TIE_LO_ESD VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH VTRIP_SEL sky130_fd_io__top_gpiov2

.ENDS

*----------------------------------------------------------
* sky130_ef_io__gpiov2_pad_wrapped
* Wrapper around sky130_ef_io__gpiov2_pad that forces
* the core-facing pins on tracks
*----------------------------------------------------------

.SUBCKT sky130_ef_io__gpiov2_pad_wrapped IN_H PAD_A_NOESD_H PAD_A_ESD_0_H PAD_A_ESD_1_H PAD DM[2] DM[1] DM[0] HLD_H_N IN INP_DIS IB_MODE_SEL ENABLE_H ENABLE_VDDA_H ENABLE_INP_H OE_N TIE_HI_ESD TIE_LO_ESD SLOW VTRIP_SEL HLD_OVR ANALOG_EN ANALOG_SEL ENABLE_VDDIO ENABLE_VSWITCH_H ANALOG_POL OUT AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

Xgpiov2_ef_q0 IN_H PAD_A_NOESD_H PAD_A_ESD_0_H PAD_A_ESD_1_H PAD DM[2] DM[1] DM[0] HLD_H_N IN INP_DIS IB_MODE_SEL ENABLE_H ENABLE_VDDA_H ENABLE_INP_H OE_N TIE_HI_ESD TIE_LO_ESD SLOW VTRIP_SEL HLD_OVR ANALOG_EN ANALOG_SEL ENABLE_VDDIO ENABLE_VSWITCH_H ANALOG_POL OUT AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q sky130_ef_io__gpiov2_pad

.ENDS

*--------------------------------------------------------------------------
* sky130_ef_io__vddio_hvc_clamped_pad
* sky130_ef_io__vddio_hvc_pad with HV clamp connections to VDDIO and VSSIO
*--------------------------------------------------------------------------

.SUBCKT sky130_ef_io__vddio_hvc_clamped_pad AMUXBUS_A AMUXBUS_B VDDIO_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying power pad (connects P_PAD and VDDIO_Q to VDDIO)
Xsky130_fd_io__top_power_hvc_base_q0 AMUXBUS_A AMUXBUS_B VDDIO VDDIO VDDIO VDDIO_PAD VSSIO VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_power_hvc_wpadv2

.ENDS

*--------------------------------------------------------------------------
* sky130_ef_io__vssio_hvc_clamped_pad
* sky130_ef_io__vssio_hvc_pad with HV clamp connections to VDDIO and VSSIO
*--------------------------------------------------------------------------

.SUBCKT sky130_ef_io__vssio_hvc_clamped_pad AMUXBUS_A AMUXBUS_B VSSIO_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying ground pad (connects G_PAD and VSSIO_Q to VSSIO)
Xsky130_fd_io__top_ground_hvc_base_q0 AMUXBUS_A AMUXBUS_B VDDIO VSSIO VSSIO_PAD VDDIO VSSIO VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_ground_hvc_wpad

.ENDS

*--------------------------------------------------------------------------
* sky130_ef_io__vdda_hvc_clamped_pad
* sky130_ef_io__vdda_hvc_pad with HV clamp connections to VDDA and VSSA
*--------------------------------------------------------------------------

.SUBCKT sky130_ef_io__vdda_hvc_clamped_pad AMUXBUS_A AMUXBUS_B VDDA_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying power pad (connects P_PAD to VDDA)
Xsky130_fd_io__top_power_hvc_base_q0 AMUXBUS_A AMUXBUS_B VDDA VDDIO VDDA VDDA_PAD VSSA VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_power_hvc_wpadv2

.ENDS

*--------------------------------------------------------------------------
* sky130_ef_io__vssa_hvc_clamped_pad
* sky130_ef_io__vssa_hvc_pad with HV clamp connections to VDDA and VSSA
*--------------------------------------------------------------------------

.SUBCKT sky130_ef_io__vssa_hvc_clamped_pad AMUXBUS_A AMUXBUS_B VSSA_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying ground pad (connects G_PAD to VSSA)
Xsky130_fd_io__top_ground_hvc_base_q0 AMUXBUS_A AMUXBUS_B VDDA VSSA VSSA_PAD VDDIO VSSA VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_ground_hvc_wpad

.ENDS

*--------------------------------------------------------------------------
* sky130_ef_io__vccd_lvc_clamped2_pad
* sky130_ef_io__vccd_lvc_pad with LV clamp connections to VCCD/VSSIO and
* VCCD/VSSD, and back-to-back diodes connecting VSSIO to VSSA
*--------------------------------------------------------------------------

.SUBCKT sky130_ef_io__vccd_lvc_clamped2_pad AMUXBUS_A AMUXBUS_B VCCD_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying power pad (connects P_PAD to VCCD)
Xsky130_fd_io__top_power_lvc_base_q0 AMUXBUS_A AMUXBUS_B VSSA VCCD VCCD VDDIO VCCD VCCD_PAD VSSIO VSSD VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_power_lvc_wpad

.ENDS

*--------------------------------------------------------------------------
* sky130_ef_io__vssd_lvc_clamped2_pad
* sky130_ef_io__vssd_lvc_pad with LV clamp connections to VCCD/VSSIO and
* VCCD/VSSD, and back-to-back diodes connecting VSSIO to VSSA
*--------------------------------------------------------------------------

.SUBCKT sky130_ef_io__vssd_lvc_clamped2_pad AMUXBUS_A AMUXBUS_B VSSD_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying ground pad (connects G_PAD to VSSD)
Xsky130_fd_io__top_ground_lvc_base_q0 AMUXBUS_A AMUXBUS_B VSSA VCCD VCCD VSSD VSSD_PAD VDDIO VSSIO VSSD VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_ground_lvc_wpad

.ENDS

*--------------------------------------------------------------------------
* sky130_ef_io__vccd_lvc_clamped3_pad
* sky130_ef_io__vccd_lvc_pad with pad and LV clamp positive connection to
* VCCD1, clamp negative connection to VSSD1, and and back-to-back diodes
* connecting VSSIO to VSSD1
*--------------------------------------------------------------------------

.SUBCKT sky130_ef_io__vccd_lvc_clamped3_pad AMUXBUS_A AMUXBUS_B VCCD_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q VCCD1 VSSD1

* Instantiate the underlying power pad (connects P_PAD to VCCD)
Xsky130_fd_io__top_power_lvc_base_q0 AMUXBUS_A AMUXBUS_B VSSD1 VCCD1 VCCD1 VDDIO VCCD1 VCCD_PAD VSSIO VSSD1 VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_power_lvc_wpad

.ENDS

*--------------------------------------------------------------------------
* sky130_ef_io__vssd_lvc_clamped3_pad
* sky130_ef_io__vssd_lvc_pad with pad and LV clamp negative connection to
* VSSD1, clamp positive connection to VCCD1, and back-to-back diodes
* connecting VSSIO to VSSD1
*--------------------------------------------------------------------------

.SUBCKT sky130_ef_io__vssd_lvc_clamped3_pad AMUXBUS_A AMUXBUS_B VSSD_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q VCCD1 VSSD1

* Instantiate the underlying ground pad (connects G_PAD to VSSD)
Xsky130_fd_io__top_ground_lvc_base_q0 AMUXBUS_A AMUXBUS_B VSSIO VCCD1 VCCD1 VSSD1 VSSD_PAD VDDIO VSSIO VSSD VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_ground_lvc_wpad

.ENDS

*--------------------------------------------------------------------------
* sky130_ef_io__vccd_lvc_clamped_pad
* sky130_ef_io__vccd_lvc_pad with LV clamp connections to VCCD and VSSD,
* and back-to-back diodes connecting VSSD to VSSIO
*--------------------------------------------------------------------------

.SUBCKT sky130_ef_io__vccd_lvc_clamped_pad AMUXBUS_A AMUXBUS_B VCCD_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying power pad (connects P_PAD to VCCD)
Xsky130_fd_io__top_power_lvc_base_q0 AMUXBUS_A AMUXBUS_B VSSIO VCCD VCCD VDDIO VCCD VCCD_PAD VSSD VSSD VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_power_lvc_wpad

.ENDS

*--------------------------------------------------------------------------
* sky130_ef_io__vssd_lvc_clamped_pad
* sky130_ef_io__vssd_lvc_pad with LV clamp connections to VCCD and VSSD,
* and back-to-back diodes connecting VSSD to VSSIO
*--------------------------------------------------------------------------

.SUBCKT sky130_ef_io__vssd_lvc_clamped_pad AMUXBUS_A AMUXBUS_B VSSD_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying ground pad (connects G_PAD to VSSD)
Xsky130_fd_io__top_ground_lvc_base_q0 AMUXBUS_A AMUXBUS_B VSSIO VCCD VCCD VSSD VSSD_PAD VDDIO VSSD VSSD VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_ground_lvc_wpad

.ENDS

*----------------------------------------------------------
* sky130_ef_io__top_power_hvc
* Power pad instantiates top_power_hvc_wpadv2 unchanged
* except for tripling the amount of metal at the core
* connection, for high-current supply applications.
*----------------------------------------------------------

.SUBCKT sky130_ef_io__top_power_hvc AMUXBUS_A AMUXBUS_B DRN_HVC P_CORE P_PAD SRC_BDY_HVC VCCD_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying power pad (connects P_PAD to VCCD)
Xsky130_fd_io__top_power_hvc_base_q0 AMUXBUS_A AMUXBUS_B DRN_HVC VDDIO P_CORE P_PAD SRC_BDY_HVC VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_power_hvc_wpadv2

.ENDS

*--------------------------------------------------------------------------
** End of included library ./pdk/sky130_ef_io.spice
** Start of included library ./pdk/sky130_ef_io.spice
* Power pads library (sky130 power pads + overlays) sky130_ef_io
* Includes corner and fill cell subcircuits

*----------------------------------------------------------
* sky130_ef_io__vccd_hvc_pad
* Power pad connects pad to VCCD with unconnected HV clamp
*----------------------------------------------------------

.SUBCKT sky130_ef_io__vccd_hvc_pad AMUXBUS_A AMUXBUS_B DRN_HVC SRC_BDY_HVC VCCD_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying power pad (connects P_PAD to VCCD)
Xsky130_fd_io__top_power_hvc_base_q0 AMUXBUS_A AMUXBUS_B DRN_HVC VDDIO VCCD VCCD_PAD SRC_BDY_HVC VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_power_hvc_wpadv2

.ENDS

*----------------------------------------------------------
* sky130_ef_io__vccd_lvc_pad
* Power pad connects pad to VCCD with unconnected LV clamp
*----------------------------------------------------------

.SUBCKT sky130_ef_io__vccd_lvc_pad AMUXBUS_A AMUXBUS_B DRN_LVC1 DRN_LVC2 SRC_BDY_LVC1 SRC_BDY_LVC2 BDY2_B2B VCCD_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying power pad (connects P_PAD to VCCD)
Xsky130_fd_io__top_power_lvc_base_q0 AMUXBUS_A AMUXBUS_B BDY2_B2B DRN_LVC1 DRN_LVC2 VDDIO VCCD VCCD_PAD SRC_BDY_LVC1 SRC_BDY_LVC2 VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_power_lvc_wpad

.ENDS

*----------------------------------------------------------
* sky130_ef_io__vdda_lvc_pad
* Power pad connects pad to VDDA with unconnected LV clamp
*----------------------------------------------------------

.SUBCKT sky130_ef_io__vdda_lvc_pad AMUXBUS_A AMUXBUS_B DRN_LVC1 DRN_LVC2 SRC_BDY_LVC1 SRC_BDY_LVC2 BDY2_B2B VDDA_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying power pad (connects P_PAD to VDDA)
Xsky130_fd_io__top_power_lvc_base_q0 AMUXBUS_A AMUXBUS_B BDY2_B2B DRN_LVC1 DRN_LVC2 VDDIO VDDA VDDA_PAD SRC_BDY_LVC1 SRC_BDY_LVC2 VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_power_lvc_wpad

.ENDS

*----------------------------------------------------------
* sky130_ef_io__vdda_lvc_pad
* Power pad connects pad to VDDA with unconnected HV clamp
*----------------------------------------------------------

.SUBCKT sky130_ef_io__vdda_hvc_pad AMUXBUS_A AMUXBUS_B DRN_HVC SRC_BDY_HVC VDDA_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying power pad (connects P_PAD to VDDA)
Xsky130_fd_io__top_power_hvc_base_q0 AMUXBUS_A AMUXBUS_B DRN_HVC VDDIO VDDA VDDA_PAD SRC_BDY_HVC VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_power_hvc_wpadv2

.ENDS

*----------------------------------------------------------
* sky130_ef_io__vddio_lvc_pad
* Power pad connects pad to VDDIO with unconnected LV clamp
*----------------------------------------------------------

.SUBCKT sky130_ef_io__vddio_lvc_pad AMUXBUS_A AMUXBUS_B DRN_LVC1 DRN_LVC2 SRC_BDY_LVC1 SRC_BDY_LVC2 BDY2_B2B VDDIO_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying power pad (connects P_PAD and VDDIO_Q to VDDIO)
Xsky130_fd_io__top_power_lvc_base_q0 AMUXBUS_A AMUXBUS_B BDY2_B2B DRN_LVC1 DRN_LVC2 VDDIO VDDIO VDDIO_PAD SRC_BDY_LVC1 SRC_BDY_LVC2 VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_power_lvc_wpad

.ENDS

*----------------------------------------------------------
* sky130_ef_io__vddio_hvc_pad
* Power pad connects pad to VDDIO with unconnected HV clamp
*----------------------------------------------------------

.SUBCKT sky130_ef_io__vddio_hvc_pad AMUXBUS_A AMUXBUS_B DRN_HVC SRC_BDY_HVC VDDIO_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying power pad (connects P_PAD and VDDIO_Q to VDDIO)
Xsky130_fd_io__top_power_hvc_base_q0 AMUXBUS_A AMUXBUS_B DRN_HVC VDDIO VDDIO VDDIO_PAD SRC_BDY_HVC VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_power_hvc_wpadv2

.ENDS

*----------------------------------------------------------
* sky130_ef_io__vssd_lvc_pad
* Ground pad connects pad to VSSD with unconnected LV clamp
*----------------------------------------------------------

.SUBCKT sky130_ef_io__vssd_lvc_pad AMUXBUS_A AMUXBUS_B DRN_LVC1 DRN_LVC2 SRC_BDY_LVC1 SRC_BDY_LVC2 BDY2_B2B VSSD_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying ground pad (connects G_PAD to VSSD)
Xsky130_fd_io__top_ground_lvc_base_q0 AMUXBUS_A AMUXBUS_B BDY2_B2B DRN_LVC1 DRN_LVC2 VSSD VSSD_PAD VDDIO SRC_BDY_LVC1 SRC_BDY_LVC2 VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_ground_lvc_wpad

.ENDS

*----------------------------------------------------------
* sky130_ef_io__vssd_hvc_pad
* Ground pad connects pad to VSSD with unconnected HV clamp
*----------------------------------------------------------

.SUBCKT sky130_ef_io__vssd_hvc_pad AMUXBUS_A AMUXBUS_B DRN_HVC SRC_BDY_HVC VSSD_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying ground pad (connects G_PAD to VSSD)
Xsky130_fd_io__top_ground_hvc_base_q0 AMUXBUS_A AMUXBUS_B DRN_HVC VSSD VSSD_PAD VDDIO SRC_BDY_HVC VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_ground_hvc_wpad

.ENDS

*----------------------------------------------------------
* sky130_ef_io__vssio_lvc_pad
* Ground pad connects pad to VSSIO with unconnected LV clamp
*----------------------------------------------------------

.SUBCKT sky130_ef_io__vssio_lvc_pad AMUXBUS_A AMUXBUS_B DRN_LVC1 DRN_LVC2 SRC_BDY_LVC1 SRC_BDY_LVC2 BDY2_B2B VSSIO_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying ground pad (connects G_PAD and VSSIO_Q to VSSIO)
Xsky130_fd_io__top_ground_lvc_base_q0 AMUXBUS_A AMUXBUS_B BDY2_B2B DRN_LVC1 DRN_LVC2 VSSIO VSSIO_PAD VDDIO SRC_BDY_LVC1 SRC_BDY_LVC2 VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_ground_lvc_wpad

.ENDS

*----------------------------------------------------------
* sky130_ef_io__vssio_hvc_pad
* Ground pad connects pad to VSSIO with unconnected HV clamp
*----------------------------------------------------------

.SUBCKT sky130_ef_io__vssio_hvc_pad AMUXBUS_A AMUXBUS_B DRN_HVC SRC_BDY_HVC VSSIO_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying ground pad (connects G_PAD and VSSIO_Q to VSSIO)
Xsky130_fd_io__top_ground_hvc_base_q0 AMUXBUS_A AMUXBUS_B DRN_HVC VSSIO VSSIO_PAD VDDIO SRC_BDY_HVC VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_ground_hvc_wpad

.ENDS

*----------------------------------------------------------
* sky130_ef_io__vssa_lvc_pad
* Ground pad connects pad to VSSA with unconnected LV clamp
*----------------------------------------------------------

.SUBCKT sky130_ef_io__vssa_lvc_pad AMUXBUS_A AMUXBUS_B DRN_LVC1 DRN_LVC2 SRC_BDY_LVC1 SRC_BDY_LVC2 BDY2_B2B VSSA_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying ground pad (connects G_PAD to VSSA)
Xsky130_fd_io__top_ground_lvc_base_q0 AMUXBUS_A AMUXBUS_B BDY2_B2B DRN_LVC1 DRN_LVC2 VSSA VSSA_PAD VDDIO SRC_BDY_LVC1 SRC_BDY_LVC2 VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_ground_lvc_wpad

.ENDS

*----------------------------------------------------------
* sky130_ef_io__vssa_lvc_pad
* Ground pad connects pad to VSSA with unconnected HV clamp
*----------------------------------------------------------

.SUBCKT sky130_ef_io__vssa_hvc_pad AMUXBUS_A AMUXBUS_B DRN_HVC SRC_BDY_HVC VSSA_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying ground pad (connects G_PAD to VSSA)
Xsky130_fd_io__top_ground_hvc_base_q0 AMUXBUS_A AMUXBUS_B DRN_HVC VSSA VSSA_PAD VDDIO SRC_BDY_HVC VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_ground_hvc_wpad
.ENDS

*----------------------------------------------------------
* sky130_ef_io__corner_pad
* Plain corner pad
*----------------------------------------------------------

.SUBCKT sky130_ef_io__corner_pad AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
* Corner pad has no active circuitry
.ENDS

*----------------------------------------------------------
* sky130_fd_io__com_bus_slice
* SkyWater padframe filler
*----------------------------------------------------------

.SUBCKT sky130_fd_io__com_bus_slice AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
* Bus filler has no active circuitry
.ENDS

*----------------------------------------------------------
* sky130_ef_io__com_bus_slice_1um
* 1um wide padframe filler
*----------------------------------------------------------

.SUBCKT sky130_ef_io__com_bus_slice_1um AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
* Bus filler has no active circuitry
.ENDS

*----------------------------------------------------------
* sky130_ef_io__com_bus_slice_5um
* 5um wide padframe filler
*----------------------------------------------------------

.SUBCKT sky130_ef_io__com_bus_slice_5um AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
* Bus filler has no active circuitry
.ENDS

*----------------------------------------------------------
* sky130_ef_io__com_bus_slice_10um
* 10um wide padframe filler
*----------------------------------------------------------

.SUBCKT sky130_ef_io__com_bus_slice_10um AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
* Bus filler has no active circuitry
.ENDS

*----------------------------------------------------------
* sky130_ef_io__com_bus_slice_20um
* 20um wide padframe filler
*----------------------------------------------------------

.SUBCKT sky130_ef_io__com_bus_slice_20um AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
* Bus filler has no active circuitry
.ENDS

*----------------------------------------------------------
* sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
* A 20um-wide padframe filler that connects VCCHIB and VCCD as well as
* VSWITCH and VDDIO
*----------------------------------------------------------

.SUBCKT sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um AMUXBUS_A AMUXBUS_B VSSA VDDA VDDIO_Q VDDIO VCCD VSSIO VSSD VSSIO_Q
* Bus filler has no active circuitry
.ENDS

*----------------------------------------------------------
* sky130_ef_io__disconnect_vdda_slice_5um
* A 5um-wide padframe filler that doesn't connect VDDA
* through it
*----------------------------------------------------------

.SUBCKT sky130_ef_io__disconnect_vdda_slice_5um AMUXBUS_A AMUXBUS_B VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
* Bus filler has no active circuitry
.ENDS

*----------------------------------------------------------
* sky130_ef_io__disconnect_vccd_slice_5um
* A 5um-wide padframe filler that doesn't connect VCCD
* through it
*----------------------------------------------------------

.SUBCKT sky130_ef_io__disconnect_vccd_slice_5um AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VSSIO VSSIO_Q
* Bus filler has no active circuitry
.ENDS

*----------------------------------------------------------
* sky130_ef_io__gpiov2_pad
* Wrapper around SkyWater gpiov2 pad
*----------------------------------------------------------

.SUBCKT sky130_ef_io__gpiov2_pad IN_H PAD_A_NOESD_H PAD_A_ESD_0_H PAD_A_ESD_1_H PAD DM[2] DM[1] DM[0] HLD_H_N IN INP_DIS IB_MODE_SEL ENABLE_H ENABLE_VDDA_H ENABLE_INP_H OE_N TIE_HI_ESD TIE_LO_ESD SLOW VTRIP_SEL HLD_OVR ANALOG_EN ANALOG_SEL ENABLE_VDDIO ENABLE_VSWITCH_H ANALOG_POL OUT AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate original version with metal4-only power bus
Xgpiov2_base_q0 AMUXBUS_A AMUXBUS_B ANALOG_EN ANALOG_POL ANALOG_SEL DM[2] DM[1] DM[0] ENABLE_H ENABLE_INP_H ENABLE_VDDA_H ENABLE_VDDIO ENABLE_VSWITCH_H HLD_H_N HLD_OVR IB_MODE_SEL IN IN_H INP_DIS OE_N OUT PAD PAD_A_ESD_0_H PAD_A_ESD_1_H PAD_A_NOESD_H SLOW TIE_HI_ESD TIE_LO_ESD VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH VTRIP_SEL sky130_fd_io__top_gpiov2

.ENDS

*----------------------------------------------------------
* sky130_ef_io__gpiov2_pad_wrapped
* Wrapper around sky130_ef_io__gpiov2_pad that forces
* the core-facing pins on tracks
*----------------------------------------------------------

.SUBCKT sky130_ef_io__gpiov2_pad_wrapped IN_H PAD_A_NOESD_H PAD_A_ESD_0_H PAD_A_ESD_1_H PAD DM[2] DM[1] DM[0] HLD_H_N IN INP_DIS IB_MODE_SEL ENABLE_H ENABLE_VDDA_H ENABLE_INP_H OE_N TIE_HI_ESD TIE_LO_ESD SLOW VTRIP_SEL HLD_OVR ANALOG_EN ANALOG_SEL ENABLE_VDDIO ENABLE_VSWITCH_H ANALOG_POL OUT AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

Xgpiov2_ef_q0 IN_H PAD_A_NOESD_H PAD_A_ESD_0_H PAD_A_ESD_1_H PAD DM[2] DM[1] DM[0] HLD_H_N IN INP_DIS IB_MODE_SEL ENABLE_H ENABLE_VDDA_H ENABLE_INP_H OE_N TIE_HI_ESD TIE_LO_ESD SLOW VTRIP_SEL HLD_OVR ANALOG_EN ANALOG_SEL ENABLE_VDDIO ENABLE_VSWITCH_H ANALOG_POL OUT AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q sky130_ef_io__gpiov2_pad

.ENDS

*--------------------------------------------------------------------------
* sky130_ef_io__vddio_hvc_clamped_pad
* sky130_ef_io__vddio_hvc_pad with HV clamp connections to VDDIO and VSSIO
*--------------------------------------------------------------------------

.SUBCKT sky130_ef_io__vddio_hvc_clamped_pad AMUXBUS_A AMUXBUS_B VDDIO_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying power pad (connects P_PAD and VDDIO_Q to VDDIO)
Xsky130_fd_io__top_power_hvc_base_q0 AMUXBUS_A AMUXBUS_B VDDIO VDDIO VDDIO VDDIO_PAD VSSIO VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_power_hvc_wpadv2

.ENDS

*--------------------------------------------------------------------------
* sky130_ef_io__vssio_hvc_clamped_pad
* sky130_ef_io__vssio_hvc_pad with HV clamp connections to VDDIO and VSSIO
*--------------------------------------------------------------------------

.SUBCKT sky130_ef_io__vssio_hvc_clamped_pad AMUXBUS_A AMUXBUS_B VSSIO_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying ground pad (connects G_PAD and VSSIO_Q to VSSIO)
Xsky130_fd_io__top_ground_hvc_base_q0 AMUXBUS_A AMUXBUS_B VDDIO VSSIO VSSIO_PAD VDDIO VSSIO VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_ground_hvc_wpad

.ENDS

*--------------------------------------------------------------------------
* sky130_ef_io__vdda_hvc_clamped_pad
* sky130_ef_io__vdda_hvc_pad with HV clamp connections to VDDA and VSSA
*--------------------------------------------------------------------------

.SUBCKT sky130_ef_io__vdda_hvc_clamped_pad AMUXBUS_A AMUXBUS_B VDDA_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying power pad (connects P_PAD to VDDA)
Xsky130_fd_io__top_power_hvc_base_q0 AMUXBUS_A AMUXBUS_B VDDA VDDIO VDDA VDDA_PAD VSSA VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_power_hvc_wpadv2

.ENDS

*--------------------------------------------------------------------------
* sky130_ef_io__vssa_hvc_clamped_pad
* sky130_ef_io__vssa_hvc_pad with HV clamp connections to VDDA and VSSA
*--------------------------------------------------------------------------

.SUBCKT sky130_ef_io__vssa_hvc_clamped_pad AMUXBUS_A AMUXBUS_B VSSA_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying ground pad (connects G_PAD to VSSA)
Xsky130_fd_io__top_ground_hvc_base_q0 AMUXBUS_A AMUXBUS_B VDDA VSSA VSSA_PAD VDDIO VSSA VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_ground_hvc_wpad

.ENDS

*--------------------------------------------------------------------------
* sky130_ef_io__vccd_lvc_clamped2_pad
* sky130_ef_io__vccd_lvc_pad with LV clamp connections to VCCD/VSSIO and
* VCCD/VSSD, and back-to-back diodes connecting VSSIO to VSSA
*--------------------------------------------------------------------------

.SUBCKT sky130_ef_io__vccd_lvc_clamped2_pad AMUXBUS_A AMUXBUS_B VCCD_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying power pad (connects P_PAD to VCCD)
Xsky130_fd_io__top_power_lvc_base_q0 AMUXBUS_A AMUXBUS_B VSSA VCCD VCCD VDDIO VCCD VCCD_PAD VSSIO VSSD VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_power_lvc_wpad

.ENDS

*--------------------------------------------------------------------------
* sky130_ef_io__vssd_lvc_clamped2_pad
* sky130_ef_io__vssd_lvc_pad with LV clamp connections to VCCD/VSSIO and
* VCCD/VSSD, and back-to-back diodes connecting VSSIO to VSSA
*--------------------------------------------------------------------------

.SUBCKT sky130_ef_io__vssd_lvc_clamped2_pad AMUXBUS_A AMUXBUS_B VSSD_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying ground pad (connects G_PAD to VSSD)
Xsky130_fd_io__top_ground_lvc_base_q0 AMUXBUS_A AMUXBUS_B VSSA VCCD VCCD VSSD VSSD_PAD VDDIO VSSIO VSSD VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_ground_lvc_wpad

.ENDS

*--------------------------------------------------------------------------
* sky130_ef_io__vccd_lvc_clamped3_pad
* sky130_ef_io__vccd_lvc_pad with pad and LV clamp positive connection to
* VCCD1, clamp negative connection to VSSD1, and and back-to-back diodes
* connecting VSSIO to VSSD1
*--------------------------------------------------------------------------

.SUBCKT sky130_ef_io__vccd_lvc_clamped3_pad AMUXBUS_A AMUXBUS_B VCCD_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q VCCD1 VSSD1

* Instantiate the underlying power pad (connects P_PAD to VCCD)
Xsky130_fd_io__top_power_lvc_base_q0 AMUXBUS_A AMUXBUS_B VSSD1 VCCD1 VCCD1 VDDIO VCCD1 VCCD_PAD VSSIO VSSD1 VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_power_lvc_wpad

.ENDS

*--------------------------------------------------------------------------
* sky130_ef_io__vssd_lvc_clamped3_pad
* sky130_ef_io__vssd_lvc_pad with pad and LV clamp negative connection to
* VSSD1, clamp positive connection to VCCD1, and back-to-back diodes
* connecting VSSIO to VSSD1
*--------------------------------------------------------------------------

.SUBCKT sky130_ef_io__vssd_lvc_clamped3_pad AMUXBUS_A AMUXBUS_B VSSD_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q VCCD1 VSSD1

* Instantiate the underlying ground pad (connects G_PAD to VSSD)
Xsky130_fd_io__top_ground_lvc_base_q0 AMUXBUS_A AMUXBUS_B VSSIO VCCD1 VCCD1 VSSD1 VSSD_PAD VDDIO VSSIO VSSD VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_ground_lvc_wpad

.ENDS

*--------------------------------------------------------------------------
* sky130_ef_io__vccd_lvc_clamped_pad
* sky130_ef_io__vccd_lvc_pad with LV clamp connections to VCCD and VSSD,
* and back-to-back diodes connecting VSSD to VSSIO
*--------------------------------------------------------------------------

.SUBCKT sky130_ef_io__vccd_lvc_clamped_pad AMUXBUS_A AMUXBUS_B VCCD_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying power pad (connects P_PAD to VCCD)
Xsky130_fd_io__top_power_lvc_base_q0 AMUXBUS_A AMUXBUS_B VSSIO VCCD VCCD VDDIO VCCD VCCD_PAD VSSD VSSD VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_power_lvc_wpad

.ENDS

*--------------------------------------------------------------------------
* sky130_ef_io__vssd_lvc_clamped_pad
* sky130_ef_io__vssd_lvc_pad with LV clamp connections to VCCD and VSSD,
* and back-to-back diodes connecting VSSD to VSSIO
*--------------------------------------------------------------------------

.SUBCKT sky130_ef_io__vssd_lvc_clamped_pad AMUXBUS_A AMUXBUS_B VSSD_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying ground pad (connects G_PAD to VSSD)
Xsky130_fd_io__top_ground_lvc_base_q0 AMUXBUS_A AMUXBUS_B VSSIO VCCD VCCD VSSD VSSD_PAD VDDIO VSSD VSSD VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_ground_lvc_wpad

.ENDS

*----------------------------------------------------------
* sky130_ef_io__top_power_hvc
* Power pad instantiates top_power_hvc_wpadv2 unchanged
* except for tripling the amount of metal at the core
* connection, for high-current supply applications.
*----------------------------------------------------------

.SUBCKT sky130_ef_io__top_power_hvc AMUXBUS_A AMUXBUS_B DRN_HVC P_CORE P_PAD SRC_BDY_HVC VCCD_PAD VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q

* Instantiate the underlying power pad (connects P_PAD to VCCD)
Xsky130_fd_io__top_power_hvc_base_q0 AMUXBUS_A AMUXBUS_B DRN_HVC VDDIO P_CORE P_PAD SRC_BDY_HVC VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH sky130_fd_io__top_power_hvc_wpadv2

.ENDS

*--------------------------------------------------------------------------
** End of included library ./pdk/sky130_ef_io.spice
** Start of included library ./pdk/sky130_fd_sc_hvl.spice
* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
X0 VPWR A2 a_469_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 X a_83_283# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X2 X a_83_283# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 a_631_107# A2 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 VGND B1 a_83_283# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X5 a_83_283# B1 a_469_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X6 a_83_283# A1 a_631_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X7 a_469_443# A1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
X0 Y B1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X1 VGND A2 a_271_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 a_56_443# A2 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X3 a_271_107# A1 Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 a_56_443# B1 Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X5 VPWR A1 a_56_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 X a_83_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X1 a_822_107# A2 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 a_316_443# B2 a_83_81# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X3 X a_83_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X4 a_316_443# A1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X5 VGND B2 a_519_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X6 a_519_107# B1 a_83_81# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X7 a_83_81# A1 a_822_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X8 a_83_81# B1 a_316_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X9 VPWR A2 a_316_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
X0 VGND B2 a_204_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X1 a_33_443# B2 Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X2 a_502_107# A2 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 a_204_107# B1 Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 Y B1 a_33_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X5 Y A1 a_502_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X6 VPWR A2 a_33_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X7 a_33_443# A1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__and2_1 A B VGND VNB VPB VPWR X
X0 VGND a_30_107# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X1 VPWR a_30_107# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X2 a_30_107# A a_183_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X3 a_183_107# B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X4 VPWR A a_30_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X5 a_30_107# B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__and3_1 A B C VGND VNB VPB VPWR X
X0 VGND a_30_517# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X1 a_201_173# B a_343_173# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X2 a_30_517# C VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X3 VPWR a_30_517# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X4 a_30_517# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X5 VPWR B a_30_517# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X6 a_30_517# A a_201_173# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X7 a_343_173# C VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__buf_1 A VGND VNB VPB VPWR X
X0 VPWR A a_84_81# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X1 X a_84_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 VGND A a_84_81# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X3 X a_84_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__buf_2 A VGND VNB VPB VPWR X
X0 VPWR A a_129_279# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X1 VPWR a_129_279# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X2 X a_129_279# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 VGND A a_129_279# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X4 X a_129_279# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X5 VGND a_129_279# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__buf_4 A VGND VNB VPB VPWR X
X0 X a_149_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X1 X a_149_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 X a_149_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X3 X a_149_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X4 VGND a_149_81# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X5 VGND A a_149_81# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X6 VPWR a_149_81# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X7 VPWR A a_149_81# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X8 VGND a_149_81# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X9 VPWR a_149_81# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__buf_8 A VGND VNB VPB VPWR X
X0 a_45_443# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X3 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X5 VGND A a_45_443# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X6 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X7 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X8 a_45_443# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X9 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X10 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X11 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X12 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X13 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X14 a_45_443# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X15 VPWR A a_45_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X16 a_45_443# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X17 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X18 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X19 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X20 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X21 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__buf_16 A VGND VNB VPB VPWR X
X0 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X2 a_183_141# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X5 VPWR A a_183_141# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X6 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X7 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X8 a_183_141# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X9 VPWR A a_183_141# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X10 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X11 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X12 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X13 VPWR A a_183_141# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X14 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X15 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X16 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X17 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X18 a_183_141# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X19 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X20 a_183_141# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X21 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X22 a_183_141# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X23 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X24 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X25 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X26 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X27 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X28 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X29 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X30 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X31 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X32 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X33 VGND A a_183_141# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X34 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X35 a_183_141# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X36 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X37 VGND A a_183_141# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X38 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X39 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X40 VGND A a_183_141# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X41 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X42 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X43 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__buf_32 A VGND VNB VPB VPWR X
X0 a_183_141# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X2 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X3 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X5 a_183_141# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X6 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X7 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X8 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X9 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X10 VPWR A a_183_141# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X11 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X12 VPWR A a_183_141# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X13 a_183_141# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X14 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X15 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X16 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X17 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X18 VPWR A a_183_141# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X19 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X20 VGND A a_183_141# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X21 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X22 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X23 VPWR A a_183_141# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X24 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X25 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X26 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X27 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X28 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X29 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X30 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X31 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X32 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X33 a_183_141# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X34 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X35 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X36 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X37 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X38 a_183_141# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X39 a_183_141# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X40 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X41 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X42 VPWR A a_183_141# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X43 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X44 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X45 a_183_141# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X46 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X47 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X48 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X49 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X50 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X51 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X52 a_183_141# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X53 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X54 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X55 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X56 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X57 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X58 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X59 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X60 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X61 VGND A a_183_141# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X62 VGND A a_183_141# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X63 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X64 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X65 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X66 a_183_141# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X67 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X68 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X69 VGND A a_183_141# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X70 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X71 VGND A a_183_141# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X72 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X73 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X74 a_183_141# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X75 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X76 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X77 X a_183_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X78 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X79 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X80 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X81 X a_183_141# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X82 VPWR a_183_141# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X83 VGND a_183_141# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__conb_1 VGND VNB VPB VPWR HI LO
R0 HI VPWR sky130_fd_pr__res_generic_po w=510000u l=45000u
R1 VGND LO sky130_fd_pr__res_generic_po w=510000u l=45000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__decap_4 VGND VNB VPB VPWR
X0 VGND VPWR VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=1e+06u
X1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=1e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__decap_8 VGND VNB VPB VPWR
X0 VGND VPWR VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=1e+06u
X1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=1e+06u
X2 VPWR VGND VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=1e+06u
X3 VGND VPWR VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=1e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__dfrbp_1 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
X0 a_1176_466# a_350_107# a_1900_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X1 a_37_107# CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X2 VGND a_2937_443# Q VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 a_2122_348# a_1900_107# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X4 VPWR RESET_B a_978_608# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X5 VGND a_37_107# a_350_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X6 a_978_608# a_350_107# a_1215_173# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X7 VPWR a_2937_443# Q VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X8 a_2412_107# a_1900_107# a_2122_348# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X9 a_978_608# a_37_107# a_1134_608# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X10 VPWR a_37_107# a_350_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X11 a_2114_107# a_2122_348# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X12 a_2937_443# a_1900_107# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X13 a_1900_107# a_350_107# a_2079_462# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X14 VPWR a_1900_107# Q_N VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X15 a_2079_462# a_2122_348# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X16 a_509_608# a_37_107# a_978_608# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X17 VGND RESET_B a_2412_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X18 VGND a_1900_107# Q_N VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X19 a_1357_173# RESET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X20 VPWR a_978_608# a_1176_466# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X21 a_1215_173# a_1176_466# a_1357_173# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X22 a_509_608# RESET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X23 VGND a_978_608# a_1176_466# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X24 a_2937_443# a_1900_107# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X25 a_509_608# a_350_107# a_978_608# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X26 VGND RESET_B a_728_173# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X27 a_37_107# CLK VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X28 a_728_173# D a_509_608# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X29 a_1900_107# a_37_107# a_2114_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X30 a_1134_608# a_1176_466# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X31 a_1176_466# a_37_107# a_1900_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X32 VPWR RESET_B a_2122_348# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X33 VPWR D a_509_608# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
X0 a_1233_173# RESET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X1 VGND RESET_B a_2387_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X2 VPWR a_921_632# a_1119_506# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X3 a_1091_173# a_1119_506# a_1233_173# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X4 a_30_107# CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X5 a_2089_107# a_2096_417# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X6 VPWR a_30_107# a_339_537# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X7 VGND RESET_B a_637_173# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X8 VPWR RESET_B a_921_632# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X9 VGND a_30_107# a_339_537# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X10 a_452_632# RESET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X11 a_2054_543# a_2096_417# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X12 a_921_632# a_339_537# a_1091_173# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X13 VPWR a_2649_207# Q VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X14 a_1875_543# a_339_537# a_2054_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X15 a_1119_506# a_30_107# a_1875_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X16 a_2387_107# a_1875_543# a_2096_417# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X17 a_2096_417# a_1875_543# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X18 a_1077_632# a_1119_506# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X19 a_30_107# CLK VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X20 a_1119_506# a_339_537# a_1875_543# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X21 VPWR D a_452_632# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X22 a_921_632# a_30_107# a_1077_632# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X23 VPWR RESET_B a_2096_417# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X24 a_637_173# D a_452_632# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X25 a_2649_207# a_1875_543# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X26 VGND a_921_632# a_1119_506# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X27 a_2649_207# a_1875_543# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X28 a_452_632# a_339_537# a_921_632# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X29 a_1875_543# a_30_107# a_2089_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X30 VGND a_2649_207# Q VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X31 a_452_632# a_30_107# a_921_632# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__dfsbp_1 CLK D SET_B VGND VNB VPB VPWR Q Q_N
X0 a_605_109# a_339_112# a_761_109# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X1 VPWR a_761_109# a_1732_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X2 a_1755_153# a_30_112# a_1874_543# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X3 a_917_109# a_959_83# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X4 VGND a_761_109# a_1642_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X5 a_1325_107# SET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X6 a_1874_543# a_339_112# a_1642_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X7 a_30_112# CLK VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X8 a_2427_107# SET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X9 VPWR a_3129_479# Q VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X10 a_3129_479# a_1874_543# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X11 VPWR a_30_112# a_339_112# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X12 VPWR a_761_109# a_959_83# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X13 VPWR a_1874_543# Q_N VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X14 a_2156_417# a_1874_543# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X15 a_2053_543# a_2156_417# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X16 VGND a_30_112# a_339_112# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X17 VGND a_3129_479# Q VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X18 VGND D a_605_109# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X19 a_1874_543# a_339_112# a_2053_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X20 a_976_543# a_959_83# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X21 a_1732_543# a_30_112# a_1874_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X22 a_761_109# a_339_112# a_917_109# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X23 a_959_83# SET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X24 VPWR SET_B a_1874_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X25 a_959_83# a_761_109# a_1325_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X26 a_2156_417# a_1874_543# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X27 a_1755_153# a_2156_417# a_2427_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X28 VPWR D a_605_109# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X29 VGND a_1874_543# Q_N VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X30 a_761_109# a_30_112# a_976_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X31 a_605_109# a_30_112# a_761_109# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X32 a_3129_479# a_1874_543# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X33 a_30_112# CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
X0 VPWR a_30_131# a_340_593# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X1 a_2553_203# a_1787_137# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X2 VPWR a_2553_203# Q VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X3 VGND a_798_107# a_1645_137# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 a_958_107# a_1000_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X5 a_1989_203# a_2031_177# a_2131_203# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X6 a_1268_251# SET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X7 a_982_529# a_1000_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X8 VPWR a_798_107# a_1000_81# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X9 a_1653_515# a_30_131# a_1787_137# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X10 VGND a_1787_137# a_2031_177# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X11 a_1787_137# a_340_593# a_1989_515# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X12 a_642_107# a_340_593# a_798_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X13 a_2553_203# a_1787_137# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X14 a_798_107# a_30_131# a_982_529# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X15 VPWR SET_B a_1787_137# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X16 a_642_107# a_30_131# a_798_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X17 a_1645_137# a_340_593# a_1787_137# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X18 VGND a_2553_203# Q VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X19 a_2031_177# a_1787_137# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X20 a_1000_81# a_798_107# a_1268_251# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X21 a_30_131# CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X22 VGND D a_642_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X23 a_2131_203# SET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X24 a_1989_515# a_2031_177# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X25 a_1000_81# SET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X26 VGND a_30_131# a_340_593# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X27 VPWR D a_642_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X28 VPWR a_798_107# a_1653_515# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X29 a_30_131# CLK VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X30 a_798_107# a_340_593# a_958_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X31 a_1787_137# a_30_131# a_1989_203# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__dfxbp_1 CLK D VGND VNB VPB VPWR Q Q_N
X0 a_1021_111# a_1063_85# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X1 a_1669_111# a_1711_85# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X2 VPWR a_865_111# a_1063_85# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X3 a_865_111# a_339_112# a_1021_111# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X4 a_1494_539# a_30_112# a_1669_111# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X5 VPWR D a_709_111# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X6 VPWR a_1494_539# a_1711_85# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X7 a_1063_85# a_339_112# a_1494_539# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X8 Q a_1711_85# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X9 VGND a_865_111# a_1063_85# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X10 a_1063_85# a_30_112# a_1494_539# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X11 VGND a_30_112# a_339_112# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X12 a_30_112# CLK VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X13 Q a_1711_85# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X14 a_2365_443# a_1711_85# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X15 a_2365_443# a_1711_85# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X16 VGND D a_709_111# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X17 VPWR a_30_112# a_339_112# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X18 a_709_111# a_339_112# a_865_111# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X19 VGND a_1494_539# a_1711_85# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X20 VPWR a_2365_443# Q_N VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X21 a_1021_539# a_1063_85# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X22 a_1669_539# a_1711_85# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X23 a_865_111# a_30_112# a_1021_539# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X24 a_1494_539# a_339_112# a_1669_539# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X25 a_30_112# CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X26 a_709_111# a_30_112# a_865_111# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X27 VGND a_2365_443# Q_N VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__dfxtp_1 CLK D VGND VNB VPB VPWR Q
X0 a_780_574# a_30_127# a_982_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X1 VPWR a_1455_543# a_1729_87# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X2 VGND a_1729_87# Q VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 a_1015_113# a_1024_371# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X4 VPWR a_780_574# a_1024_371# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X5 a_1455_543# a_339_559# a_1731_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X6 VGND a_1455_543# a_1729_87# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X7 a_780_574# a_339_559# a_1015_113# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X8 a_30_127# CLK VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X9 a_1455_543# a_30_127# a_1687_113# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X10 a_605_563# a_30_127# a_780_574# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X11 a_1024_371# a_30_127# a_1455_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X12 a_1024_371# a_339_559# a_1455_543# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X13 a_605_563# a_339_559# a_780_574# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X14 a_30_127# CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X15 VGND a_780_574# a_1024_371# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X16 VPWR a_1729_87# Q VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X17 VPWR D a_605_563# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X18 VGND a_30_127# a_339_559# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X19 VGND D a_605_563# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X20 a_982_543# a_1024_371# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X21 a_1687_113# a_1729_87# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X22 a_1731_543# a_1729_87# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X23 VPWR a_30_127# a_339_559# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__diode_2 DIODE VGND VNB VPB VPWR
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_11v0 pj=5.88e+06u area=6.072e+11p
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__dlclkp_1 CLK GATE VGND VNB VPB VPWR GCLK
X0 a_303_311# a_239_419# a_1027_159# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X1 a_189_159# a_231_71# a_303_311# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X2 VGND a_1438_171# GCLK VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 VGND GATE a_189_159# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X4 VGND a_303_311# a_1069_133# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X5 a_189_445# a_239_419# a_303_311# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X6 VPWR GATE a_189_445# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X7 a_239_419# a_231_71# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X8 VPWR a_1438_171# GCLK VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X9 a_1438_171# CLK VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X10 a_239_419# a_231_71# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X11 a_1027_457# a_1069_133# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X12 a_1591_171# CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X13 VPWR a_1069_133# a_1438_171# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X14 VPWR CLK a_231_71# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X15 a_303_311# a_231_71# a_1027_457# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X16 VPWR a_303_311# a_1069_133# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X17 VGND CLK a_231_71# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X18 a_1438_171# a_1069_133# a_1591_171# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X19 a_1027_159# a_1069_133# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__dlrtp_1 D GATE RESET_B VGND VNB VPB VPWR Q
X0 a_1096_491# a_1138_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X1 a_775_491# a_345_107# a_917_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X2 a_1096_107# a_1138_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X3 a_917_107# a_462_107# a_1096_491# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X4 a_775_107# a_462_107# a_917_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X5 VPWR a_917_107# a_1138_81# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X6 a_462_107# a_345_107# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X7 a_1138_81# a_917_107# a_1512_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X8 a_917_107# a_345_107# a_1096_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X9 a_462_107# a_345_107# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X10 VPWR a_1138_81# Q VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X11 a_1138_81# RESET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X12 a_32_107# D VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X13 VPWR a_32_107# a_775_491# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X14 VGND GATE a_345_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X15 a_32_107# D VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X16 VGND a_32_107# a_775_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X17 VGND a_1138_81# Q VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X18 VPWR GATE a_345_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X19 a_1512_107# RESET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__dlxtp_1 D GATE VGND VNB VPB VPWR Q
X0 a_650_107# a_384_107# a_806_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X1 a_30_443# GATE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X2 a_962_107# a_1004_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X3 VPWR D a_650_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X4 VGND D a_650_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X5 VGND a_806_107# Q VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X6 a_1014_587# a_1004_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X7 VPWR a_806_107# Q VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X8 a_806_107# a_30_443# a_962_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X9 a_1004_81# a_806_107# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X10 a_30_443# GATE VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X11 VPWR a_30_443# a_384_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X12 a_806_107# a_384_107# a_1014_587# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X13 a_650_107# a_30_443# a_806_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X14 a_1004_81# a_806_107# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X15 VGND a_30_443# a_384_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__einvn_1 A TE_B VGND VNB VPB VPWR Z
X0 VGND a_30_173# a_437_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X1 a_30_173# TE_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X2 a_437_107# A Z VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 VPWR TE_B a_413_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X4 a_30_173# TE_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X5 a_413_443# A Z VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__einvp_1 A TE VGND VNB VPB VPWR Z
X0 a_413_443# A Z VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 a_30_189# TE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X2 a_30_189# TE VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X3 VGND TE a_413_123# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 a_413_123# A Z VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X5 VPWR a_30_189# a_413_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__fill_1 VGND VNB VPB VPWR
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__fill_2 VGND VNB VPB VPWR
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__fill_4 VGND VNB VPB VPWR
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__fill_8 VGND VNB VPB VPWR
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__inv_1 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__inv_2 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X2 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__inv_4 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X4 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X5 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X6 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X7 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__inv_8 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X4 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X6 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X7 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X8 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X9 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X10 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X11 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X12 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X13 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X14 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X15 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__inv_16 A VGND VNB VPB VPWR Y
X0 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X1 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X6 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X7 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X8 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X9 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X10 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X11 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X12 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X13 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X14 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X15 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X16 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X17 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X18 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X19 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X20 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X21 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X22 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X23 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X24 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X25 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X26 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X27 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X28 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X29 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X30 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X31 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__lsbufhv2hv_hl_1 A LOWHVPWR VGND VNB VPB VPWR X
X0 X a_662_81# LOWHVPWR LOWHVPWR sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 LOWHVPWR A a_662_81# LOWHVPWR sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X2 X a_662_81# a_762_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 a_762_107# A a_662_81# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__lsbufhv2hv_lh_1 A LOWHVPWR VGND VNB VPB VPWR X
X0 a_847_1221# a_626_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 a_1353_107# a_935_141# a_779_141# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X2 VPWR a_1353_107# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X3 a_847_1221# a_626_141# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X4 a_1353_107# a_847_1221# a_1793_563# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=1e+06u
X5 a_1353_107# a_935_141# a_779_141# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X6 a_626_141# A LOWHVPWR LOWHVPWR sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X7 VGND a_626_141# a_847_1221# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X8 VGND a_1353_107# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X9 a_626_141# A a_779_141# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X10 LOWHVPWR a_626_141# a_935_141# LOWHVPWR sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X11 a_779_141# a_935_141# a_1353_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X12 a_847_1221# a_1353_107# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=1e+06u
X13 a_779_141# a_935_141# a_1353_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X14 VGND a_626_141# a_847_1221# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X15 a_779_141# a_626_141# a_935_141# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__lsbufhv2lv_1 A LVPWR VGND VNB VPB VPWR X

X1  VPWR		a_30_1337# 	a_30_207# 	VPB 	sky130_fd_pr__pfet_g5v0d10v5  w=420000u l=500000u
X10 VPWR       		A          	a_30_1337# 	VPB 	sky130_fd_pr__pfet_g5v0d10v5  w=420000u l=500000u
X11 a_30_1337# 		A 		VGND 		VNB 	sky130_fd_pr__nfet_g5v0d10v5  w=420000u l=500000u
X0  a_30_207# 		a_30_1337#      VGND 	VNB 	sky130_fd_pr__nfet_g5v0d10v5  w=420000u l=500000u
X3  a_389_1337#		a_30_1337# 	VGND 		VNB 	sky130_fd_pr__nfet_g5v0d10v5  w=750000u l=500000u
X4  a_389_1337#		a_30_1337# 	VGND 		VNB 	sky130_fd_pr__nfet_g5v0d10v5  w=750000u l=500000u
X7  VGND		a_30_207# 	a_389_141# 	VNB 	sky130_fd_pr__nfet_g5v0d10v5  w=750000u l=500000u
X13 a_389_141# 		a_30_207#       VGND      VNB     sky130_fd_pr__nfet_g5v0d10v5  w=750000u l=500000u
X8  a_389_141# 		a_30_207#       VGND      VNB     sky130_fd_pr__nfet_g5v0d10v5  w=750000u l=500000u
X9  a_389_141# 		a_30_207#       VGND      VNB     sky130_fd_pr__nfet_g5v0d10v5  w=750000u l=500000u
X14 VGND 		a_30_1337# 	a_389_1337#	VNB	sky130_fd_pr__nfet_g5v0d10v5  w=750000u l=500000u
X15 VGND 		a_30_1337# 	a_389_1337# 	VNB 	sky130_fd_pr__nfet_g5v0d10v5  w=750000u l=500000u
X5  X 			a_389_141# 	LVPWR 		LVPWR 	sky130_fd_pr__pfet_01v8_hvt   w=1.12e+06u l=150000u
X6  a_389_141# 		a_389_1337# 	LVPWR 		LVPWR 	sky130_fd_pr__pfet_01v8_hvt   w=1.12e+06u l=150000u
X12 LVPWR 		a_389_141# 	a_389_1337# 	LVPWR 	sky130_fd_pr__pfet_01v8_hvt   w=1.12e+06u l=150000u
X2  X 			a_389_141# 	VGND 	VNB 	sky130_fd_pr__nfet_01v8       w=740000u   l=150000u

.ends



******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__lsbufhv2lv_simple_1 A LVPWR VGND VNB VPB VPWR X
X0 X a_662_81# a_762_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X1 a_762_107# A a_662_81# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X2 X a_662_81# LVPWR LVPWR sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X3 LVPWR A a_662_81# LVPWR sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__lsbuflv2hv_1 A LVPWR VGND VNB VPB VPWR X
X0 VGND a_404_1133# a_504_1221# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 a_686_151# a_772_151# a_1197_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X2 a_1711_885# a_504_1221# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X3 a_1711_885# a_504_1221# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 a_404_1133# A a_686_151# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 VPWR a_1711_885# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X6 a_404_1133# A LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X7 VGND a_404_1133# a_504_1221# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X8 a_504_1221# a_404_1133# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X9 a_1197_107# a_504_1221# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=1e+06u
X10 a_686_151# a_772_151# a_1197_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X11 a_686_151# a_404_1133# a_772_151# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 LVPWR a_404_1133# a_772_151# LVPWR sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X13 a_686_151# a_772_151# a_1197_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X14 VGND a_404_1133# a_504_1221# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X15 a_504_1221# a_1197_107# a_1606_563# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=1e+06u
X16 a_504_1221# a_404_1133# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X17 VGND a_1711_885# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X18 a_1197_107# a_772_151# a_686_151# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X19 a_1197_107# a_772_151# a_686_151# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__lsbuflv2hv_clkiso_hlkg_3 A SLEEP_B LVPWR VGND VNB VPB VPWR X
X0 VPWR a_262_107# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X1 VGND a_528_1171# a_362_1243# VNB sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X2 a_362_133# a_528_1171# a_1472_1171# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X3 a_362_1243# a_528_1171# VGND VNB sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X4 a_362_1243# a_840_107# a_1410_571# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X5 a_1472_1171# a_528_1171# a_362_133# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X6 a_940_485# a_2092_381# a_1410_571# VPB sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X7 a_1472_1171# a_528_1171# LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X8 a_840_107# a_1472_1171# VGND VNB sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X9 VGND a_1472_1171# a_840_107# VNB sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X10 a_940_485# a_2092_381# a_1410_571# VPB sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X11 a_528_1171# a_3617_1198# LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X12 VGND a_528_1171# a_362_1243# VNB sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X13 X a_262_107# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X14 LVPWR a_3617_1198# a_528_1171# LVPWR sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X15 a_362_133# a_528_1171# a_1472_1171# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X16 a_1472_1171# a_528_1171# a_362_133# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X17 a_3617_1198# A LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X18 a_362_133# a_840_107# a_262_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
X19 X a_262_107# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X20 LVPWR a_3617_1198# a_528_1171# LVPWR sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X21 a_528_1171# a_3617_1198# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X22 a_262_107# a_840_107# a_362_133# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
X23 a_1410_571# a_2092_381# a_940_485# VPB sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X24 a_840_107# a_2092_381# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X25 a_1472_1171# a_528_1171# LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X26 a_362_133# a_262_107# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
X27 a_840_107# a_1472_1171# VGND VNB sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X28 VGND a_3617_1198# a_528_1171# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X29 LVPWR a_528_1171# a_1472_1171# LVPWR sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X30 a_2092_381# SLEEP_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X31 a_528_1171# a_3617_1198# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X32 VGND a_3617_1198# a_528_1171# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X33 LVPWR a_528_1171# a_1472_1171# LVPWR sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X34 a_940_485# a_840_107# a_262_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X35 a_362_1243# a_528_1171# VGND VNB sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X36 VGND VGND a_362_1243# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X37 VGND a_1472_1171# a_840_107# VNB sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X38 a_2092_381# SLEEP_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X39 a_528_1171# a_3617_1198# LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X40 a_3617_1198# A VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X41 LVPWR A a_3617_1198# LVPWR sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X42 VGND A a_3617_1198# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X43 X a_262_107# a_362_133# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
X44 a_262_107# a_840_107# a_940_485# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X45 a_1410_571# a_362_1243# a_840_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X46 a_1410_571# a_2092_381# a_940_485# VPB sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X47 X a_262_107# a_362_133# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__lsbuflv2hv_isosrchvaon_1 A SLEEP_B LVPWR VGND VNB VPB VPWR X
X0 a_176_993# a_229_967# a_341_485# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=2e+06u
X1 a_341_183# SLEEP_B a_507_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 X a_229_967# a_341_485# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X3 a_188_1293# a_553_1225# a_229_967# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
X4 a_341_183# A a_241_1225# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X5 a_188_1293# a_241_1225# a_176_993# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
X6 a_341_485# SLEEP_B a_507_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X7 a_188_1293# SLEEP_B a_341_183# VNB sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X8 a_553_1225# a_241_1225# LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X9 a_553_1225# a_241_1225# VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X10 a_341_183# SLEEP_B a_188_1293# VNB sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X11 a_176_993# a_241_1225# a_188_1293# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
X12 a_341_485# a_176_993# a_229_967# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=2e+06u
X13 X a_229_967# a_341_183# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X14 a_176_993# a_507_107# a_341_183# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=800000u
X15 LVPWR A a_241_1225# LVPWR sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X16 a_229_967# a_553_1225# a_188_1293# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__lsbuflv2hv_symmetric_1 A LVPWR VGND VNB VPB VPWR X
X0 a_1400_777# a_1406_429# a_1197_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 VGND a_1406_429# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 a_1406_429# a_816_1221# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X3 a_573_897# A a_686_151# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 a_573_897# A LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X5 a_1606_563# a_816_1221# a_1400_777# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=1e+06u
X6 VGND a_573_897# a_816_1221# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X7 a_816_1221# a_1400_777# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X8 a_816_1221# a_573_897# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X9 a_686_151# a_573_897# a_772_151# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 LVPWR a_573_897# a_772_151# LVPWR sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X11 a_686_151# a_772_151# a_1197_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X12 a_816_1221# a_1406_429# a_1606_563# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=1e+06u
X13 VPWR a_1400_777# a_816_1221# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X14 VPWR a_1406_429# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X15 a_1406_429# a_816_1221# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X16 a_1197_107# a_772_151# a_686_151# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X17 a_1400_777# a_1406_429# a_1606_563# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X18 a_1197_107# a_1406_429# a_1400_777# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__mux2_1 A0 A1 S VGND VNB VPB VPWR X
X0 X a_94_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X1 a_671_107# a_713_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X2 a_373_491# A0 a_94_81# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X3 X a_94_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X4 a_373_107# A1 a_94_81# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X5 a_94_81# A1 a_671_491# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X6 a_94_81# A0 a_671_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X7 VPWR S a_373_491# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X8 VPWR S a_713_81# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X9 a_671_491# a_713_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X10 VGND S a_373_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X11 VGND S a_713_81# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
X0 a_30_107# S0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X1 a_30_107# S0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X2 a_1097_627# a_1681_89# a_1669_615# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X3 a_1281_107# A0 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X4 a_955_627# a_30_107# a_1097_627# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X5 a_481_107# S0 a_637_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X6 a_1253_627# A0 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X7 a_983_107# S0 a_1097_627# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X8 VGND a_1669_615# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X9 a_481_107# a_30_107# a_637_627# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X10 a_637_627# A3 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X11 VPWR a_1669_615# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X12 a_1097_627# S1 a_1669_615# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X13 a_1681_89# S1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X14 VGND A2 a_339_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X15 a_339_107# a_30_107# a_481_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X16 VGND A1 a_983_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X17 VPWR A1 a_955_627# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X18 VPWR A2 a_339_627# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X19 a_1669_615# a_1681_89# a_481_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X20 a_1097_627# a_30_107# a_1281_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X21 a_339_627# S0 a_481_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X22 a_1097_627# S0 a_1253_627# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X23 a_1681_89# S1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X24 a_637_107# A3 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X25 a_1669_615# S1 a_481_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__nand2_1 A B VGND VNB VPB VPWR Y
X0 VPWR B Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 VGND B a_233_111# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 a_233_111# A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__nand3_1 A B C VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 VGND C a_243_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 VPWR C Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X3 a_385_107# A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 a_243_107# B a_385_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X5 Y B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__nor2_1 A B VGND VNB VPB VPWR Y
X0 VPWR A a_251_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 Y B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 a_251_443# B Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__nor3_1 A B C VGND VNB VPB VPWR Y
X0 a_347_443# C Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 Y B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 a_205_443# B a_347_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X3 VGND C Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X5 VPWR A a_205_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
X0 a_83_87# A2 a_602_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 a_460_107# A2 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 a_83_87# B1 a_460_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 X a_83_87# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 VGND A1 a_460_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X5 X a_83_87# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X6 a_602_443# A1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X7 VPWR B1 a_83_87# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
X0 a_30_107# A1 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X1 VGND A2 a_30_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 a_205_443# A2 Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X3 a_30_107# B1 Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 Y B1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X5 VPWR A1 a_205_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 a_354_107# A2 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X1 a_87_81# A2 a_831_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X2 X a_87_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 VGND A1 a_354_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 X a_87_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X5 VPWR B1 a_533_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X6 a_354_107# B1 a_87_81# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X7 a_831_443# A1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X8 a_87_81# B2 a_354_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X9 a_533_443# B2 a_87_81# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
X0 a_207_443# B2 Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 a_520_443# A1 VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X2 Y B2 a_36_113# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 VGND A1 a_36_113# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 VPWR B1 a_207_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X5 a_36_113# A2 VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X6 a_36_113# B1 Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X7 Y A2 a_520_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__or2_1 A B VGND VNB VPB VPWR X
X0 VPWR a_84_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 a_241_443# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X2 a_84_443# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X3 VGND B a_84_443# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X4 a_84_443# B a_241_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X5 VGND a_84_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__or3_1 A B C VGND VNB VPB VPWR X
X0 VGND a_30_107# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X1 VPWR a_30_107# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X2 a_30_107# C VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X3 a_30_107# C a_190_464# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X4 a_341_464# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X5 a_30_107# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X6 VGND B a_30_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X7 a_190_464# B a_341_464# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__probe_p_8 A VGND VNB VPB VPWR X
X0 a_45_443# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X3 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X5 VGND A a_45_443# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X6 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X7 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X8 a_45_443# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X9 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X10 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X11 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X12 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X13 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X14 a_45_443# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X15 VPWR A a_45_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X16 a_45_443# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X17 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X18 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X19 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X20 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X21 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__probec_p_8 A VGND VNB VPB VPWR X
X0 a_45_443# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X3 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X5 VGND A a_45_443# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X6 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X7 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X8 a_45_443# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X9 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X10 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X11 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X12 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X13 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X14 a_45_443# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X15 VPWR A a_45_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X16 a_45_443# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X17 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X18 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X19 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X20 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X21 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__schmittbuf_1 A VGND VNB VPB VPWR X
X0 a_117_181# A a_231_463# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X1 a_117_181# A a_217_207# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X2 a_78_463# VGND VNB sky130_fd_pr__res_generic_nd__hv w=290000u l=1.355e+06u
X3 a_64_207# VPWR VPB sky130_fd_pr__res_generic_pd__hv w=290000u l=3.11e+06u
X4 a_231_463# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X5 a_64_207# a_117_181# a_217_207# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X6 VGND a_117_181# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X7 VPWR a_117_181# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X8 a_217_207# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X9 a_78_463# a_117_181# a_231_463# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__sdfrbp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q Q_N
X0 a_3098_107# a_2624_107# a_2841_81# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X1 VPWR SCD a_794_655# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X2 a_1999_126# a_2014_537# a_2141_126# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X3 VGND a_2624_107# Q_N VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 a_1972_659# a_2014_537# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X5 a_2871_543# a_2841_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X6 VGND CLK a_1290_126# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X7 a_2799_107# a_2841_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X8 a_2624_107# a_1290_126# a_2799_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X9 VPWR a_1290_126# a_1569_126# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X10 a_339_655# D a_496_655# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X11 a_1816_659# a_1290_126# a_1972_659# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X12 VPWR a_1816_659# a_2014_537# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X13 VPWR RESET_B a_2841_81# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X14 a_794_655# a_222_131# a_339_655# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X15 a_339_655# SCE a_816_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X16 VPWR CLK a_1290_126# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X17 VPWR RESET_B a_1816_659# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X18 VGND a_1816_659# a_2014_537# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X19 VGND SCE a_222_131# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X20 a_2841_81# a_2624_107# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X21 a_3613_443# a_2624_107# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X22 a_2141_126# RESET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X23 a_361_107# D a_518_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X24 a_496_655# SCE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X25 a_339_655# RESET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X26 VGND a_1290_126# a_1569_126# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X27 a_2014_537# a_1569_126# a_2624_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X28 a_2624_107# a_1569_126# a_2871_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X29 a_518_107# a_222_131# a_339_655# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X30 a_2014_537# a_1290_126# a_2624_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X31 a_361_107# RESET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X32 VGND RESET_B a_3098_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X33 a_1816_659# a_1569_126# a_1999_126# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X34 a_3613_443# a_2624_107# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X35 VPWR a_3613_443# Q VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X36 VPWR SCE a_222_131# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X37 a_339_655# a_1290_126# a_1816_659# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X38 VPWR a_2624_107# Q_N VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X39 VGND a_3613_443# Q VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X40 a_339_655# a_1569_126# a_1816_659# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X41 a_816_107# SCD a_361_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__sdfrtp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
X0 VPWR SCE a_116_451# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X1 VGND SCE a_116_451# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X2 a_1510_100# a_1212_471# a_2360_115# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 a_2574_543# a_2616_417# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X4 VGND RESET_B a_2904_181# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X5 a_1212_100# CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X6 VGND a_3417_443# Q VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X7 a_294_126# SCE a_65_649# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X8 VPWR a_3417_443# Q VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X9 a_1610_126# RESET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X10 a_3417_443# a_2360_115# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X11 a_524_649# D a_65_649# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X12 a_2360_115# a_1212_100# a_2539_181# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X13 a_137_126# RESET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X14 a_2539_181# a_2616_417# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X15 a_222_649# SCD VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X16 VPWR CLK a_1212_100# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X17 a_65_649# RESET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X18 a_1468_641# a_1510_100# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X19 VPWR RESET_B a_2616_417# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X20 a_3417_443# a_2360_115# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X21 a_65_649# a_116_451# a_592_126# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X22 a_1312_126# a_1212_100# a_1468_641# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X23 VPWR a_1312_126# a_1510_100# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X24 VGND a_1312_126# a_1510_100# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X25 a_1468_126# a_1510_100# a_1610_126# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X26 a_2904_181# a_2360_115# a_2616_417# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X27 VPWR SCE a_524_649# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X28 a_65_649# a_1212_471# a_1312_126# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X29 VPWR RESET_B a_1312_126# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X30 a_2360_115# a_1212_471# a_2574_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X31 a_1212_471# a_1212_100# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X32 a_1312_126# a_1212_471# a_1468_126# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X33 a_1212_471# a_1212_100# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X34 a_137_126# SCD a_294_126# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X35 a_65_649# a_116_451# a_222_649# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X36 a_2616_417# a_2360_115# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X37 a_65_649# a_1212_100# a_1312_126# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X38 a_592_126# D a_137_126# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X39 a_1510_100# a_1212_100# a_2360_115# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__sdfsbp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
X0 a_641_569# SCD VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X1 VGND a_972_569# a_1243_116# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X2 a_2501_543# a_972_569# a_2715_173# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X3 a_485_569# a_1243_116# a_1513_120# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X4 a_1711_94# a_1513_120# a_2077_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X5 VGND D a_348_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X6 VPWR a_2501_543# Q_N VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X7 a_348_107# a_30_569# a_485_569# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X8 a_2857_173# SET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X9 VPWR CLK a_972_569# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X10 a_343_569# D a_485_569# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X11 a_1513_120# a_972_569# a_1710_556# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X12 a_2394_107# a_1243_116# a_2501_543# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X13 a_2501_543# a_1243_116# a_2687_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X14 a_2729_463# a_2501_543# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X15 a_3609_173# a_2501_543# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X16 VPWR a_3609_173# Q VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X17 VPWR SET_B a_2501_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X18 a_646_107# SCD VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X19 a_3609_173# a_2501_543# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X20 a_485_569# a_30_569# a_641_569# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X21 a_30_569# SCE VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X22 VPWR a_972_569# a_1243_116# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X23 VGND a_3609_173# Q VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X24 a_2729_463# a_2501_543# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X25 VGND CLK a_972_569# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X26 a_1669_120# a_1711_94# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X27 a_2715_173# a_2729_463# a_2857_173# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X28 a_30_569# SCE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X29 a_1711_94# SET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X30 a_1513_120# a_1243_116# a_1669_120# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X31 VPWR SCE a_343_569# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X32 a_2687_543# a_2729_463# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X33 VGND a_2501_543# Q_N VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X34 a_2359_543# a_972_569# a_2501_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X35 a_1710_556# a_1711_94# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X36 a_485_569# a_972_569# a_1513_120# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X37 a_485_569# SCE a_646_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X38 a_2077_107# SET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X39 VPWR a_1513_120# a_1711_94# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X40 VPWR a_1513_120# a_2359_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X41 VGND a_1513_120# a_2394_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__sdfstp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
X0 VGND a_2477_543# a_2698_421# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X1 a_2352_107# a_1201_123# a_2477_543# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 VGND a_3321_173# Q VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 a_30_107# SCE VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X4 a_1471_113# a_1201_123# a_1627_113# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X5 VPWR SCE a_339_569# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X6 VPWR a_1471_113# a_1669_87# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X7 a_1471_113# a_935_107# a_1686_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X8 VGND CLK a_935_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X9 a_2477_543# a_935_107# a_2669_173# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X10 a_339_569# D a_481_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X11 a_481_107# a_1201_123# a_1471_113# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X12 VPWR a_1471_113# a_2335_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X13 a_481_107# a_935_107# a_1471_113# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X14 a_1669_87# SET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X15 a_481_107# SCE a_637_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X16 a_2812_173# SET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X17 VPWR CLK a_935_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X18 a_637_569# SCD VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X19 a_2656_543# a_2698_421# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X20 VGND a_1471_113# a_2352_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X21 a_1686_543# a_1669_87# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X22 a_30_107# SCE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X23 a_2035_107# SET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X24 a_1627_113# a_1669_87# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X25 VPWR SET_B a_2477_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X26 VGND D a_339_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X27 a_1669_87# a_1471_113# a_2035_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X28 a_339_107# a_30_107# a_481_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X29 VPWR a_3321_173# Q VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X30 a_2698_421# a_2477_543# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X31 VGND a_935_107# a_1201_123# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X32 a_2669_173# a_2698_421# a_2812_173# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X33 a_3321_173# a_2477_543# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X34 a_3321_173# a_2477_543# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X35 a_481_107# a_30_107# a_637_569# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X36 VPWR a_935_107# a_1201_123# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X37 a_2477_543# a_1201_123# a_2656_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X38 a_2335_543# a_935_107# a_2477_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X39 a_637_107# SCD VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__sdfxbp_1 CLK D SCD SCE VGND VNB VPB VPWR Q Q_N
X0 a_1528_579# a_1570_457# a_1124_81# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X1 a_425_107# SCE a_567_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X2 VGND a_2518_445# a_2789_147# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 a_2365_445# a_2789_147# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X4 VGND CLK a_1570_457# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X5 a_30_515# SCE VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X6 a_567_107# a_30_515# a_723_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X7 VPWR a_2789_147# a_3531_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X8 a_2518_445# a_1570_457# a_2747_173# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X9 a_268_659# a_30_515# a_567_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X10 VPWR CLK a_1570_457# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X11 a_567_107# a_1570_457# a_1124_81# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X12 VGND SCD a_425_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X13 a_567_107# D a_581_659# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X14 VGND a_1067_107# a_1454_173# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X15 VGND a_3531_107# Q_N VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X16 a_268_659# SCD VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X17 a_1067_107# a_1726_453# a_2518_445# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X18 a_1067_107# a_1124_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X19 a_1124_81# a_1726_453# a_567_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X20 VPWR a_3531_107# Q_N VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X21 a_1726_453# a_1570_457# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X22 a_723_107# D VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X23 Q a_2789_147# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X24 a_1124_81# a_1726_453# a_1454_173# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X25 a_30_515# SCE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X26 a_1067_107# a_1124_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X27 a_2747_173# a_2789_147# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X28 VGND a_2789_147# a_3531_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X29 VPWR a_2518_445# a_2789_147# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X30 Q a_2789_147# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X31 a_2365_445# a_1726_453# a_2518_445# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X32 a_1726_453# a_1570_457# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X33 VPWR a_1067_107# a_1528_579# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X34 VPWR SCE a_581_659# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X35 a_2518_445# a_1570_457# a_1067_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__sdfxtp_1 CLK D SCD SCE VGND VNB VPB VPWR Q
X0 VPWR a_2123_543# a_2352_81# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X1 VPWR CLK a_938_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X2 a_342_107# a_30_593# a_484_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X3 a_2123_543# a_938_107# a_2310_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X4 a_484_107# a_30_593# a_641_593# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X5 Q a_2352_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X6 a_1688_81# a_1204_107# a_2123_543# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X7 a_30_593# SCE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X8 a_484_107# SCE a_640_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X9 a_1490_107# a_1204_107# a_1646_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X10 a_1490_107# a_938_107# a_1646_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X11 VPWR SCE a_343_593# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X12 a_2123_543# a_1204_107# a_2302_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X13 VGND a_938_107# a_1204_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X14 a_1688_81# a_938_107# a_2123_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X15 a_30_593# SCE VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X16 VGND D a_342_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X17 VGND CLK a_938_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X18 a_484_107# a_938_107# a_1490_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X19 a_2310_107# a_2352_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X20 a_484_107# a_1204_107# a_1490_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X21 a_2302_543# a_2352_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X22 a_641_593# SCD VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X23 a_640_107# SCD VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X24 a_1646_107# a_1688_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X25 VGND a_1490_107# a_1688_81# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X26 VPWR a_1490_107# a_1688_81# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X27 Q a_2352_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X28 a_1646_543# a_1688_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X29 a_343_593# D a_484_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X30 VPWR a_938_107# a_1204_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X31 VGND a_2123_543# a_2352_81# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__sdlclkp_1 CLK GATE SCE VGND VNB VPB VPWR GCLK
X0 VGND a_1630_171# GCLK VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X1 a_1783_171# CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X2 a_58_159# a_423_71# a_495_311# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X3 VPWR a_1261_133# a_1630_171# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X4 VPWR SCE a_219_457# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X5 VPWR CLK a_423_71# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X6 VPWR a_1630_171# GCLK VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X7 a_431_431# a_423_71# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X8 VPWR a_495_311# a_1261_133# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X9 VGND CLK a_423_71# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X10 a_1630_171# a_1261_133# a_1783_171# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X11 a_58_159# SCE VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X12 a_219_457# GATE a_58_159# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X13 a_495_311# a_423_71# a_1219_457# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X14 a_1219_457# a_1261_133# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X15 VGND a_495_311# a_1261_133# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X16 a_58_159# a_431_431# a_495_311# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X17 a_1630_171# CLK VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X18 VGND GATE a_58_159# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X19 a_495_311# a_431_431# a_1219_159# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X20 a_431_431# a_423_71# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X21 a_1219_159# a_1261_133# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__sdlxtp_1 D GATE SCD SCE VGND VNB VPB VPWR Q
X0 a_1724_593# a_1678_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X1 a_1480_107# a_944_107# a_1636_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X2 a_489_107# SCE a_645_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X3 a_1678_81# a_1480_107# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X4 a_489_107# a_30_587# a_660_587# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X5 a_489_107# a_1214_107# a_1480_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X6 VGND D a_347_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X7 a_1480_107# a_1214_107# a_1724_593# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X8 VPWR a_944_107# a_1214_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X9 a_489_107# a_944_107# a_1480_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X10 VPWR SCE a_362_587# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X11 VPWR a_1480_107# Q VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X12 VPWR GATE a_944_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X13 a_1636_107# a_1678_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X14 VGND GATE a_944_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X15 VGND a_944_107# a_1214_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X16 a_660_587# SCD VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X17 a_645_107# SCD VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X18 a_30_587# SCE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X19 a_30_587# SCE VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X20 a_347_107# a_30_587# a_489_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X21 a_1678_81# a_1480_107# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X22 VGND a_1480_107# Q VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X23 a_362_587# D a_489_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__xnor2_1 A B VGND VNB VPB VPWR Y
X0 VGND A a_523_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X1 VPWR A a_539_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X2 VPWR B a_30_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X3 a_539_443# B Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X4 a_222_107# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X5 a_523_107# a_30_107# Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X6 a_523_107# B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X7 Y a_30_107# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X8 a_30_107# B a_222_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X9 a_30_107# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__xor2_1 A B VGND VNB VPB VPWR X
X0 X a_30_443# a_531_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 VGND B a_30_443# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 a_30_443# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 a_30_443# B a_187_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X4 a_617_107# B X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X5 a_187_443# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X6 a_531_443# B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X7 X a_30_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X8 VPWR A a_531_443# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X9 VGND A a_617_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
.ends


******* EOF

** End of included library ./pdk/sky130_fd_sc_hvl.spice
** Start of included library ./pdk/sky130_fd_sc_hd.spice
* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 a_489_413# B2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 VGND A1_N a_226_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_76_199# B2 a_556_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VPWR A1_N a_226_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_226_297# A2_N a_226_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 VGND a_226_47# a_76_199# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 X a_76_199# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 X a_76_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_76_199# a_226_47# a_489_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 a_226_47# A2_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VPWR B1 a_489_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 a_556_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 VGND A1_N a_313_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 X a_82_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_82_21# a_313_47# a_574_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X3 a_82_21# B2 a_646_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VGND a_313_47# a_82_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VPWR a_82_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VPWR B1 a_574_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 a_574_369# B2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X8 VPWR A1_N a_313_297# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 a_313_297# A2_N a_313_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X10 VGND a_82_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_646_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 X a_82_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_313_47# A2_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 VGND A2_N a_415_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VGND a_193_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VGND a_415_21# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR a_193_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VGND a_193_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_193_47# a_415_21# a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_415_21# A2_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_109_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_193_47# a_415_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 X a_193_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VGND A1_N a_415_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VPWR a_193_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_193_47# B2 a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_717_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_109_47# B2 a_193_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_27_297# B2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 VPWR A1_N a_717_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 VGND B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 a_415_21# A2_N a_717_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_27_297# a_415_21# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 VPWR B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 a_415_21# A1_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 a_717_297# A2_N a_415_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X24 X a_193_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 X a_193_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 X a_193_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
X0 a_109_297# A2_N a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_481_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 Y B2 a_481_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 Y a_109_47# a_397_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VPWR B1 a_397_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_397_297# B2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_109_47# A2_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VGND A1_N a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VPWR A1_N a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VGND a_109_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
X0 a_136_47# B2 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VPWR B2 a_54_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_442_21# A2_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 Y a_442_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VGND A2_N a_442_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VGND A1_N a_442_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_54_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VGND a_442_21# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_662_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_442_21# A1_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_136_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VPWR B1 a_54_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VPWR A1_N a_662_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 Y a_442_21# a_54_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_442_21# A2_N a_662_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 Y B2 a_136_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_54_297# B2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 VGND B1 a_136_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 a_54_297# a_442_21# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_662_297# A2_N a_442_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
X0 Y a_751_21# a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VPWR A1_N a_1139_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_751_21# A2_N a_1139_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 Y B2 a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VGND A1_N a_751_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 Y B2 a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_1139_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_751_21# A2_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_27_297# a_751_21# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VPWR B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_109_47# B2 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VGND A2_N a_751_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 Y a_751_21# a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 VGND a_751_21# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_751_21# A2_N a_1139_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 VGND A2_N a_751_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 a_27_297# B2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 a_27_297# a_751_21# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_109_47# B2 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_1139_297# A2_N a_751_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 Y a_751_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 a_751_21# A1_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 Y a_751_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 VGND a_751_21# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 VGND B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 a_109_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X28 VGND B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 VGND A1_N a_751_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 a_27_297# B2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X31 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X32 a_1139_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X33 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X34 a_1139_297# A2_N a_751_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X35 a_109_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X36 a_751_21# A1_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X37 a_751_21# A2_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X38 VPWR B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X39 VPWR A1_N a_1139_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
X0 VPWR a_215_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_215_297# a_27_413# a_298_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VPWR A2 a_298_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_298_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_215_297# A1 a_382_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_27_413# B1_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_27_413# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VGND a_215_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_382_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VGND a_27_413# a_215_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
X0 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_79_21# A1 a_581_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VPWR B1_N a_297_93# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 VGND a_297_93# a_79_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_485_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_581_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_79_21# a_297_93# a_485_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VPWR A2 a_485_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 VGND B1_N a_297_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
X0 a_861_47# A1 a_205_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_205_21# A1 a_1021_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_205_21# a_42_47# a_603_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VPWR A1 a_603_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_42_47# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VPWR a_205_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 X a_205_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_603_297# a_42_47# a_205_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_603_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 X a_205_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VPWR A2 a_603_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_205_21# a_42_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VPWR a_205_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 X a_205_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 VGND A2 a_861_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_1021_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VGND a_42_47# a_205_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 VGND a_205_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 X a_205_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 a_42_47# B1_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_603_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 VGND a_205_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a21boi_0 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 a_27_47# B1_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_400_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_300_369# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X3 Y a_27_47# a_300_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X4 VGND a_27_47# Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 Y A1 a_400_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VPWR A2 a_300_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 a_27_47# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 a_384_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VGND a_27_413# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_300_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 Y a_27_413# a_300_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_27_413# B1_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 Y A1 a_384_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_27_413# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VPWR A2 a_300_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 Y A1 a_637_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_61_47# B1_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 Y a_61_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VGND A2 a_479_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_217_297# a_61_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_217_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_637_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 Y a_61_47# a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VPWR A1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 VGND a_61_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_479_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VPWR B1_N a_61_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 a_223_297# a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_223_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_658_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR A2 a_223_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VGND A2 a_658_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_658_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR A1 a_223_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_658_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VGND a_27_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 Y A1 a_658_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_223_297# a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 Y a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 Y a_27_47# a_223_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VGND A2 a_658_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_223_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_658_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_223_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 VPWR A1 a_223_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 VGND a_27_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 Y A1 a_658_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_27_47# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 Y a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 Y a_27_47# a_223_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 a_27_47# B1_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 VPWR A2 a_223_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 a_223_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
X0 a_384_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 X a_81_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_81_21# B1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VGND B1 a_81_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_299_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VPWR A2 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 X a_81_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_81_21# A1 a_384_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
X0 a_80_199# A1 a_458_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 X a_80_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VPWR a_80_199# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VGND a_80_199# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VGND B1 a_80_199# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 X a_80_199# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR A2 a_386_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_458_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_80_199# B1 a_386_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_386_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
X0 VPWR A2 a_483_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VGND a_84_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_483_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_741_47# A1 a_84_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_84_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VGND A2 a_741_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR a_84_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VGND B1 a_84_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 X a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_84_21# B1 a_483_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 X a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 VPWR a_84_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_483_297# B1 a_84_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_483_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 VGND a_84_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_901_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 X a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 X a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 a_84_21# A1 a_901_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 VPWR A1 a_483_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
X0 a_199_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_113_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 Y B1 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VPWR A2 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 Y A1 a_199_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
X0 VGND A2 a_114_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_285_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_114_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 Y A1 a_285_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
X0 VGND A2 a_462_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 Y B1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_28_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_28_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_28_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VPWR A1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VPWR A1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 Y B1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_28_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 VPWR A2 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_28_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_462_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_28_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 VPWR A2 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 VGND A2 a_462_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 a_462_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 Y A1 a_462_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 a_462_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 a_462_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 Y A1 a_462_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 a_109_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VPWR A1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_373_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_109_47# B1 a_27_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_27_297# A1 a_373_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VGND B2 a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_27_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_109_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_109_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_109_47# B1 a_27_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR A1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VGND B2 a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_27_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_27_297# A1 a_381_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_109_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_381_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 a_484_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 X a_96_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_96_21# B2 a_484_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VGND B2 a_566_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VGND a_96_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VPWR a_96_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VPWR A2 a_484_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_918_47# A1 a_96_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 X a_96_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VPWR a_96_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_484_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 X a_96_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VGND a_96_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_918_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VPWR A1 a_484_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_96_21# B1 a_566_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VGND A2 a_918_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 a_484_297# B2 a_96_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 a_96_21# A1 a_918_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 a_484_297# B1 a_96_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 a_566_47# B1 a_96_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 a_96_21# B1 a_484_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 a_566_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 X a_96_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
X0 a_109_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_109_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VPWR A1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_381_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VGND B2 a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 Y B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 Y A1 a_381_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_109_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
X0 VGND A2 a_467_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 Y A1 a_467_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VPWR A1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_467_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_467_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_109_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 Y B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_109_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_109_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
X0 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_803_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_803_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_803_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VGND A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 a_803_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X24 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 Y A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 VGND A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X30 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X31 Y A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 a_80_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 X a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_209_47# A2 a_303_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 X a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_303_47# A1 a_80_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VPWR A1 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_209_297# B1 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VGND A3 a_209_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_209_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VPWR A3 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 a_277_47# A2 a_361_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_361_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_79_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VGND A3 a_277_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VPWR A1 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_277_297# B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VPWR A3 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_277_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 VGND B1 a_277_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_361_47# A2 a_445_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_277_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 X a_277_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 X a_277_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_277_47# A1 a_361_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_277_47# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VPWR a_277_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 X a_277_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VGND a_277_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VPWR a_277_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 VGND a_277_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_193_47# A1 a_277_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_27_297# B1 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 X a_277_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_109_47# A2 a_193_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 VGND A3 a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 a_445_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
X0 a_109_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_181_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VPWR A1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_109_47# A2 a_181_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VGND A3 a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR A3 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_109_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
X0 a_277_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_277_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_27_47# A2 a_277_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 Y A1 a_277_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
X0 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 Y A1 a_445_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_27_47# A2 a_445_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_27_47# A2 a_445_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 Y A1 a_445_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_445_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X24 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 a_445_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 a_445_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X30 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X31 a_445_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 a_93_21# B2 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 X a_93_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_250_297# B1 a_93_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_256_47# A2 a_346_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 X a_93_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VGND A3 a_256_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_93_21# B1 a_584_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VPWR A1 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_346_47# A1 a_93_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_250_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VPWR A3 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_584_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 a_549_47# A2 a_665_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VGND B2 a_352_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_299_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_21_199# B1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_299_297# B2 a_21_199# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_352_47# B1 a_21_199# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_21_199# A1 a_549_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_299_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 X a_21_199# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VGND a_21_199# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VPWR A2 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 X a_21_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VPWR a_21_199# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_665_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 a_445_297# B2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_635_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_79_21# B1 a_1142_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VGND A3 a_445_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_445_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_445_47# A2 a_635_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_1142_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_445_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_445_297# B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_635_47# A2 a_445_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VGND B2 a_1142_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VPWR A1 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 a_445_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 a_1142_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 a_445_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 VPWR A3 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 a_79_21# B1 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X24 a_79_21# B2 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 a_79_21# A1 a_635_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 VPWR A2 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
X0 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_309_47# A2 a_383_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_109_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_383_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 Y A1 a_309_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VGND B2 a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
X0 a_730_47# A2 a_478_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 Y A1 a_478_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VGND A3 a_730_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_478_47# A2 a_730_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_730_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 a_478_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
X0 a_803_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_803_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VGND A3 a_1249_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_1249_47# A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_1249_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 a_1249_47# A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X24 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X28 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 VGND A3 a_1249_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X31 a_803_47# A2 a_1249_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X32 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X33 a_803_47# A2 a_1249_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X34 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X35 Y A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X36 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X37 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X38 a_1249_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X39 Y A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
X0 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VPWR A4 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_79_21# B1 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VPWR A2 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_297_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_297_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_465_47# A3 a_561_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_561_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_381_47# A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_79_21# A1 a_381_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
X0 a_549_47# A2 a_665_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VPWR A3 a_381_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_381_297# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_79_21# B1 a_381_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_465_47# A3 a_549_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VPWR A1 a_381_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VGND A4 a_465_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_381_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_79_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_665_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
X0 a_467_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_889_47# A3 a_1079_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_639_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR A1 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VPWR A2 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_1079_47# A3 a_889_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_467_297# B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_467_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_467_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VPWR A3 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_1079_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_79_21# B1 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_889_47# A2 a_639_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_79_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_467_297# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 VPWR A4 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 a_639_47# A2 a_889_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X24 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 a_79_21# A1 a_639_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 VGND A4 a_1079_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
X0 a_336_47# A2 a_428_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_109_297# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_236_47# A3 a_336_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_428_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VGND A4 a_236_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VPWR A3 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_109_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VPWR A1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a41oi_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
X0 a_317_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_149_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_567_47# A2 a_317_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR A4 a_149_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_149_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_149_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_149_297# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_757_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 Y B1 a_149_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VPWR A1 a_149_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VPWR A3 a_149_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_317_47# A2 a_567_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_757_47# A3 a_567_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VPWR A2 a_149_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_567_47# A3 a_757_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_149_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 Y A1 a_317_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 VGND A4 a_757_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
X0 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 Y A1 a_493_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VGND A4 a_1269_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 Y A1 a_493_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_493_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VPWR A4 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_1269_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_27_297# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_27_297# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_911_47# A2 a_493_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_911_47# A3 a_1269_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_911_47# A2 a_493_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 a_911_47# A3 a_1269_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 VPWR A4 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 a_493_47# A2 a_911_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 a_493_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 a_1269_47# A3 a_911_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X28 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X29 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 VGND A4 a_1269_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X32 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X33 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X34 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X35 a_1269_47# A3 a_911_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X36 a_1269_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X37 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X38 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X39 a_493_47# A2 a_911_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 VGND A2 a_300_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 X a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 X a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_300_47# A1 a_80_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_80_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_472_297# C1 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VGND C1 a_80_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VPWR A1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_217_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_217_297# B1 a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_299_297# B1 a_585_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_585_297# C1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_348_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VGND A2 a_348_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_79_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VGND C1 a_79_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 a_555_297# C1 a_79_204# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_473_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_1123_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_79_204# C1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VPWR A1 a_473_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 X a_79_204# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VPWR a_79_204# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_951_47# A1 a_79_204# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VGND C1 a_79_204# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VGND a_79_204# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VGND A2 a_951_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_727_297# B1 a_473_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 X a_79_204# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VGND a_79_204# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_79_204# C1 a_727_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 VGND B1 a_79_204# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_79_204# A1 a_1123_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 a_473_297# B1 a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 VPWR a_79_204# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 X a_79_204# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_473_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 VPWR A2 a_473_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 X a_79_204# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 a_79_204# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
X0 VGND A2 a_139_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_311_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VPWR A1 a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_56_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_56_297# B1 a_311_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_139_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
X0 a_292_297# B1 a_37_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_37_297# B1 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VPWR A2 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VGND A2 a_485_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_485_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 Y A1 a_485_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_485_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VPWR A1 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_292_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 Y C1 a_37_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_37_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_292_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
X0 Y C1 a_781_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 Y A1 a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 Y A1 a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_27_297# B1 a_949_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_109_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_781_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_949_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_781_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_1301_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_27_297# B1 a_781_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 a_109_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 VGND A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 a_109_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 Y C1 a_1301_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 VGND A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X28 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X29 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X30 a_109_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 VPWR A1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_193_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_205_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_465_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_27_47# A1 a_465_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_193_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_27_47# C1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_27_47# C1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_109_297# B2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VGND B2 a_205_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 VPWR A1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_193_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_205_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_465_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_27_47# A1 a_465_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_193_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_27_47# C1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_27_47# C1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_109_297# B2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VGND B2 a_205_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 a_79_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_79_21# C1 a_804_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_804_297# B2 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VGND A2 a_445_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_79_21# B1 a_1053_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_445_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_445_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_445_297# B2 a_804_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_445_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VPWR A1 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_445_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VGND B2 a_1053_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_79_21# A1 a_445_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_445_297# B1 a_804_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_1053_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 a_804_297# B1 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 VPWR A2 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X24 VGND C1 a_79_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 a_804_297# C1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 a_1053_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
X0 VGND B2 a_204_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_465_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VPWR A1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_204_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 Y A1 a_465_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_193_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 Y C1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_193_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_109_297# B2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
X0 VPWR A1 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_383_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_735_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR A2 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_27_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 Y A1 a_735_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_301_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND B2 a_383_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VGND A2 a_735_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_27_297# B1 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_27_297# B2 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_301_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_301_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_735_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_383_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_301_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 Y B1 a_383_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 Y C1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
X0 a_471_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_1241_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 Y C1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 Y C1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_27_297# B1 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_471_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_27_297# B1 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VGND A2 a_1241_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_27_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_471_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_27_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_453_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_471_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 a_471_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 Y A1 a_1241_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 VGND A2 a_1241_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 VGND B2 a_453_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_471_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 VGND B2 a_453_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 a_453_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 VPWR A1 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X24 VPWR A1 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 a_453_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 a_1241_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 a_1241_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 a_27_297# B2 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X30 VPWR A2 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X31 a_471_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X32 a_1241_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X33 a_471_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X34 VPWR A2 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X35 Y B1 a_453_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X36 a_27_297# B2 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X37 Y B1 a_453_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X38 Y A1 a_1241_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X39 a_453_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a222oi_1 A1 A2 B1 B2 C1 C2 VGND VNB VPB VPWR Y
X0 VGND B2 a_393_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X1 VPWR A2 a_311_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_109_297# B1 a_311_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_311_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_311_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_109_47# C2 VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X6 Y A1 a_561_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X7 a_561_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X8 a_393_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X9 Y C1 a_109_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X10 Y C1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_109_297# C2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 VPWR A1 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VGND A3 a_208_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_75_199# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_544_297# C1 a_75_199# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_201_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 X a_75_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_208_47# A2 a_315_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VPWR A3 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND C1 a_75_199# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 X a_75_199# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_315_47# A1 a_75_199# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_201_297# B1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 a_319_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_79_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VGND A3 a_319_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_319_297# B1 a_635_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_319_47# A2 a_417_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_635_297# C1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_417_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VPWR A1 a_319_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VGND C1 a_79_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VPWR A3 a_319_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VPWR A1 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_109_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_277_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_277_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_109_47# A1 a_1059_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VPWR A2 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_861_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_1059_47# A2 a_861_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VGND B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VGND A3 a_861_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_277_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 a_109_47# C1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 a_1059_47# A1 a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 a_27_297# B1 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 VGND C1 a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 VPWR A3 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 a_27_297# C1 a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 a_861_47# A2 a_1059_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 a_109_47# C1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 a_277_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
X0 a_376_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VPWR A1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_109_47# A2 a_194_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_194_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VGND A3 a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR A3 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_109_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_109_297# B1 a_376_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
X0 a_109_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 Y C1 a_641_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_277_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_109_297# B1 a_641_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_277_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_641_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VPWR A1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_27_47# A2 a_277_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 Y A1 a_277_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_641_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 VPWR A3 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 a_109_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
X0 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_109_297# B1 a_1139_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 Y A1 a_445_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_27_47# A2 a_445_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_27_47# A2 a_445_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_1139_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 Y A1 a_445_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VPWR A1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_109_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_1139_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_109_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 Y C1 a_1139_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 Y C1 a_1139_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 VPWR A1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_445_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 a_1139_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 VPWR A3 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X29 VPWR A3 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X30 a_1139_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X31 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X32 a_109_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X33 a_445_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X34 a_445_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X35 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X36 a_109_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X37 a_109_297# B1 a_1139_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X38 a_445_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X39 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
X0 VGND D1 a_85_193# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 X a_85_193# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_516_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_414_297# B1 a_516_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_660_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VPWR A2 a_516_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_85_193# C1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 X a_85_193# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND B1 a_85_193# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_85_193# A1 a_660_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_85_193# D1 a_334_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_334_297# C1 a_414_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
X0 a_86_235# A1 a_715_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VGND a_86_235# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_715_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VGND D1 a_86_235# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_86_235# C1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VPWR a_86_235# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VGND B1 a_86_235# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VPWR A2 a_607_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 X a_86_235# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_607_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_499_297# B1 a_607_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_86_235# D1 a_427_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_427_297# C1 a_499_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 X a_86_235# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
X0 a_477_297# B1 a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_44_47# A1 a_770_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_44_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VGND a_44_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_44_47# D1 a_30_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 X a_44_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR A1 a_477_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VPWR a_44_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_285_297# B1 a_477_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VGND B1 a_44_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_770_47# A1 a_44_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_30_297# D1 a_44_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VGND D1 a_44_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VGND C1 a_44_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VGND A2 a_770_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_30_297# C1 a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 a_477_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 VPWR a_44_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 VGND a_44_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 VPWR A2 a_477_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 X a_44_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 X a_44_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 a_44_47# C1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 a_770_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 a_285_297# C1 a_30_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 X a_44_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 a_477_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 a_44_47# D1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a2111oi_0 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
X0 VPWR A2 a_313_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X1 Y A1 a_427_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_313_369# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X3 a_241_369# B1 a_313_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X4 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 Y D1 a_169_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X6 VGND D1 Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_169_369# C1 a_241_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 a_427_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
X0 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_316_297# B1 a_420_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 Y A1 a_568_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 Y D1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_420_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_568_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VGND D1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_217_297# C1 a_316_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VPWR A2 a_420_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
X0 VGND D1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_467_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_923_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_467_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 Y D1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_28_297# C1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_28_297# B1 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 Y D1 a_287_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_115_297# D1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_467_297# B1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VPWR A1 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_287_297# C1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 VPWR A2 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 VGND A2 a_923_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 a_684_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 Y A1 a_684_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
X0 VPWR A1 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_821_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 Y D1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_821_297# B1 a_455_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_28_297# D1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_455_297# B1 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_821_297# B1 a_455_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_1205_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 Y D1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_28_297# C1 a_455_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_28_297# D1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VGND D1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_455_297# B1 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 a_821_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 a_821_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 Y D1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 a_28_297# C1 a_455_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 a_455_297# C1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 VGND D1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 Y A1 a_1205_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 a_1205_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 a_1205_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 VPWR A2 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 a_821_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 VGND A2 a_1205_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 VPWR A1 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X32 a_455_297# C1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X33 Y D1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X34 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X35 a_1205_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X36 Y A1 a_1205_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X37 VGND A2 a_1205_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X38 VPWR A2 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X39 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__and2_0 A B VGND VNB VPB VPWR X
X0 a_40_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_123_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_40_47# A a_123_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VGND a_40_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VPWR A a_40_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 VPWR a_40_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
X0 VGND a_59_75# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VPWR A a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_59_75# A a_145_75# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_59_75# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_145_75# B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VPWR a_59_75# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
X0 VPWR a_61_75# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VPWR A a_61_75# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_147_75# B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_61_75# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 VGND a_61_75# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 X a_61_75# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_61_75# A a_147_75# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 X a_61_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
X0 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_110_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_27_47# A a_110_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
X0 a_207_413# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 VPWR a_207_413# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VGND a_207_413# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_207_413# a_27_413# a_297_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_27_413# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 VPWR a_27_413# a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 VGND A_N a_27_413# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_297_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
X0 VPWR a_27_413# a_212_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_212_413# a_27_413# a_297_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VPWR a_212_413# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VGND a_212_413# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 X a_212_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_212_413# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_27_413# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VGND A_N a_27_413# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_297_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 X a_212_413# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
X0 VPWR A_N a_33_199# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VGND A_N a_33_199# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_27_47# a_33_199# a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VPWR a_33_199# a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_109_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
X0 a_181_47# C VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_109_47# B a_181_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_27_47# A a_109_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
X0 X a_29_311# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 X a_29_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_184_53# C VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_29_311# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 VGND a_29_311# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_112_53# B a_184_53# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_29_311# A a_112_53# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VPWR a_29_311# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VPWR B a_29_311# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 a_29_311# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
X0 a_185_47# B a_294_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 X a_94_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VPWR B a_94_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_94_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_94_47# A a_185_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_94_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VGND a_94_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 X a_94_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VPWR a_94_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_294_47# C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 X a_94_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VGND a_94_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 X a_94_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VPWR a_94_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
X0 a_209_311# a_109_93# a_296_53# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VGND a_209_311# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VGND A_N a_109_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VPWR a_209_311# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VPWR A_N a_109_93# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_368_53# C VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VPWR B a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_209_311# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_296_53# B a_368_53# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_209_311# a_109_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
X0 a_373_53# C VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 X a_215_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_215_311# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_215_311# a_109_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 VPWR a_215_311# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_301_53# B a_373_53# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VPWR B a_215_311# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VGND A_N a_109_53# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_215_311# a_109_53# a_301_53# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 X a_215_311# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VGND a_215_311# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VPWR A_N a_109_53# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
X0 X a_56_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_257_47# C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VGND a_56_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR B a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 X a_56_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 X a_56_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VPWR A_N a_98_199# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_56_297# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND a_56_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_56_297# a_98_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_56_297# a_98_199# a_152_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VGND A_N a_98_199# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VPWR a_56_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 X a_56_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_152_47# B a_257_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 VPWR a_56_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
X0 a_197_47# C a_303_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_303_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_27_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_109_47# B a_197_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 a_27_47# A a_109_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
X0 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_109_47# B a_198_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_27_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 a_27_47# A a_109_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_304_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_198_47# C a_304_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
X0 a_27_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_285_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_109_47# B a_188_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_27_47# A a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_188_47# C a_285_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
X0 VPWR a_193_413# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_193_413# a_27_47# a_297_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_193_413# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 VPWR C a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_369_47# C a_469_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_27_47# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_193_413# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VGND a_193_413# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VPWR a_27_47# a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 a_27_47# A_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_297_47# B a_369_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_469_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
X0 VPWR a_193_413# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_193_413# a_27_413# a_297_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_193_413# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 VPWR C a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 VGND a_193_413# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_369_47# C a_469_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_27_413# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_193_413# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 VPWR a_27_413# a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 X a_193_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_469_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VGND A_N a_27_413# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_297_47# B a_369_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 X a_193_413# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
X0 a_174_21# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 X a_174_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VGND a_174_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_815_47# a_27_47# a_174_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_617_47# C a_701_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VPWR D a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 X a_174_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 X a_174_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_27_47# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 X a_174_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_174_21# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 VPWR a_174_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VGND a_174_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VPWR a_174_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_27_47# A_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_701_47# B a_815_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VGND D a_617_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 VPWR B a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
X0 VPWR B_N a_223_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_343_93# a_223_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 VGND B_N a_223_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VPWR C a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_515_93# C a_615_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_27_47# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 VPWR a_343_93# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_343_93# a_27_47# a_429_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_429_93# a_223_47# a_515_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_343_93# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_27_47# A_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_615_93# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VPWR a_27_47# a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X13 VGND a_343_93# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
X0 X a_174_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_174_21# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 VGND a_174_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_174_21# a_27_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VPWR B_N a_505_280# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_548_47# C a_639_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VPWR C a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_174_21# a_505_280# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_639_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VPWR a_27_47# a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 X a_174_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_27_47# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X12 VPWR a_174_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_27_47# A_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_476_47# a_505_280# a_548_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 VGND B_N a_505_280# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
X0 VPWR a_27_47# a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_174_21# a_832_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 X a_174_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_556_47# C a_652_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VPWR A_N a_832_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 VGND a_174_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VGND D a_556_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_766_47# a_832_21# a_174_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_652_47# a_27_47# a_766_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 X a_174_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 X a_174_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_27_47# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X12 X a_174_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VPWR a_174_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 VGND a_174_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 VPWR a_174_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 a_27_47# B_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 VGND A_N a_832_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 VPWR D a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_174_21# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
X0 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X1 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
X2 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X3 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
X0 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_161_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VPWR A a_161_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_161_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VGND A a_161_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
X0 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X28 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X29 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X30 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__buf_16 A VGND VNB VPB VPWR X
X0 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X32 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X33 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X34 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X35 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X36 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X37 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X38 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X39 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X40 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X41 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X42 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X43 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__bufbuf_8 A VGND VNB VPB VPWR X
X0 X a_318_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 X a_318_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 X a_318_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VGND a_318_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 X a_318_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND a_318_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR a_318_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 X a_318_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VPWR a_318_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_318_47# a_206_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 X a_318_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VGND a_27_47# a_206_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VGND a_206_47# a_318_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_318_47# a_206_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 X a_318_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_318_47# a_206_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 VPWR a_27_47# a_206_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 VGND a_318_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X20 VPWR a_206_47# a_318_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 VPWR a_318_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 VGND a_318_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 VPWR a_318_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X24 X a_318_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 a_318_47# a_206_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__bufbuf_16 A VGND VNB VPB VPWR X
X0 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VGND a_215_47# a_549_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_549_47# a_215_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_215_47# a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_549_47# a_215_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VPWR a_215_47# a_549_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_215_47# a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 a_215_47# a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_549_47# a_215_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X24 VPWR a_109_47# a_215_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 VGND a_215_47# a_549_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X29 VGND a_215_47# a_549_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X32 a_549_47# a_215_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X33 a_215_47# a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X34 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X35 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X36 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X37 VPWR a_215_47# a_549_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X38 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X39 VPWR a_215_47# a_549_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X40 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X41 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X42 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X43 VGND a_109_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X44 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X45 a_549_47# a_215_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X46 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X47 a_549_47# a_215_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X48 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X49 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X50 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X51 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__bufinv_8 A VGND VNB VPB VPWR Y
X0 VGND a_215_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VGND a_215_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 Y a_215_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_215_47# a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 Y a_215_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VPWR a_215_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_215_47# a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_215_47# a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 Y a_215_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 Y a_215_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VPWR a_109_47# a_215_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 VGND a_215_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VPWR a_215_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VGND a_215_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 Y a_215_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_215_47# a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VPWR a_215_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 VPWR a_215_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 VGND a_109_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 Y a_215_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 Y a_215_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 Y a_215_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
X0 VPWR a_361_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 Y a_361_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_361_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_361_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VGND a_361_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VGND a_361_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 Y a_361_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VPWR a_27_47# a_361_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 Y a_361_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VGND a_361_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VPWR a_27_47# a_361_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 VGND a_27_47# a_361_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VPWR a_361_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 Y a_361_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VPWR a_361_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 Y a_361_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_361_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 VPWR a_361_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 a_361_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 Y a_361_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 VGND a_27_47# a_361_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 Y a_361_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 VGND a_361_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 VGND a_361_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 Y a_361_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 Y a_361_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 VGND a_361_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 Y a_361_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 VPWR a_361_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X29 a_361_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 VGND a_361_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X32 VGND a_361_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X33 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X34 Y a_361_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X35 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X36 Y a_361_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X37 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X38 Y a_361_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X39 VPWR a_361_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X40 Y a_361_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X41 Y a_361_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X42 a_361_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X43 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X44 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X45 VPWR a_361_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X46 VPWR a_361_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X47 VGND a_27_47# a_361_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X48 VPWR a_27_47# a_361_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X49 Y a_361_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
X0 VGND A a_75_212# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X1 X a_75_212# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
X2 X a_75_212# VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X3 VPWR A a_75_212# VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
X0 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
X0 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
X0 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X29 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X30 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X32 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X33 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X34 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X36 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X37 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X38 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X39 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__clkdlybuf4s15_1 A VGND VNB VPB VPWR X
X0 a_394_47# a_282_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=150000u
X1 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VPWR a_27_47# a_282_47# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=150000u
X3 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VGND a_394_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VPWR a_394_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VGND a_27_47# a_282_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_394_47# a_282_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__clkdlybuf4s15_2 A VGND VNB VPB VPWR X
X0 a_362_333# a_228_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VPWR a_27_47# a_228_47# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=150000u
X3 VPWR a_362_333# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VGND a_27_47# a_228_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_362_333# a_228_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=150000u
X6 X a_362_333# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VGND a_362_333# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 X a_362_333# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__clkdlybuf4s18_1 A VGND VNB VPB VPWR X
X0 a_394_47# a_282_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X1 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VGND a_394_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VPWR a_394_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VPWR a_27_47# a_282_47# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X6 VGND a_27_47# a_282_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=180000u
X7 a_394_47# a_282_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=180000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__clkdlybuf4s18_2 A VGND VNB VPB VPWR X
X0 a_334_47# a_227_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X1 VPWR a_27_47# a_227_47# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X2 VPWR a_334_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 X a_334_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_334_47# a_227_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=180000u
X6 VGND a_27_47# a_227_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=180000u
X7 VGND a_334_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 X a_334_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
X0 a_355_47# a_244_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=250000u
X1 VPWR a_27_47# a_244_47# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=250000u
X2 VPWR a_355_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_355_47# a_244_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=250000u
X5 VGND a_27_47# a_244_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=250000u
X6 VGND a_355_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__clkdlybuf4s25_2 A VGND VNB VPB VPWR X
X0 VPWR a_331_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 X a_331_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 X a_331_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VPWR a_27_47# a_225_47# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=250000u
X6 a_331_47# a_225_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=250000u
X7 VGND a_331_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_331_47# a_225_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=250000u
X9 VGND a_27_47# a_225_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=250000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VNB VPB VPWR X
X0 a_390_47# a_283_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=500000u
X1 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VPWR a_27_47# a_283_47# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=500000u
X3 VGND a_27_47# a_283_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=500000u
X4 VPWR a_390_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND a_390_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_390_47# a_283_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=500000u
X7 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__clkdlybuf4s50_2 A VGND VNB VPB VPWR X
X0 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VPWR a_27_47# a_283_47# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=500000u
X2 X a_390_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VGND a_27_47# a_283_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=500000u
X4 a_390_47# a_283_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=500000u
X5 X a_390_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VPWR a_390_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VGND a_390_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_390_47# a_283_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=500000u
X9 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__clkinv_16 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X28 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X30 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X31 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X32 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X33 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X35 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X36 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X37 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X38 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X39 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__clkinvlp_2 A VGND VNB VPB VPWR Y
X0 a_150_67# A Y VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X3 VGND A a_150_67# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 a_110_47# A Y VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X2 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X4 Y A a_268_47# VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X6 a_268_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X7 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
R0 VGND LO sky130_fd_pr__res_generic_po w=480000u l=45000u
R1 HI VPWR sky130_fd_pr__res_generic_po w=480000u l=45000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=870000u l=590000u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=590000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=870000u l=1.05e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=1.05e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=870000u l=1.97e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=1.97e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=870000u l=2.89e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=2.89e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=870000u l=4.73e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=4.73e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dfbbn_1 CLK_N D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
X0 VGND a_647_21# a_1159_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X1 a_2136_47# a_1415_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 a_647_21# a_941_21# a_791_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X3 a_1256_413# a_27_47# a_1340_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_473_413# a_27_47# a_581_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X5 a_381_47# a_193_47# a_473_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X6 VPWR D a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VPWR SET_B a_647_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 VPWR a_647_21# a_1112_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X9 a_581_47# a_647_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_1159_47# a_27_47# a_1256_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X11 a_941_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X12 a_1363_47# a_1415_315# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 VGND SET_B a_791_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_891_329# a_941_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X15 VPWR SET_B a_1415_315# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X16 a_2136_47# a_1415_315# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_791_47# a_473_413# a_647_21# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X18 a_557_413# a_647_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X19 a_647_21# a_473_413# a_891_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X20 a_1415_315# a_1256_413# a_1672_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X21 a_1672_329# a_941_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X22 VGND a_2136_47# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 a_1340_413# a_1415_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X24 VGND a_1415_315# Q_N VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 a_473_413# a_193_47# a_557_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X26 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 VPWR a_2136_47# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X28 a_27_47# CLK_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 a_27_47# CLK_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X30 a_381_47# a_27_47# a_473_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X31 a_1415_315# a_941_21# a_1555_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X32 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X33 VGND D a_381_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 VGND SET_B a_1555_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 a_1256_413# a_193_47# a_1363_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X36 a_1112_329# a_193_47# a_1256_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X37 a_1555_47# a_1256_413# a_1415_315# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X38 a_941_21# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X39 VPWR a_1415_315# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dfbbn_2 CLK_N D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
X0 a_944_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X1 Q_N a_1431_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_1257_47# a_193_47# a_1366_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X3 a_2236_47# a_1431_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_1115_329# a_193_47# a_1257_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 Q a_2236_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_476_47# a_193_47# a_560_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_584_47# a_650_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_650_21# a_944_21# a_790_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X9 a_1366_47# a_1431_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VGND a_1431_21# Q_N VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VGND a_2236_47# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_381_47# a_193_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X13 a_1431_21# a_944_21# a_1547_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X14 VPWR D a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 a_1257_47# a_27_47# a_1343_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X16 a_2236_47# a_1431_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X17 a_1162_47# a_27_47# a_1257_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X18 a_476_47# a_27_47# a_584_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X19 Q_N a_1431_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_894_329# a_944_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X21 a_790_47# a_476_47# a_650_21# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X22 VPWR a_1431_21# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 a_1547_47# a_1257_47# a_1431_21# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X24 VPWR SET_B a_650_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X25 VPWR a_650_21# a_1115_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X26 VGND SET_B a_1547_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 VPWR SET_B a_1431_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X28 VGND SET_B a_790_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 a_650_21# a_476_47# a_894_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X30 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 a_27_47# CLK_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X32 a_27_47# CLK_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X33 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X34 VGND D a_381_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 Q a_2236_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X36 a_560_413# a_650_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X37 VGND a_650_21# a_1162_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X38 a_1343_413# a_1431_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X39 a_1431_21# a_1257_47# a_1665_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X40 a_1665_329# a_944_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X41 a_944_21# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X42 a_381_47# a_27_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X43 VPWR a_2236_47# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dfbbp_1 CLK D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
X0 a_1364_47# a_1429_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_2136_47# a_1429_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 VGND SET_B a_1545_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_788_47# a_474_413# a_648_21# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X4 a_1255_47# a_193_47# a_1341_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_381_47# a_27_47# a_474_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X6 VPWR D a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VPWR SET_B a_648_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 VPWR a_648_21# a_1113_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X9 a_942_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X10 a_2136_47# a_1429_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_892_329# a_942_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X12 VPWR SET_B a_1429_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X13 VGND SET_B a_788_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 VGND a_648_21# a_1160_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X15 a_558_413# a_648_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X16 a_648_21# a_474_413# a_892_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X17 a_1341_413# a_1429_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X18 VGND a_2136_47# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 VGND a_1429_21# Q_N VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_1255_47# a_27_47# a_1364_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X21 a_474_413# a_27_47# a_558_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X22 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 VPWR a_2136_47# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X24 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 a_648_21# a_942_21# a_788_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X26 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X27 a_1429_21# a_1255_47# a_1663_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X28 a_1663_329# a_942_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X29 a_1429_21# a_942_21# a_1545_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X30 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X31 a_381_47# a_193_47# a_474_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X32 VGND D a_381_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X33 a_1160_47# a_193_47# a_1255_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X34 a_474_413# a_193_47# a_582_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X35 a_1545_47# a_1255_47# a_1429_21# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X36 a_942_21# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X37 a_1113_329# a_27_47# a_1255_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X38 a_582_47# a_648_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X39 VPWR a_1429_21# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dfrbp_1 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
X0 a_1270_413# a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 VPWR a_543_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X2 VGND a_543_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X3 VPWR a_1847_47# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VGND D a_448_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_1108_47# a_193_47# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_1217_47# a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_448_47# a_27_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X8 a_1847_47# a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_448_47# a_193_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 a_543_47# a_193_47# a_639_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X12 a_1108_47# a_27_47# a_1217_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X13 a_1462_47# a_1108_47# a_1283_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_543_47# a_27_47# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X16 a_805_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_761_289# a_193_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X18 VPWR RESET_B a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X19 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X22 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X23 a_1283_21# a_1108_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X24 a_1847_47# a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X25 VGND RESET_B a_1462_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 VPWR D a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X27 a_651_413# a_761_289# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X28 a_761_289# a_27_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X29 VGND a_1847_47# Q_N VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 VPWR RESET_B a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X31 a_639_47# a_761_289# a_805_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dfrbp_2 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
X0 a_1270_413# a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 Q_N a_1659_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR a_543_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X4 VGND a_543_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X5 VGND D a_448_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_1108_47# a_193_47# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VPWR a_1659_47# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_1217_47# a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_448_47# a_27_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X10 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_448_47# a_193_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X13 a_543_47# a_193_47# a_639_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X14 a_1108_47# a_27_47# a_1217_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X15 a_1462_47# a_1108_47# a_1283_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_1659_47# a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X17 a_1659_47# a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_543_47# a_27_47# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X19 a_805_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_761_289# a_193_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X21 VPWR RESET_B a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X22 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 VGND a_1659_47# Q_N VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X26 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X27 a_1283_21# a_1108_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X28 VGND RESET_B a_1462_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 VPWR D a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X30 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X31 a_651_413# a_761_289# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X32 a_761_289# a_27_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X33 VPWR RESET_B a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X34 a_639_47# a_761_289# a_805_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 Q_N a_1659_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
X0 a_1270_413# a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 VPWR a_543_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X2 VGND a_543_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X3 VGND D a_448_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_1108_47# a_27_47# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_1217_47# a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_448_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X8 a_448_47# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 a_543_47# a_27_47# a_639_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X10 a_1108_47# a_193_47# a_1217_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X11 a_1462_47# a_1108_47# a_1283_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_543_47# a_193_47# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X13 a_805_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_761_289# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X15 VPWR RESET_B a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X16 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_27_47# CLK_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_27_47# CLK_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X19 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X21 a_1283_21# a_1108_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X22 VGND RESET_B a_1462_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 VPWR D a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X24 a_651_413# a_761_289# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X25 a_761_289# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X26 VPWR RESET_B a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X27 a_639_47# a_761_289# a_805_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
X0 a_1270_413# a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 VPWR a_543_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X2 VGND a_543_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X3 VGND D a_448_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_1108_47# a_193_47# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_1217_47# a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_448_47# a_27_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X8 a_448_47# a_193_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 a_543_47# a_193_47# a_639_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X10 a_1108_47# a_27_47# a_1217_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X11 a_1462_47# a_1108_47# a_1283_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_543_47# a_27_47# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X13 a_805_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_761_289# a_193_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X15 VPWR RESET_B a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X16 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X19 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X21 a_1283_21# a_1108_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X22 VGND RESET_B a_1462_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 VPWR D a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X24 a_651_413# a_761_289# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X25 a_761_289# a_27_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X26 VPWR RESET_B a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X27 a_639_47# a_761_289# a_805_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
X0 a_1270_413# a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VPWR a_543_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X3 VGND a_543_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X4 VGND D a_448_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_1108_47# a_193_47# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_1217_47# a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_448_47# a_27_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X9 a_448_47# a_193_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_543_47# a_193_47# a_639_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X11 a_1108_47# a_27_47# a_1217_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X12 a_1462_47# a_1108_47# a_1283_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_543_47# a_27_47# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X14 a_805_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 a_761_289# a_193_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X17 VPWR RESET_B a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X18 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X21 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X23 a_1283_21# a_1108_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X24 VGND RESET_B a_1462_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 VPWR D a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X26 a_651_413# a_761_289# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X27 a_761_289# a_27_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X28 VPWR RESET_B a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X29 a_639_47# a_761_289# a_805_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
X0 a_1270_413# a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 VPWR a_543_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X2 VGND a_543_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X3 VGND D a_448_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_1108_47# a_193_47# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_1217_47# a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_448_47# a_27_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X8 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_448_47# a_193_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_543_47# a_193_47# a_639_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X11 a_1108_47# a_27_47# a_1217_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X12 a_1462_47# a_1108_47# a_1283_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_543_47# a_27_47# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X16 a_805_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_761_289# a_193_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X20 VPWR RESET_B a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X21 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X25 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X26 a_1283_21# a_1108_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X27 VGND RESET_B a_1462_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 VPWR D a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X29 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 a_651_413# a_761_289# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X31 a_761_289# a_27_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X32 VPWR RESET_B a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X33 a_639_47# a_761_289# a_805_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dfsbp_1 CLK D SET_B VGND VNB VPB VPWR Q Q_N
X0 a_562_413# a_652_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_956_413# a_27_47# a_1028_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_381_47# a_193_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 VPWR a_1028_413# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_1028_413# a_193_47# a_1136_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_1028_413# a_27_47# a_1224_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_1786_47# a_1028_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 a_476_47# a_27_47# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_381_47# a_27_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X9 VGND a_476_47# a_1056_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_1028_413# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 a_1056_47# a_193_47# a_1028_413# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VGND a_1028_413# a_1178_261# VNB sky130_fd_pr__nfet_01v8 w=540000u l=150000u
X13 VPWR a_1786_47# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_1296_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 VGND a_1028_413# Q_N VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VPWR SET_B a_652_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X17 a_796_47# a_476_47# a_652_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 VPWR a_476_47# a_956_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X19 a_586_47# a_652_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 VPWR D a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X21 VPWR a_1028_413# a_1178_261# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X22 a_652_21# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X23 a_1136_413# a_1178_261# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X24 a_476_47# a_193_47# a_586_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X25 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X28 a_1224_47# a_1178_261# a_1296_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 a_1786_47# a_1028_413# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X30 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X31 VGND D a_381_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X32 VGND SET_B a_796_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X33 VGND a_1786_47# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dfsbp_2 CLK D SET_B VGND VNB VPB VPWR Q Q_N
X0 a_562_413# a_652_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_956_413# a_27_47# a_1028_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_381_47# a_193_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 VPWR a_1028_413# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_1028_413# a_193_47# a_1136_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_1028_413# a_27_47# a_1224_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_476_47# a_27_47# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_381_47# a_27_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X8 VGND a_476_47# a_1056_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_1028_413# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 VPWR a_1870_47# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_1056_47# a_193_47# a_1028_413# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VGND a_1028_413# a_1178_261# VNB sky130_fd_pr__nfet_01v8 w=540000u l=150000u
X13 Q_N a_1028_413# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_1296_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 VGND a_1028_413# Q_N VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_1870_47# a_1028_413# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 VPWR SET_B a_652_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X18 a_796_47# a_476_47# a_652_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 VPWR a_476_47# a_956_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X20 a_1870_47# a_1028_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 a_586_47# a_652_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 VPWR D a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X23 VPWR a_1028_413# a_1178_261# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X24 a_652_21# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X25 a_1136_413# a_1178_261# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X26 a_476_47# a_193_47# a_586_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X27 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X30 VGND a_1870_47# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 a_1224_47# a_1178_261# a_1296_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X32 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X33 VGND D a_381_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X34 VGND SET_B a_796_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 Q a_1870_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X36 Q a_1870_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X37 Q_N a_1028_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
X0 a_562_413# a_652_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_1296_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_381_47# a_193_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_1602_47# a_1032_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X4 a_1140_413# a_1182_261# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_1032_413# a_27_47# a_1224_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VGND a_1032_413# a_1182_261# VNB sky130_fd_pr__nfet_01v8 w=540000u l=150000u
X7 a_476_47# a_27_47# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_381_47# a_27_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X9 VGND a_476_47# a_1056_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_1602_47# a_1032_413# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_1056_47# a_193_47# a_1032_413# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VPWR SET_B a_652_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X13 a_796_47# a_476_47# a_652_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 VPWR a_476_47# a_956_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 a_586_47# a_652_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 VPWR D a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X17 a_652_21# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X18 a_1032_413# a_193_47# a_1140_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X19 VGND a_1602_47# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_476_47# a_193_47# a_586_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X21 a_1032_413# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X22 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_956_413# a_27_47# a_1032_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X24 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X26 VPWR a_1032_413# a_1182_261# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X27 a_1224_47# a_1182_261# a_1296_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X29 VGND D a_381_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X30 VGND SET_B a_796_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 VPWR a_1602_47# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
X0 a_562_413# a_652_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_956_413# a_27_47# a_1028_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_1300_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_381_47# a_193_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 VGND a_1602_47# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_1028_413# a_193_47# a_1136_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 VPWR a_1602_47# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VGND a_1028_413# a_1178_261# VNB sky130_fd_pr__nfet_01v8 w=540000u l=150000u
X8 a_476_47# a_27_47# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 a_381_47# a_27_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X10 VGND a_476_47# a_1056_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_1028_413# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X12 a_1602_47# a_1028_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_1602_47# a_1028_413# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 Q a_1602_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_1056_47# a_193_47# a_1028_413# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_1228_47# a_1178_261# a_1300_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 VPWR SET_B a_652_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X18 a_796_47# a_476_47# a_652_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 VPWR a_476_47# a_956_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X20 VPWR a_1028_413# a_1178_261# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X21 a_586_47# a_652_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 VPWR D a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X23 a_652_21# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X24 a_1136_413# a_1178_261# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X25 a_476_47# a_193_47# a_586_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X26 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X29 Q a_1602_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X31 VGND D a_381_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X32 VGND SET_B a_796_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X33 a_1028_413# a_27_47# a_1228_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
X0 a_562_413# a_652_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_956_413# a_27_47# a_1028_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_381_47# a_193_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_1028_413# a_193_47# a_1136_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_1028_413# a_27_47# a_1224_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 Q a_1598_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VPWR a_1598_47# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_476_47# a_27_47# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_381_47# a_27_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X9 VGND a_476_47# a_1056_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_1028_413# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 a_1056_47# a_193_47# a_1028_413# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VGND a_1028_413# a_1178_261# VNB sky130_fd_pr__nfet_01v8 w=540000u l=150000u
X13 VGND a_1598_47# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_1296_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_1598_47# a_1028_413# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 VPWR SET_B a_652_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X17 a_796_47# a_476_47# a_652_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 VPWR a_476_47# a_956_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X19 a_586_47# a_652_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 VPWR D a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X21 VPWR a_1028_413# a_1178_261# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X22 a_652_21# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X23 a_1136_413# a_1178_261# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X24 Q a_1598_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 Q a_1598_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 a_476_47# a_193_47# a_586_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X27 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 Q a_1598_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X30 VGND a_1598_47# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X32 VPWR a_1598_47# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X33 VPWR a_1598_47# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X34 a_1224_47# a_1178_261# a_1296_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X36 VGND D a_381_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X37 VGND SET_B a_796_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X38 VGND a_1598_47# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X39 a_1598_47# a_1028_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dfxbp_1 CLK D VGND VNB VPB VPWR Q Q_N
X0 a_1490_369# a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X1 a_891_413# a_193_47# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_466_413# a_27_47# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_634_159# a_27_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 VGND a_1490_369# Q_N VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_381_47# a_193_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 VPWR D a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VPWR a_466_413# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt w=750000u l=150000u
X8 VGND a_466_413# a_634_159# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X9 a_1017_47# a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_561_413# a_634_159# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 a_891_413# a_27_47# a_1017_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X12 VPWR a_1059_315# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_634_159# a_193_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X14 a_592_47# a_634_159# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 VGND a_1059_315# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_466_413# a_193_47# a_592_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X17 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_381_47# a_27_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X19 a_1059_315# a_891_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X22 a_1059_315# a_891_413# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 a_1490_369# a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X25 VGND D a_381_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 a_975_413# a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X27 VPWR a_1490_369# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dfxbp_2 CLK D VGND VNB VPB VPWR Q Q_N
X0 a_891_413# a_193_47# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 VGND a_1589_47# Q_N VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_466_413# a_27_47# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_634_159# a_27_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_1589_47# a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 VPWR a_1589_47# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_381_47# a_193_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VPWR D a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 VPWR a_466_413# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt w=750000u l=150000u
X9 VGND a_466_413# a_634_159# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X10 a_1017_47# a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 Q_N a_1589_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_1589_47# a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_561_413# a_634_159# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X16 a_891_413# a_27_47# a_1017_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X17 VPWR a_1059_315# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 a_634_159# a_193_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X19 a_592_47# a_634_159# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 VGND a_1059_315# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 a_466_413# a_193_47# a_592_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X22 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_381_47# a_27_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X24 a_1059_315# a_891_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X27 a_1059_315# a_891_413# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 Q_N a_1589_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X30 VGND D a_381_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 a_975_413# a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
X0 a_891_413# a_193_47# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_1059_315# a_891_413# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_466_413# a_27_47# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_634_159# a_27_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_381_47# a_193_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 VPWR D a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 VPWR a_466_413# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt w=750000u l=150000u
X7 VGND a_466_413# a_634_159# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X8 a_1017_47# a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_1059_315# a_891_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_561_413# a_634_159# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 VPWR a_1059_315# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_891_413# a_27_47# a_1017_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X13 a_634_159# a_193_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X14 a_592_47# a_634_159# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_466_413# a_193_47# a_592_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X16 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_381_47# a_27_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X18 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X20 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X21 VGND D a_381_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_975_413# a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X23 VGND a_1059_315# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
X0 a_891_413# a_193_47# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_1059_315# a_891_413# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_466_413# a_27_47# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_634_159# a_27_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_381_47# a_193_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 VPWR D a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 VPWR a_466_413# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt w=750000u l=150000u
X7 VGND a_466_413# a_634_159# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X8 a_1017_47# a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_1059_315# a_891_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_561_413# a_634_159# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X12 VPWR a_1059_315# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_891_413# a_27_47# a_1017_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X14 a_634_159# a_193_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X15 a_592_47# a_634_159# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_466_413# a_193_47# a_592_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X17 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_381_47# a_27_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X19 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X21 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X23 VGND D a_381_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 a_975_413# a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X25 VGND a_1059_315# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
X0 a_891_413# a_193_47# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_1062_300# a_891_413# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 Q a_1062_300# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_475_413# a_193_47# a_572_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X4 a_1062_300# a_891_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VPWR a_1062_300# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_634_183# a_27_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 Q a_1062_300# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND a_1062_300# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_381_47# a_27_47# a_475_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X10 VPWR D a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 VPWR a_475_413# a_634_183# VPB sky130_fd_pr__pfet_01v8_hvt w=750000u l=150000u
X12 VPWR a_1062_300# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_572_47# a_634_183# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_975_413# a_1062_300# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 a_1020_47# a_1062_300# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_891_413# a_27_47# a_1020_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X17 VGND a_475_413# a_634_183# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X18 a_475_413# a_27_47# a_568_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X19 a_568_413# a_634_183# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X20 Q a_1062_300# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X24 VGND a_1062_300# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X26 VGND D a_381_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 a_634_183# a_193_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X28 a_381_47# a_193_47# a_475_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X29 Q a_1062_300# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=5.36e+06u area=4.347e+11p
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dlclkp_1 CLK GATE VGND VNB VPB VPWR GCLK
X0 a_957_369# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X1 VGND a_957_369# GCLK VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_642_307# a_476_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_476_413# a_27_47# a_600_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_600_413# a_642_307# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 VGND GATE a_396_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VPWR GATE a_381_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 a_476_413# a_193_47# a_651_47# VNB sky130_fd_pr__nfet_01v8 w=390000u l=150000u
X8 a_957_369# a_642_307# a_1042_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VPWR a_642_307# a_957_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X10 a_396_119# a_27_47# a_476_413# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_1042_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X15 a_651_47# a_642_307# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X17 VGND a_476_413# a_642_307# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 VPWR a_957_369# GCLK VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_381_369# a_193_47# a_476_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dlclkp_2 CLK GATE VGND VNB VPB VPWR GCLK
X0 a_381_369# a_193_47# a_477_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_957_369# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 VGND GATE a_397_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_643_307# a_477_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VGND a_957_369# GCLK VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 GCLK a_957_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_477_413# a_193_47# a_652_47# VNB sky130_fd_pr__nfet_01v8 w=390000u l=150000u
X7 VGND a_477_413# a_643_307# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_477_413# a_27_47# a_601_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 a_601_413# a_643_307# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 VPWR GATE a_381_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X11 a_397_119# a_27_47# a_477_413# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_652_47# a_643_307# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 VPWR a_643_307# a_957_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X14 GCLK a_957_369# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X19 a_957_369# a_643_307# a_1041_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 VPWR a_957_369# GCLK VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 a_1041_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dlclkp_4 CLK GATE VGND VNB VPB VPWR GCLK
X0 a_381_369# a_193_47# a_477_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_1046_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VGND a_953_297# GCLK VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_477_413# a_193_47# a_575_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X4 VPWR GATE a_381_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 a_575_47# a_627_153# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VGND a_953_297# GCLK VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_627_153# a_477_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_953_297# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_953_297# a_627_153# a_1046_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 GCLK a_953_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VPWR a_953_297# GCLK VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_381_47# a_27_47# a_477_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X13 VPWR a_627_153# a_953_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_627_153# a_477_413# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 GCLK a_953_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 GCLK a_953_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X21 VGND GATE a_381_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_477_413# a_27_47# a_585_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X23 a_585_413# a_627_153# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X24 VPWR a_953_297# GCLK VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 GCLK a_953_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dlrbn_1 D GATE_N RESET_B VGND VNB VPB VPWR Q Q_N
X0 a_561_413# a_27_47# a_682_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_682_413# a_724_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_724_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_561_413# a_193_47# a_659_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X4 VGND a_724_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VPWR a_299_47# a_465_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X6 a_465_369# a_193_47# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_942_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_659_47# a_724_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_1308_47# a_724_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_299_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X11 a_724_21# a_561_413# a_942_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VPWR a_724_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VGND a_1308_47# Q_N VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VGND a_299_47# a_465_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_27_47# GATE_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_27_47# GATE_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 VPWR a_561_413# a_724_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_465_47# a_27_47# a_561_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X20 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X21 a_299_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 VPWR a_1308_47# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 a_1308_47# a_724_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dlrbn_2 D GATE_N RESET_B VGND VNB VPB VPWR Q Q_N
X0 a_561_413# a_27_47# a_682_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_682_413# a_724_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 VPWR a_724_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_561_413# a_193_47# a_659_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X4 VPWR a_299_47# a_465_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 a_465_369# a_193_47# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_724_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_659_47# a_724_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_1313_47# a_724_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 Q a_724_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_299_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X11 Q_N a_1313_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_724_21# a_561_413# a_942_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VPWR a_1313_47# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 Q_N a_1313_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_942_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VGND a_299_47# a_465_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 Q a_724_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_27_47# GATE_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_27_47# GATE_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X21 VPWR a_561_413# a_724_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 a_465_47# a_27_47# a_561_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X23 a_1313_47# a_724_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X25 a_299_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 VGND a_724_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 VGND a_1313_47# Q_N VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dlrbp_1 D GATE RESET_B VGND VNB VPB VPWR Q Q_N
X0 a_560_47# a_193_47# a_645_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_645_413# a_711_307# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 VGND a_711_307# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR a_299_47# a_465_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X4 a_465_369# a_27_47# a_560_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_1308_47# a_711_307# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_299_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 VPWR a_560_47# a_711_307# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_560_47# a_27_47# a_658_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X9 a_941_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_658_47# a_711_307# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VPWR a_711_307# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_711_307# a_560_47# a_941_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VGND a_1308_47# Q_N VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VGND a_299_47# a_465_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_27_47# GATE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_27_47# GATE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X19 a_299_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_711_307# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 a_465_47# a_193_47# a_560_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X22 VPWR a_1308_47# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 a_1308_47# a_711_307# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dlrbp_2 D GATE RESET_B VGND VNB VPB VPWR Q Q_N
X0 a_561_413# a_193_47# a_645_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 VGND a_1316_47# Q_N VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_645_413# a_711_307# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_561_413# a_27_47# a_659_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X4 a_942_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VGND a_711_307# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR a_299_47# a_465_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 a_465_369# a_27_47# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_659_47# a_711_307# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_711_307# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 Q a_711_307# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_299_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X12 a_711_307# a_561_413# a_942_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_1316_47# a_711_307# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X14 Q_N a_1316_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 VPWR a_1316_47# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 Q a_711_307# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 VGND a_299_47# a_465_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_27_47# GATE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_27_47# GATE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X21 VPWR a_561_413# a_711_307# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 a_465_47# a_193_47# a_561_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X23 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X24 a_299_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 a_1316_47# a_711_307# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 VPWR a_711_307# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 Q_N a_1316_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dlrtn_1 D GATE_N RESET_B VGND VNB VPB VPWR Q
X0 a_561_413# a_27_47# a_682_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_682_413# a_724_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_561_413# a_193_47# a_659_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X3 VGND a_724_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VPWR a_299_47# a_465_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 a_465_369# a_193_47# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_724_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_659_47# a_724_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_299_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 a_724_21# a_561_413# a_942_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_942_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VGND a_299_47# a_465_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_27_47# GATE_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_27_47# GATE_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X15 VPWR a_561_413# a_724_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 a_465_47# a_27_47# a_561_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X17 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 a_299_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 VPWR a_724_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dlrtn_2 D GATE_N RESET_B VGND VNB VPB VPWR Q
X0 a_560_47# a_27_47# a_645_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_645_413# a_711_307# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 Q a_711_307# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR a_299_47# a_465_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X4 a_465_369# a_193_47# a_560_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 VGND a_711_307# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_299_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 VPWR a_560_47# a_711_307# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_560_47# a_193_47# a_658_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X9 VPWR a_711_307# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_658_47# a_711_307# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_711_307# a_560_47# a_941_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VGND a_299_47# a_465_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_27_47# GATE_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_27_47# GATE_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X16 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X17 a_299_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_465_47# a_27_47# a_560_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X19 Q a_711_307# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 a_941_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 a_711_307# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dlrtn_4 D GATE_N RESET_B VGND VNB VPB VPWR Q
X0 a_562_413# a_27_47# a_683_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_683_413# a_725_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_725_21# a_562_413# a_943_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VGND a_725_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VPWR a_300_47# a_466_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 a_466_369# a_193_47# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_725_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 Q a_725_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_300_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 a_943_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 Q a_725_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 Q a_725_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VGND a_300_47# a_466_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 Q a_725_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_466_47# a_27_47# a_562_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X15 a_300_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_562_413# a_193_47# a_660_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X17 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_27_47# GATE_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 VPWR a_725_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 a_27_47# GATE_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X21 VGND a_725_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X23 VPWR a_562_413# a_725_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X24 a_660_47# a_725_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 VPWR a_725_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dlrtp_1 D GATE RESET_B VGND VNB VPB VPWR Q
X0 VPWR a_560_425# a_711_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_711_21# a_560_425# a_929_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_711_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VPWR a_299_47# a_465_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X4 a_299_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 a_654_47# a_711_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VPWR a_711_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_465_369# a_27_47# a_560_425# VPB sky130_fd_pr__pfet_01v8_hvt w=360000u l=150000u
X8 a_465_47# a_193_47# a_560_425# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_560_425# a_27_47# a_654_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_664_425# a_711_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 VGND a_299_47# a_465_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_27_47# GATE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_27_47# GATE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X15 VGND a_711_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X17 a_560_425# a_193_47# a_664_425# VPB sky130_fd_pr__pfet_01v8_hvt w=360000u l=150000u
X18 a_299_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_929_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dlrtp_2 D GATE RESET_B VGND VNB VPB VPWR Q
X0 a_560_47# a_193_47# a_644_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_644_413# a_711_307# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_711_307# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 Q a_711_307# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_465_369# a_27_47# a_560_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 VPWR a_299_47# a_465_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X6 a_940_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VGND a_711_307# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_299_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 VPWR a_711_307# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_560_47# a_27_47# a_657_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X11 VGND a_299_47# a_465_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VPWR a_560_47# a_711_307# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_27_47# GATE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_27_47# GATE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X16 a_657_47# a_711_307# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 a_299_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_465_47# a_193_47# a_560_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X20 a_711_307# a_560_47# a_940_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 Q a_711_307# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dlrtp_4 D GATE RESET_B VGND VNB VPB VPWR Q
X0 a_562_413# a_193_47# a_683_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_683_413# a_725_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_725_21# a_562_413# a_943_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VGND a_725_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VPWR a_300_47# a_466_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 a_466_369# a_27_47# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_725_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 Q a_725_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_300_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 a_943_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 Q a_725_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 Q a_725_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VGND a_300_47# a_466_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 Q a_725_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_466_47# a_193_47# a_562_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X15 a_300_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_562_413# a_27_47# a_660_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X17 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_27_47# GATE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 VPWR a_725_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 a_27_47# GATE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X21 VGND a_725_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X23 VPWR a_562_413# a_725_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X24 a_660_47# a_725_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 VPWR a_725_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dlxbn_1 D GATE_N VGND VNB VPB VPWR Q Q_N
X0 VGND a_1124_47# Q_N VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_716_21# a_560_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VGND a_716_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_560_47# a_27_47# a_674_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_674_413# a_716_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_470_369# a_193_47# a_560_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_560_47# a_193_47# a_651_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X7 VPWR a_716_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_299_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 a_1124_47# a_716_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X10 VPWR a_299_47# a_470_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X11 VGND a_299_47# a_465_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_27_47# GATE_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 VPWR a_1124_47# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_27_47# GATE_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X16 a_651_47# a_716_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 a_299_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_465_47# a_27_47# a_560_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X20 a_716_21# a_560_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 a_1124_47# a_716_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dlxbn_2 D GATE_N VGND VNB VPB VPWR Q Q_N
X0 VPWR a_728_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_663_47# a_728_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VGND a_1223_47# Q_N VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_728_21# a_565_413# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_565_413# a_27_47# a_686_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_686_413# a_728_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 VPWR a_303_47# a_469_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 a_469_369# a_193_47# a_565_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 Q a_728_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_303_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X10 VGND a_728_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VGND a_303_47# a_469_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_469_47# a_27_47# a_565_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X13 a_565_413# a_193_47# a_663_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X14 Q_N a_1223_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_303_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_27_47# GATE_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_27_47# GATE_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X19 a_1223_47# a_728_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X20 Q a_728_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X22 Q_N a_1223_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 a_1223_47# a_728_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 VPWR a_1223_47# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 a_728_21# a_565_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dlxbp_1 D GATE VGND VNB VPB VPWR Q Q_N
X0 VGND a_1124_47# Q_N VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_716_21# a_560_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_560_47# a_193_47# a_648_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_467_369# a_27_47# a_560_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 VPWR a_299_47# a_467_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 VGND a_716_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_648_413# a_716_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_299_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X8 a_560_47# a_27_47# a_651_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X9 VPWR a_716_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_1124_47# a_716_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X11 VGND a_299_47# a_465_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_27_47# GATE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 VPWR a_1124_47# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_27_47# GATE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X16 a_651_47# a_716_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 a_299_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_465_47# a_193_47# a_560_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X20 a_716_21# a_560_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 a_1124_47# a_716_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dlxtn_1 D GATE_N VGND VNB VPB VPWR Q
X0 a_560_47# a_27_47# a_644_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_715_21# a_560_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_650_47# a_715_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_465_369# a_193_47# a_560_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 VPWR a_715_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VPWR a_299_47# a_465_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X6 a_715_21# a_560_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_299_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X8 a_644_413# a_715_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 VGND a_299_47# a_465_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_560_47# a_193_47# a_650_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X12 a_27_47# GATE_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_27_47# GATE_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X14 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X15 a_299_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_465_47# a_27_47# a_560_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X17 VGND a_715_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dlxtn_2 D GATE_N VGND VNB VPB VPWR Q
X0 VPWR a_728_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_663_47# a_728_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_728_21# a_565_413# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_565_413# a_27_47# a_686_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_686_413# a_728_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 VPWR a_303_47# a_469_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X6 a_469_369# a_193_47# a_565_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 Q a_728_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_303_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 VGND a_728_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VGND a_303_47# a_469_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_469_47# a_27_47# a_565_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X12 a_565_413# a_193_47# a_663_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X13 a_303_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_27_47# GATE_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_27_47# GATE_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X17 Q a_728_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X19 a_728_21# a_565_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dlxtn_4 D GATE_N VGND VNB VPB VPWR Q
X0 a_561_413# a_27_47# a_682_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_682_413# a_724_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 VGND a_724_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_561_413# a_193_47# a_659_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X4 Q a_724_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 Q a_724_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR a_299_47# a_465_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 a_465_369# a_193_47# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_659_47# a_724_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VPWR a_724_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_299_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X11 VPWR a_724_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_724_21# a_561_413# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_724_21# a_561_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 VGND a_724_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 VGND a_299_47# a_465_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_27_47# GATE_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 Q a_724_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_27_47# GATE_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X20 a_465_47# a_27_47# a_561_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X21 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X22 a_299_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 Q a_724_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dlxtp_1 D GATE VGND VNB VPB VPWR Q
X0 a_560_47# a_193_47# a_644_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_713_21# a_560_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_560_47# a_27_47# a_659_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X3 a_465_369# a_27_47# a_560_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 VPWR a_299_47# a_465_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 a_644_413# a_713_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_713_21# a_560_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_299_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X8 VGND a_713_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VGND a_299_47# a_465_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_659_47# a_713_21# VGND VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X11 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_27_47# GATE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_27_47# GATE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X14 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X15 a_299_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_465_47# a_193_47# a_560_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X17 VPWR a_713_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
X0 VPWR a_299_93# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_299_93# a_193_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_299_93# a_193_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 VGND a_299_93# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dlygate4sd2_1 A VGND VNB VPB VPWR X
X0 a_327_47# a_221_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=180000u
X1 a_327_47# a_221_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X2 VGND a_327_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR a_49_47# a_221_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X4 a_49_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VGND a_49_47# a_221_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=180000u
X6 a_49_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VPWR a_327_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
X0 a_391_47# a_285_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=500000u
X1 VPWR a_49_47# a_285_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=500000u
X2 a_49_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VPWR a_391_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VGND a_391_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VGND a_49_47# a_285_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=500000u
X6 a_391_47# a_285_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=500000u
X7 a_49_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
X0 a_381_47# X VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_381_47# X VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_664_47# a_558_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_62_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VPWR a_664_47# a_841_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND a_381_47# a_558_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VGND a_62_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VPWR a_62_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_664_47# a_558_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_62_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 VPWR a_381_47# a_558_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 VGND a_664_47# a_841_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dlymetal6s4s_1 A VGND VNB VPB VPWR X
X0 a_664_47# X VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_345_47# a_239_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_62_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VGND a_345_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VPWR a_664_47# a_841_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_345_47# a_239_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 VGND a_62_47# a_239_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VPWR a_62_47# a_239_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_664_47# X VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VPWR a_345_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_62_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 VGND a_664_47# a_841_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dlymetal6s6s_1 A VGND VNB VPB VPWR X
X0 a_346_47# a_240_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_63_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VPWR a_63_47# a_240_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VPWR a_629_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VGND a_346_47# a_523_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VGND a_63_47# a_240_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_629_47# a_523_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_629_47# a_523_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VGND a_629_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_346_47# a_240_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 VPWR a_346_47# a_523_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_63_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
X0 VGND TE_B a_193_369# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VGND a_193_369# a_531_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_531_47# a_27_47# Z VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR TE_B a_383_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_383_297# a_27_47# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X6 VPWR TE_B a_193_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__ebufn_2 A TE_B VGND VNB VPB VPWR Z
X0 VGND TE_B a_214_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_392_47# a_27_47# Z VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VPWR TE_B a_214_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X3 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X4 Z a_27_47# a_320_309# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND a_214_47# a_392_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR TE_B a_320_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X7 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_320_309# a_27_47# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_392_47# a_214_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_320_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X11 Z a_27_47# a_392_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__ebufn_4 A TE_B VGND VNB VPB VPWR Z
X0 a_393_47# a_214_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VGND TE_B a_214_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 Z a_27_47# a_320_309# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 Z a_27_47# a_393_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 Z a_27_47# a_320_309# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND a_214_47# a_393_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 Z a_27_47# a_393_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VGND a_214_47# a_393_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VPWR TE_B a_214_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_320_309# a_27_47# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_393_47# a_214_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VPWR TE_B a_320_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X12 VPWR TE_B a_320_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X13 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_320_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X16 a_320_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X17 a_393_47# a_27_47# Z VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 a_320_309# a_27_47# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_393_47# a_27_47# Z VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
X0 a_407_309# a_116_47# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VPWR TE_B a_407_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X2 a_455_47# a_116_47# Z VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_455_47# a_116_47# Z VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VPWR TE_B a_407_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X5 VPWR TE_B a_407_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X6 Z a_116_47# a_407_309# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 Z a_116_47# a_407_309# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND a_301_47# a_455_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 Z a_116_47# a_455_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VGND a_301_47# a_455_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_455_47# a_301_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VPWR TE_B a_407_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X13 a_455_47# a_301_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_116_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_407_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X16 VGND a_301_47# a_455_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 VPWR A a_116_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 a_407_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X19 VGND A a_116_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_116_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 a_455_47# a_116_47# Z VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 Z a_116_47# a_407_309# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 VGND a_301_47# a_455_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 Z a_116_47# a_455_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 a_407_309# a_116_47# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 Z a_116_47# a_455_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 VPWR TE_B a_301_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X28 VGND TE_B a_301_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 a_455_47# a_301_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 a_455_47# a_116_47# Z VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 a_407_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X32 Z a_116_47# a_407_309# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X33 a_455_47# a_301_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X34 a_407_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X35 a_407_309# a_116_47# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X36 Z a_116_47# a_455_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X37 a_407_309# a_116_47# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__edfxbp_1 CLK D DE VGND VNB VPB VPWR Q Q_N
X0 a_986_413# a_27_47# a_1077_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 VGND a_1591_413# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_729_47# a_791_264# a_299_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VGND a_986_413# a_1150_159# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X4 a_299_47# D a_381_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 a_381_369# a_423_343# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X6 a_791_264# a_1591_413# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_1591_413# a_193_47# a_1675_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 VGND a_1150_159# a_1514_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VPWR DE a_729_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X10 VPWR a_986_413# a_1150_159# VPB sky130_fd_pr__pfet_01v8_hvt w=750000u l=150000u
X11 a_381_47# DE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_1500_413# a_27_47# a_1591_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X13 a_1675_413# a_791_264# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X14 a_729_369# a_791_264# a_299_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X15 a_423_343# DE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 VPWR a_1591_413# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 a_1101_47# a_1150_159# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_791_264# a_1591_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X19 a_1077_413# a_1150_159# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X20 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 a_299_47# a_27_47# a_986_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X22 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 VGND a_423_343# a_729_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 a_986_413# a_193_47# a_1101_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X25 VGND a_791_264# Q_N VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X27 VPWR a_791_264# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X28 a_1591_413# a_27_47# a_1717_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X29 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X30 a_299_47# a_193_47# a_986_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X31 a_299_47# D a_381_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X32 a_423_343# DE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X33 a_1514_47# a_193_47# a_1591_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X34 VPWR a_1150_159# a_1500_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X35 a_1717_47# a_791_264# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__edfxtp_1 CLK D DE VGND VNB VPB VPWR Q
X0 a_986_413# a_27_47# a_1077_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_791_264# a_1591_413# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_729_47# a_791_264# a_299_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_791_264# a_1591_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X4 VGND a_986_413# a_1150_159# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X5 a_299_47# D a_381_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X6 a_381_369# a_423_343# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 a_1591_413# a_193_47# a_1675_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 VGND a_1150_159# a_1514_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VGND a_1591_413# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VPWR DE a_729_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X11 VPWR a_986_413# a_1150_159# VPB sky130_fd_pr__pfet_01v8_hvt w=750000u l=150000u
X12 a_381_47# DE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_1500_413# a_27_47# a_1591_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X14 a_1675_413# a_791_264# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 a_729_369# a_791_264# a_299_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X16 a_423_343# DE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_1101_47# a_1150_159# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_1077_413# a_1150_159# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X19 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_299_47# a_27_47# a_986_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X21 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 VGND a_423_343# a_729_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_986_413# a_193_47# a_1101_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X24 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X25 a_1591_413# a_27_47# a_1717_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X26 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X27 a_299_47# a_193_47# a_986_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X28 a_299_47# D a_381_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 a_423_343# DE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X30 a_1514_47# a_193_47# a_1591_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X31 VPWR a_1591_413# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X32 VPWR a_1150_159# a_1500_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X33 a_1717_47# a_791_264# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__einvn_0 A TE_B VGND VNB VPB VPWR Z
X0 a_30_47# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 VPWR TE_B a_215_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 a_215_369# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X3 a_215_47# A Z VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_30_47# TE_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VGND a_30_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__einvn_1 A TE_B VGND VNB VPB VPWR Z
X0 a_204_297# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_27_47# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 VGND a_27_47# a_286_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR TE_B a_204_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_27_47# TE_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_286_47# A Z VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__einvn_2 A TE_B VGND VNB VPB VPWR Z
X0 VGND a_27_47# a_214_120# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 Z A a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_204_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X3 a_214_120# A Z VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VPWR TE_B a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X5 a_204_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_214_120# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_27_47# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X8 a_27_47# TE_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 Z A a_214_120# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__einvn_4 A TE_B VGND VNB VPB VPWR Z
X0 Z A a_215_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_215_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_204_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_204_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X4 a_204_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X5 VPWR TE_B a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X6 VPWR TE_B a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X7 Z A a_215_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 Z A a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VGND a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 Z A a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_215_47# A Z VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_215_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_215_47# A Z VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_204_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_27_47# TE_B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_27_47# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 VGND a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__einvn_8 A TE_B VGND VNB VPB VPWR Z
X0 VGND a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 Z A a_215_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 Z A a_215_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_215_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_215_47# A Z VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_215_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_215_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_204_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_204_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X9 Z A a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_204_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X11 Z A a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_215_47# A Z VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VPWR TE_B a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X14 a_215_47# A Z VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 VGND a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VPWR TE_B a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X17 VPWR TE_B a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X18 VGND a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 Z A a_215_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 Z A a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 a_215_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 a_27_47# TE_B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 a_204_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X24 a_204_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 Z A a_215_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 VPWR TE_B a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X27 a_204_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X28 a_27_47# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X29 VGND a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 a_204_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X31 Z A a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X32 a_215_47# A Z VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X33 a_204_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__einvp_1 A TE VGND VNB VPB VPWR Z
X0 a_276_297# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VGND TE a_204_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_27_47# TE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_204_47# A Z VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VPWR a_27_47# a_276_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_27_47# TE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__einvp_2 A TE VGND VNB VPB VPWR Z
X0 a_215_309# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X1 a_204_47# TE VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_215_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VGND TE a_204_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_204_47# A Z VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VPWR a_27_47# a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X6 Z A a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_27_47# TE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X8 a_27_47# TE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 Z A a_204_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__einvp_4 A TE VGND VNB VPB VPWR Z
X0 VPWR a_27_47# a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X1 VGND TE a_193_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 Z A a_193_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_215_309# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X4 a_215_309# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X5 a_193_47# TE VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_215_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VPWR a_27_47# a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X8 Z A a_193_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 Z A a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 Z A a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_193_47# A Z VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VGND TE a_193_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_193_47# A Z VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_215_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_27_47# TE VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_27_47# TE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 a_193_47# TE VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__einvp_8 A TE VGND VNB VPB VPWR Z
X0 VPWR a_27_47# a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X1 VGND TE a_193_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 Z A a_193_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_215_309# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X4 Z A a_193_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_215_309# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X6 a_215_309# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X7 a_193_47# TE VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_193_47# A Z VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VPWR a_27_47# a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X10 a_215_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_193_47# TE VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 Z A a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 Z A a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_193_47# A Z VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 VGND TE a_193_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_193_47# A Z VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 VPWR a_27_47# a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X18 VGND TE a_193_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 VPWR a_27_47# a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X20 Z A a_193_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 a_215_309# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=150000u
X22 Z A a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 VGND TE a_193_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 a_27_47# TE VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 a_215_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 a_215_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 Z A a_193_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 a_215_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X29 a_27_47# TE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X30 a_193_47# TE VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 a_193_47# TE VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X32 Z A a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X33 a_193_47# A Z VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__fa_1 A B CIN VGND VNB VPB VPWR COUT SUM
X0 VGND A a_208_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VGND B a_382_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_1163_413# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_208_413# B a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_382_413# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 VPWR A a_738_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_76_199# CIN a_382_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_738_413# CIN VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_995_47# CIN a_1091_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 VPWR B a_382_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_1091_413# B a_1163_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 VGND A a_738_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_382_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 VGND B a_738_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 VPWR a_995_47# SUM VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_738_47# CIN VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_738_47# a_76_199# a_995_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_76_199# CIN a_382_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_1091_47# B a_1163_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_738_413# a_76_199# a_995_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X20 VGND a_995_47# SUM VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 VPWR B a_738_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X22 a_1163_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 VPWR A a_208_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X24 COUT a_76_199# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 COUT a_76_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 a_208_47# B a_76_199# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 a_995_47# CIN a_1091_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__fa_2 A B CIN VGND VNB VPB VPWR COUT SUM
X0 a_80_21# CIN a_473_371# VPB sky130_fd_pr__pfet_01v8_hvt w=630000u l=150000u
X1 a_289_371# B a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt w=630000u l=150000u
X2 a_1086_47# CIN a_1171_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X3 a_829_47# CIN VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VPWR B a_473_371# VPB sky130_fd_pr__pfet_01v8_hvt w=630000u l=150000u
X5 VGND A a_294_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_80_21# CIN a_473_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VPWR a_80_21# COUT VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND a_1086_47# SUM VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VGND a_80_21# COUT VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_1266_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_1194_47# B a_1266_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 COUT a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VGND B a_829_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_294_47# B a_80_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 VPWR a_1086_47# SUM VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 SUM a_1086_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 VGND B a_473_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 VPWR A a_289_371# VPB sky130_fd_pr__pfet_01v8_hvt w=630000u l=150000u
X19 a_829_47# a_80_21# a_1086_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 VPWR B a_829_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X21 SUM a_1086_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 VPWR A a_829_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X23 a_1086_47# CIN a_1194_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 a_829_369# a_80_21# a_1086_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X25 a_1266_371# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=630000u l=150000u
X26 a_829_369# CIN VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X27 a_473_371# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=630000u l=150000u
X28 a_1171_369# B a_1266_371# VPB sky130_fd_pr__pfet_01v8_hvt w=630000u l=150000u
X29 VGND A a_829_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X30 COUT a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X31 a_473_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__fa_4 A B CIN VGND VNB VPB VPWR COUT SUM
X0 a_79_21# CIN a_658_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X1 a_456_371# B a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=630000u l=150000u
X2 VPWR a_1271_47# SUM VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VPWR B a_1014_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X4 a_658_369# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 a_1271_47# CIN a_1356_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X6 COUT a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_1014_369# a_79_21# a_1271_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X8 a_461_47# B a_79_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VGND B a_658_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_1356_369# B a_1451_371# VPB sky130_fd_pr__pfet_01v8_hvt w=630000u l=150000u
X11 a_79_21# CIN a_658_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_1379_47# B a_1451_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 VGND a_1271_47# SUM VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VGND B a_1014_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 SUM a_1271_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_1451_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 VGND A a_1014_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 SUM a_1271_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 VPWR B a_658_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X20 VGND a_79_21# COUT VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 VPWR A a_456_371# VPB sky130_fd_pr__pfet_01v8_hvt w=630000u l=150000u
X22 a_1014_47# a_79_21# a_1271_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_1014_369# CIN VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X24 COUT a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 SUM a_1271_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 VPWR a_79_21# COUT VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 VGND a_79_21# COUT VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 VPWR a_79_21# COUT VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X29 VPWR A a_1014_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X30 SUM a_1271_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X31 VGND a_1271_47# SUM VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X32 COUT a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X33 VGND A a_461_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 a_1014_47# CIN VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 COUT a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X36 a_1451_371# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=630000u l=150000u
X37 VPWR a_1271_47# SUM VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X38 a_658_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X39 a_1271_47# CIN a_1379_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__fah_1 A B CI VGND VNB VPB VPWR COUT SUM
X0 a_1332_297# a_1008_47# a_1262_49# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X1 a_1332_297# a_1008_47# a_508_297# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X2 COUT a_1332_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_719_47# a_508_297# a_310_49# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X4 a_1262_49# a_1008_47# a_1617_49# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X5 a_1262_49# CI VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VGND A a_67_199# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X7 a_719_47# a_508_297# a_27_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X8 a_27_47# a_67_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_310_49# A VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X10 a_1262_49# CI VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X11 a_27_47# a_508_297# a_1008_47# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X12 a_1617_49# a_719_47# a_1262_49# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X13 a_310_49# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_310_49# a_508_297# a_1008_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X15 a_1640_380# a_1008_47# a_1617_49# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X16 a_1008_47# B a_310_49# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X17 a_1617_49# a_719_47# a_1640_380# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X18 VPWR B a_508_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_508_297# a_719_47# a_1332_297# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X20 VPWR A a_67_199# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 VGND B a_508_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 VGND a_1262_49# a_1640_380# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X23 a_27_47# a_67_199# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 VPWR a_1617_49# SUM VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 a_27_47# B a_719_47# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X26 a_1008_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X27 VPWR a_1262_49# a_1640_380# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X28 VGND a_1617_49# SUM VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 COUT a_1332_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X30 a_310_49# B a_719_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X31 a_1262_49# a_719_47# a_1332_297# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__fahcin_1 A B CIN VGND VNB VPB VPWR COUT SUM
X0 VGND CIN a_1636_315# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_1251_49# CIN VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_67_199# a_489_21# a_721_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X3 a_1565_49# a_721_47# a_1647_49# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X4 a_1565_49# a_1636_315# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X5 a_1251_49# CIN VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X6 a_1647_49# a_434_49# a_1565_49# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X7 a_489_21# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_27_47# a_67_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_1565_49# a_1636_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VPWR CIN a_1636_315# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_27_47# a_67_199# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X12 VGND a_489_21# a_1142_49# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X13 VGND a_1647_49# SUM VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VPWR A a_67_199# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_721_47# B a_67_199# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X16 a_434_49# a_489_21# a_67_199# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X17 a_1142_49# a_434_49# COUT VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X18 a_67_199# B a_434_49# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X19 a_434_49# a_489_21# a_27_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X20 a_27_47# a_489_21# a_721_47# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X21 a_1647_49# a_434_49# a_1636_315# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X22 a_489_21# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 a_721_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X24 a_1251_49# a_434_49# COUT VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X25 COUT a_721_47# a_1142_49# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X26 COUT a_721_47# a_1251_49# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X27 VPWR a_489_21# a_1142_49# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X28 VPWR a_1647_49# SUM VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X29 VGND A a_67_199# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 a_27_47# B a_434_49# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X31 a_1636_315# a_721_47# a_1647_49# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__fahcon_1 A B CI VGND VNB VPB VPWR COUT_N SUM
X0 COUT_N a_726_47# a_1261_49# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X1 VPWR B a_1144_49# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_1261_49# CI VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_28_47# a_67_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_726_47# B a_67_199# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X5 a_28_47# a_67_199# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X6 a_1710_49# a_434_49# a_1589_49# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X7 a_1261_49# a_434_49# COUT_N VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X8 VPWR A a_67_199# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 COUT_N a_726_47# a_1144_49# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X10 VPWR CI a_1589_49# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 VPWR a_1710_49# SUM VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_434_49# a_488_21# a_67_199# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X13 a_1634_315# a_726_47# a_1710_49# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X14 a_726_47# B a_28_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X15 a_488_21# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VGND CI a_1589_49# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 a_1634_315# a_1589_49# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X18 a_1261_49# CI VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X19 a_67_199# B a_434_49# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X20 a_1710_49# a_434_49# a_1634_315# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X21 a_1144_49# a_434_49# COUT_N VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X22 a_67_199# a_488_21# a_726_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X23 VGND B a_1144_49# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X24 VGND a_1710_49# SUM VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 a_28_47# a_488_21# a_726_47# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X26 a_488_21# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 a_434_49# a_488_21# a_28_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X28 a_1589_49# a_726_47# a_1710_49# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X29 VGND A a_67_199# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 a_28_47# B a_434_49# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X31 a_1634_315# a_1589_49# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__fill_4 VGND VNB VPB VPWR
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__fill_8 VGND VNB VPB VPWR
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__ha_1 A B VGND VNB VPB VPWR COUT SUM
X0 a_250_199# B a_674_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_79_21# a_250_199# a_297_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_250_199# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 VPWR a_250_199# COUT VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VGND A a_297_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_79_21# B a_376_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_376_413# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 SUM a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_674_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 SUM a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VPWR a_250_199# a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 a_297_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VGND a_250_199# COUT VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VPWR B a_250_199# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__ha_2 A B VGND VNB VPB VPWR COUT SUM
X0 VPWR a_342_199# COUT VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_766_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 SUM a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_389_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 COUT a_342_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND a_342_199# COUT VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_79_21# B a_468_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 a_468_369# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X8 VPWR a_342_199# a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 a_342_199# B a_766_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_79_21# a_342_199# a_389_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 SUM a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VGND a_79_21# SUM VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VPWR B a_342_199# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X14 VPWR a_79_21# SUM VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_342_199# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X16 COUT a_342_199# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 VGND A a_389_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__ha_4 A B VGND VNB VPB VPWR COUT SUM
X0 VGND a_514_199# COUT VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_890_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_514_199# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_717_297# B a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_79_21# a_514_199# a_467_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 SUM a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_1167_47# B a_514_199# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 COUT a_514_199# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_79_21# B a_890_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_467_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_79_21# a_514_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_514_199# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VGND A a_1167_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_1325_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VPWR B a_514_199# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_467_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_467_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 a_514_199# B a_1325_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 VGND a_79_21# SUM VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 a_467_47# a_514_199# a_79_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 VGND a_514_199# COUT VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 VPWR a_514_199# COUT VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 VPWR a_514_199# COUT VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 VGND B a_467_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 COUT a_514_199# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 SUM a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 VPWR a_79_21# SUM VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 VPWR A a_717_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X28 VGND a_79_21# SUM VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 COUT a_514_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X30 COUT a_514_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X31 VPWR a_79_21# SUM VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X32 SUM a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X33 SUM a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X34 VPWR a_514_199# a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X35 VPWR A a_514_199# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
X0 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
X0 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
X0 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X24 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X28 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X29 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_bleeder_1 SHORT VGND VNB VPB VPWR
X0 a_291_105# SHORT a_363_105# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X1 a_219_105# SHORT a_291_105# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X2 VGND SHORT a_147_105# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X3 a_363_105# SHORT VPWR VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X4 a_147_105# SHORT a_219_105# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_clkbufkapwr_1 A KAPWR VGND VNB VPB VPWR X
X0 VGND A a_75_212# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X1 X a_75_212# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
X2 X a_75_212# VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X3 KAPWR A a_75_212# VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_clkbufkapwr_2 A KAPWR VGND VNB VPB VPWR X
X0 a_27_47# A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 X a_27_47# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 KAPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_clkbufkapwr_4 A KAPWR VGND VNB VPB VPWR X
X0 KAPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 X a_27_47# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_27_47# A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 X a_27_47# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 KAPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_clkbufkapwr_8 A KAPWR VGND VNB VPB VPWR X
X0 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_110_47# A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 KAPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 X a_110_47# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 KAPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 KAPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 X a_110_47# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 KAPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 KAPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 X a_110_47# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 X a_110_47# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_clkbufkapwr_16 A KAPWR VGND VNB VPB VPWR X
X0 KAPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_110_47# A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 KAPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 X a_110_47# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 KAPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_110_47# A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 KAPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 KAPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 X a_110_47# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 X a_110_47# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 X a_110_47# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 KAPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X24 KAPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 X a_110_47# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 KAPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X29 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X30 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 X a_110_47# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X32 X a_110_47# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X33 X a_110_47# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X34 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 KAPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X36 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X37 KAPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X38 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X39 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_clkinvkapwr_1 A KAPWR VGND VNB VPB VPWR Y
X0 Y A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 KAPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_clkinvkapwr_2 A KAPWR VGND VNB VPB VPWR Y
X0 Y A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 KAPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 Y A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_clkinvkapwr_4 A KAPWR VGND VNB VPB VPWR Y
X0 KAPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 Y A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 KAPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 Y A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 Y A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 KAPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_clkinvkapwr_8 A KAPWR VGND VNB VPB VPWR Y
X0 Y A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 Y A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 Y A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 Y A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 KAPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 KAPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 KAPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 KAPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 KAPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 KAPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 Y A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 Y A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_clkinvkapwr_16 A KAPWR VGND VNB VPB VPWR Y
X0 Y A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 KAPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 KAPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 Y A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 Y A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 KAPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 KAPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 KAPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 Y A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 KAPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 KAPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 KAPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 Y A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 Y A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 KAPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 Y A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 Y A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 Y A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X28 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 KAPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X30 Y A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X31 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X32 KAPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X33 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 Y A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X35 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X36 Y A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X37 KAPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X38 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X39 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_decapkapwr_3 KAPWR VGND VNB VPB VPWR
X0 KAPWR VGND KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=870000u l=590000u
X1 VGND KAPWR VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=590000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_decapkapwr_4 KAPWR VGND VNB VPB VPWR
X0 KAPWR VGND KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=870000u l=1.05e+06u
X1 VGND KAPWR VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=1.05e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_decapkapwr_6 KAPWR VGND VNB VPB VPWR
X0 KAPWR VGND KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=870000u l=1.97e+06u
X1 VGND KAPWR VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=1.97e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_decapkapwr_8 KAPWR VGND VNB VPB VPWR
X0 KAPWR VGND KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=870000u l=2.89e+06u
X1 VGND KAPWR VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=2.89e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_decapkapwr_12 KAPWR VGND VNB VPB VPWR
X0 KAPWR VGND KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=870000u l=4.73e+06u
X1 VGND KAPWR VGND VNB sky130_fd_pr__nfet_01v8 w=550000u l=4.73e+06u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_inputiso0n_1 A SLEEP_B VGND VNB VPB VPWR X
X0 VGND a_59_75# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VPWR A a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_59_75# A a_145_75# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_59_75# SLEEP_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_145_75# SLEEP_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VPWR a_59_75# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_inputiso0p_1 A SLEEP VGND VNB VPB VPWR X
X0 a_207_413# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 VPWR a_207_413# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VGND a_207_413# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_207_413# a_27_413# a_297_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_27_413# SLEEP VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 VPWR a_27_413# a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 VGND SLEEP a_27_413# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_297_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_inputiso1n_1 A SLEEP_B VGND VNB VPB VPWR X
X0 a_219_297# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_27_53# SLEEP_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VGND a_27_53# a_219_297# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VGND a_219_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_219_297# a_27_53# a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_301_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 VPWR SLEEP_B a_27_53# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VPWR a_219_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_inputiso1p_1 A SLEEP VGND VNB VPB VPWR X
X0 a_150_297# SLEEP VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 VGND a_68_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_68_297# SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_68_297# A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 VPWR a_68_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_inputisolatch_1 D SLEEP_B VGND VNB VPB VPWR Q
X0 a_560_413# a_629_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 VPWR a_476_47# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_575_47# a_629_21# VGND VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X3 a_476_47# a_193_47# a_560_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_476_47# a_27_47# a_575_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X5 a_381_47# a_193_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X6 VGND a_476_47# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VPWR D a_381_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X8 a_27_47# SLEEP_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=550000u l=150000u
X9 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=550000u l=150000u
X10 a_629_21# a_476_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_27_47# SLEEP_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 VGND D a_381_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_629_21# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_381_369# a_27_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_isobufsrc_1 A SLEEP VGND VNB VPB VPWR X
X0 a_74_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 X a_74_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_74_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VPWR SLEEP a_265_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_265_297# a_74_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_isobufsrc_2 A SLEEP VGND VNB VPB VPWR X
X0 X a_251_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VPWR SLEEP a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 X a_251_21# a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VGND a_251_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_27_297# a_251_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_27_297# SLEEP VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_251_21# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_251_21# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_isobufsrc_4 A SLEEP VGND VNB VPB VPWR X
X0 a_27_297# a_419_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VPWR SLEEP a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VPWR SLEEP a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 X a_419_21# a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_27_297# SLEEP VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_27_297# SLEEP VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 X a_419_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_27_297# a_419_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 X a_419_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_419_21# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 X a_419_21# a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_419_21# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VGND a_419_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 VGND a_419_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_isobufsrc_8 A SLEEP VGND VNB VPB VPWR X
X0 a_321_297# SLEEP X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 X a_123_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 X a_123_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VPWR A a_123_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND a_123_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR a_123_297# a_321_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_321_297# a_123_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 X a_123_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_321_297# a_123_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_321_297# a_123_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_321_297# SLEEP X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_321_297# SLEEP X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VPWR a_123_297# a_321_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 X a_123_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 X SLEEP a_321_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_123_297# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 X SLEEP a_321_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 VGND a_123_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 VGND A a_123_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 VGND a_123_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 VGND a_123_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 VPWR a_123_297# a_321_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 VPWR a_123_297# a_321_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X29 a_123_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X30 X SLEEP a_321_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X31 X SLEEP a_321_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X32 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X33 a_321_297# a_123_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X34 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X35 a_321_297# SLEEP X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_isobufsrc_16 A SLEEP VGND VNB VPB VPWR X
X0 X SLEEP a_505_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VGND a_143_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VPWR A a_143_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_505_297# a_143_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 X a_143_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 X a_143_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_505_297# a_143_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_143_297# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_505_297# SLEEP X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 X a_143_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VPWR a_143_297# a_505_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 X SLEEP a_505_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VPWR a_143_297# a_505_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 VPWR a_143_297# a_505_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 VGND A a_143_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 VPWR a_143_297# a_505_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 VGND a_143_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 X SLEEP a_505_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 a_505_297# SLEEP X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 a_505_297# SLEEP X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X24 X a_143_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 a_143_297# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 X a_143_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 X SLEEP a_505_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X29 a_143_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X30 a_143_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X31 a_505_297# a_143_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X32 X SLEEP a_505_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X33 VGND a_143_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X34 X SLEEP a_505_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X35 a_505_297# SLEEP X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X36 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X37 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X38 VPWR A a_143_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X39 VPWR a_143_297# a_505_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X40 a_505_297# SLEEP X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X41 X a_143_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X42 VPWR a_143_297# a_505_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X43 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X44 VPWR a_143_297# a_505_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X45 X a_143_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X46 VPWR a_143_297# a_505_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X47 a_505_297# a_143_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X48 VGND a_143_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X49 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X50 a_505_297# a_143_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X51 VGND A a_143_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X52 VGND a_143_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X53 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X54 X SLEEP a_505_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X55 VGND a_143_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X56 VGND a_143_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X57 a_505_297# a_143_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X58 a_505_297# a_143_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X59 a_505_297# SLEEP X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X60 X a_143_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X61 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X62 a_505_297# SLEEP X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X63 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X64 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X65 a_505_297# SLEEP X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X66 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X67 VGND a_143_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X68 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X69 a_505_297# a_143_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X70 X SLEEP a_505_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X71 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_isobufsrckapwr_16 A SLEEP KAPWR VGND VNB VPB VPWR X
X0 VGND a_1122_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VPWR SLEEP a_255_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 KAPWR a_1122_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VGND a_341_47# a_1122_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VGND a_1122_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 X a_1122_47# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_341_47# SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 X a_1122_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 KAPWR a_341_47# a_1122_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VPWR A a_147_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 X a_1122_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VGND SLEEP a_341_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 X a_1122_47# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 X a_1122_47# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_1122_47# a_341_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_255_297# a_147_47# a_341_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 KAPWR a_1122_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 VGND a_341_47# a_1122_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 VGND a_1122_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_1122_47# a_341_47# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 a_341_47# a_147_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 X a_1122_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_1122_47# a_341_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 VGND A a_147_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 X a_1122_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 VGND a_1122_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 KAPWR a_1122_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 X a_1122_47# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X28 KAPWR a_1122_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X29 VGND a_147_47# a_341_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 a_255_297# a_147_47# a_341_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X31 X a_1122_47# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X32 KAPWR a_1122_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X33 X a_1122_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 a_255_297# SLEEP VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X35 X a_1122_47# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X36 a_255_297# SLEEP VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X37 VGND a_1122_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X38 a_341_47# a_147_47# a_255_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X39 X a_1122_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X40 VGND a_1122_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X41 a_341_47# a_147_47# a_255_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X42 VGND a_147_47# a_341_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X43 VGND SLEEP a_341_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X44 X a_1122_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X45 VPWR SLEEP a_255_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X46 KAPWR a_1122_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X47 X a_1122_47# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X48 KAPWR a_1122_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X49 X a_1122_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X50 a_1122_47# a_341_47# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X51 KAPWR a_1122_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X52 X a_1122_47# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X53 VGND a_1122_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X54 KAPWR a_341_47# a_1122_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X55 a_341_47# a_147_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X56 a_341_47# SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X57 VGND a_1122_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_1 A VGND VPB VPWRIN VPWR X
X0 VPWR a_1028_32# X VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
X1 a_714_58# A VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_714_58# a_620_911# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
X3 a_620_911# a_505_297# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_620_911# a_505_297# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VPWRIN A a_505_297# VPWRIN sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VPWR a_620_911# a_1028_32# VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
X7 VGND a_505_297# a_620_911# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VGND a_505_297# a_620_911# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VGND A a_714_58# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_714_58# A VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VGND a_620_911# a_1028_32# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_620_911# a_714_58# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
X13 VGND a_1028_32# X VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VGND A a_505_297# VGND sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 VGND A a_714_58# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_2 A VGND VPB VPWRIN VPWR X
X0 VGND a_1032_911# X VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 X a_1032_911# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 X a_1032_911# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_714_47# a_620_911# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
X4 a_620_911# a_505_297# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_620_911# a_505_297# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VGND A a_714_47# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VPWRIN A a_505_297# VPWRIN sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_714_47# A VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VPWR a_1032_911# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VPWR a_620_911# a_1032_911# VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
X11 VGND a_505_297# a_620_911# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VGND a_505_297# a_620_911# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VGND A a_714_47# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_714_47# A VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 VGND a_620_911# a_1032_911# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_620_911# a_714_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
X17 VGND A a_505_297# VGND sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_4 A VGND VPB VPWRIN VPWR X
X0 VGND a_1032_911# X VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 X a_1032_911# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VPWR a_1032_911# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 X a_1032_911# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_714_47# a_620_911# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
X5 a_620_911# a_505_297# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_620_911# a_505_297# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 X a_1032_911# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND A a_714_47# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VPWRIN A a_505_297# VPWRIN sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_714_47# A VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VPWR a_1032_911# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VPWR a_620_911# a_1032_911# VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
X13 VGND a_1032_911# X VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VGND a_505_297# a_620_911# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 X a_1032_911# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VGND a_505_297# a_620_911# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 VGND A a_714_47# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 a_714_47# A VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 VGND a_620_911# a_1032_911# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_620_911# a_714_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
X21 VGND A a_505_297# VGND sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_4 A LOWLVPWR VGND VNB VPB VPWR X
X0 a_424_82# a_1032_911# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 X a_1032_911# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VPWR a_1032_911# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 X a_1032_911# a_424_82# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_714_47# a_620_911# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
X5 a_620_911# a_505_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_620_911# a_505_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 X a_1032_911# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_424_82# A a_714_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 LOWLVPWR A a_505_297# LOWLVPWR sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_714_47# A a_424_82# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VPWR a_1032_911# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VPWR a_620_911# a_1032_911# VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
X13 a_424_82# a_1032_911# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VGND a_505_297# a_620_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 X a_1032_911# a_424_82# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VGND a_505_297# a_620_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 a_424_82# A a_714_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 a_714_47# A a_424_82# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 VGND a_620_911# a_1032_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_620_911# a_714_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
X21 a_424_82# A a_505_297# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_1 A LOWLVPWR VGND VPB VPWR X
X0 VPWR a_1028_32# X VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
X1 a_714_58# A VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_714_58# a_620_911# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
X3 a_620_911# a_505_297# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_620_911# a_505_297# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 LOWLVPWR A a_505_297# LOWLVPWR sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VPWR a_620_911# a_1028_32# VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
X7 VGND a_505_297# a_620_911# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VGND a_505_297# a_620_911# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VGND A a_714_58# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_714_58# A VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VGND a_620_911# a_1028_32# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_620_911# a_714_58# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
X13 VGND a_1028_32# X VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VGND A a_505_297# VGND sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 VGND A a_714_58# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_2 A LOWLVPWR VGND VPB VPWR X
X0 VGND a_1032_911# X VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 X a_1032_911# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 X a_1032_911# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_714_47# a_620_911# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
X4 a_620_911# a_505_297# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_620_911# a_505_297# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VGND A a_714_47# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 LOWLVPWR A a_505_297# LOWLVPWR sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_714_47# A VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VPWR a_1032_911# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VPWR a_620_911# a_1032_911# VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
X11 VGND a_505_297# a_620_911# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VGND a_505_297# a_620_911# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VGND A a_714_47# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_714_47# A VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 VGND a_620_911# a_1032_911# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_620_911# a_714_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
X17 VGND A a_505_297# VGND sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_4 A LOWLVPWR VGND VPB VPWR X
X0 VGND a_1032_911# X VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 X a_1032_911# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VPWR a_1032_911# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 X a_1032_911# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_714_47# a_620_911# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
X5 a_620_911# a_505_297# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_620_911# a_505_297# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 X a_1032_911# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND A a_714_47# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 LOWLVPWR A a_505_297# LOWLVPWR sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_714_47# A VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VPWR a_1032_911# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VPWR a_620_911# a_1032_911# VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
X13 VGND a_1032_911# X VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VGND a_505_297# a_620_911# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 X a_1032_911# VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VGND a_505_297# a_620_911# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 VGND A a_714_47# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 a_714_47# A VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 VGND a_620_911# a_1032_911# VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_620_911# a_714_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
X21 VGND A a_505_297# VGND sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0






.subckt sky130_fd_sc_hd__macro_sparecell VGND VNB VPB VPWR LO
Xsky130_fd_sc_hd__nand2_2_1 sky130_fd_sc_hd__nor2_2_1/B LO LO VPB VNB VGND VPWR sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__nand2_2_0 sky130_fd_sc_hd__nor2_2_0/A LO LO VPB VNB VGND VPWR sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__inv_2_0 sky130_fd_sc_hd__inv_2_0/A sky130_fd_sc_hd__inv_2_0/Y VPB VNB VPWR VGND sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_1 sky130_fd_sc_hd__inv_2_1/A sky130_fd_sc_hd__inv_2_1/Y VPB VNB VPWR VGND sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__nor2_2_0 sky130_fd_sc_hd__nor2_2_0/A sky130_fd_sc_hd__inv_2_0/A sky130_fd_sc_hd__nor2_2_0/A VPB VNB VGND VPWR sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__nor2_2_1 sky130_fd_sc_hd__nor2_2_1/B sky130_fd_sc_hd__inv_2_1/A sky130_fd_sc_hd__nor2_2_1/B VPB VNB VGND VPWR sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__conb_1_0 VPB VNB VGND VPWR sky130_fd_sc_hd__conb_1_0/HI LO sky130_fd_sc_hd__conb_1
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__maj3_1 A B C VGND VNB VPB VPWR X
X0 a_109_341# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_265_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_27_47# B a_421_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VGND A a_265_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_27_47# B a_421_341# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_421_341# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_421_47# C VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_27_47# C a_109_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_27_47# C a_109_341# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X12 VPWR A a_265_341# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X13 a_265_341# B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__maj3_2 A B C VGND VNB VPB VPWR X
X0 a_129_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_47_47# C a_129_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 VPWR A a_285_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X3 a_285_369# B a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X4 a_47_47# B a_441_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_441_47# C VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_129_369# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 a_47_47# C a_129_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_47_47# B a_441_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 X a_47_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 X a_47_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_285_47# B a_47_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VGND a_47_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VPWR a_47_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_441_369# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X15 VGND A a_285_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__maj3_4 A B C VGND VNB VPB VPWR X
X0 X a_47_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 X a_47_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_47_297# C a_151_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR a_47_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_47_297# B a_482_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 X a_47_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_151_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_151_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_314_47# B a_47_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_314_297# B a_47_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VGND a_47_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_47_297# C a_151_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VPWR A a_314_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VGND A a_314_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 X a_47_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_47_297# B a_482_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 a_482_297# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 a_482_47# C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 VGND a_47_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 VPWR a_47_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
X0 VPWR S a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_76_199# A0 a_439_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_535_374# a_505_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 VPWR S a_505_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_76_199# A1 a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_218_47# A1 a_76_199# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_218_374# A0 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 X a_76_199# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 X a_76_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VGND S a_218_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VGND S a_505_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_439_47# a_505_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
X0 VGND a_257_199# a_288_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_306_369# A1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 a_288_47# A0 a_79_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_79_21# A1 a_578_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VPWR S a_257_199# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 a_79_21# A0 a_591_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X6 VGND S a_257_199# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_591_369# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X8 a_578_47# S VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VPWR a_257_199# a_306_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X13 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
X0 X a_396_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 X a_396_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VGND a_396_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_206_47# A0 a_396_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_396_47# A1 a_204_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_314_297# A0 a_396_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_490_47# S VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_314_297# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 X a_396_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VGND a_27_47# a_206_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_396_47# A1 a_490_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VGND a_396_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VPWR a_396_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VPWR a_27_47# a_204_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 VPWR a_396_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_27_47# S VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_27_47# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 X a_396_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
X0 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VGND S a_792_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X2 a_1302_47# A0 a_79_21# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X3 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_79_21# A1 a_792_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X5 a_1302_297# A1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_1302_297# a_1259_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VPWR S a_792_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_792_297# A0 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_792_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_792_47# S VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X14 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 VPWR S a_1259_199# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 VGND S a_1259_199# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 a_79_21# A0 a_1302_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X20 a_792_297# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 VGND a_1259_199# a_1302_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X25 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 VPWR a_1259_199# a_1302_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 a_1302_47# a_1259_199# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X28 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X29 a_79_21# A0 a_792_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X30 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X31 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X32 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X33 a_79_21# A1 a_1302_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__mux2i_1 A0 A1 S VGND VNB VPB VPWR Y
X0 a_283_205# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VPWR S a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_27_297# A0 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VGND S a_193_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_204_297# a_283_205# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_27_47# a_283_205# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_283_205# S VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 Y A1 a_204_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 Y A1 a_193_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_27_47# A0 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__mux2i_2 A0 A1 S VGND VNB VPB VPWR Y
X0 a_361_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_193_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 Y A0 a_361_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VGND a_27_47# a_361_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 Y A1 a_361_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 Y A0 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_361_47# A0 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_361_297# A1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_193_47# S VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VGND S a_193_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_193_297# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_193_297# A0 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_27_47# S VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 Y A1 a_193_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_361_297# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_27_47# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 VPWR S a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 VPWR a_27_47# a_361_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__mux2i_4 A0 A1 S VGND VNB VPB VPWR Y
X0 VGND S a_445_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 Y A1 a_445_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VGND a_1191_21# a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 Y A1 a_445_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VPWR a_1191_21# a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND S a_445_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_445_297# A1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_445_297# A1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_109_47# A0 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 Y A1 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_445_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VPWR S a_1191_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_109_297# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VPWR S a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 Y A0 a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_109_297# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 a_109_47# A0 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 Y A0 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 Y A0 a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 VPWR S a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 VGND a_1191_21# a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 Y A1 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 a_445_297# a_1191_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 Y A0 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X24 VPWR a_1191_21# a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 a_109_297# A0 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 a_445_47# S VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 a_445_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 a_109_47# a_1191_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 VGND S a_1191_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 a_109_297# A0 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X31 a_109_47# a_1191_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X32 a_445_297# a_1191_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X33 a_445_47# S VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
X0 a_277_47# S1 a_1478_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_757_363# S0 a_750_97# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_668_97# S0 a_750_97# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_750_97# S1 a_1478_413# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VPWR A2 a_757_363# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_277_47# S0 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_1478_413# a_1290_413# a_277_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_277_47# S0 a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_923_363# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 VPWR a_1478_413# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_27_413# a_247_21# a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 a_668_97# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VGND a_1478_413# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_193_47# a_247_21# a_277_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_247_21# S0 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_27_413# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X16 VPWR A0 a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X17 a_1478_413# a_1290_413# a_750_97# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X18 a_247_21# S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X19 a_750_97# a_247_21# a_923_363# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X20 VPWR S1 a_1290_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X21 VGND A0 a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 VGND A2 a_834_97# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 a_750_97# a_247_21# a_834_97# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 VGND S1 a_1290_413# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
X0 VPWR A1 a_1060_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X1 a_193_47# a_27_47# a_288_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X2 VPWR a_788_316# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_1279_413# A0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X4 VGND a_788_316# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 X a_788_316# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_288_47# S1 a_788_316# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_193_369# S0 a_288_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_372_413# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 a_872_316# a_27_47# a_1281_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X10 a_288_47# a_27_47# a_372_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 VGND A1 a_1064_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VPWR S1 a_600_345# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X13 a_872_316# S0 a_1279_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X14 a_27_47# S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X15 VPWR A2 a_193_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X16 VGND A2 a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_288_47# a_600_345# a_788_316# VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=150000u
X18 a_397_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_27_47# S0 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_1060_369# a_27_47# a_872_316# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X21 VGND S1 a_600_345# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_1281_47# A0 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 X a_788_316# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 a_288_47# S0 a_397_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X25 a_788_316# S1 a_872_316# VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=150000u
X26 a_788_316# a_600_345# a_872_316# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 a_1064_47# S0 a_872_316# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__mux4_4 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
X0 VPWR A1 a_1061_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X1 a_288_47# S1 a_789_316# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_193_47# a_27_47# a_288_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X3 X a_789_316# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_873_316# a_27_47# a_1282_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X5 a_1280_413# A0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X6 VPWR a_789_316# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VGND a_789_316# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VGND A1 a_1065_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_193_369# S0 a_288_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 X a_789_316# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_398_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 X a_789_316# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VGND S1 a_601_345# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_373_413# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X15 a_288_47# S0 a_398_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X16 a_1282_47# A0 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 X a_789_316# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 a_288_47# a_27_47# a_373_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X19 VPWR a_789_316# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 a_789_316# a_601_345# a_873_316# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 a_27_47# S0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X22 VPWR A2 a_193_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X23 VPWR S1 a_601_345# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X24 a_1065_47# S0 a_873_316# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X25 VGND A2 a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 a_27_47# S0 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 a_288_47# a_601_345# a_789_316# VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=150000u
X28 a_1061_369# a_27_47# a_873_316# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X29 a_789_316# S1 a_873_316# VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=150000u
X30 VGND a_789_316# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 a_873_316# S0 a_1280_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VGND B a_113_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_113_47# A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
X0 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
X0 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X28 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X29 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X30 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
X0 a_206_47# a_27_93# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_27_93# A_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VGND B a_206_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_27_93# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 Y a_27_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
X0 a_229_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 Y a_27_93# a_229_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_27_93# A_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_229_47# a_27_93# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_27_93# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VPWR a_27_93# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 Y a_27_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VGND B a_229_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
X0 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VGND B a_215_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_215_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_215_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_215_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VGND B a_215_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 Y a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_215_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_27_47# A_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_27_47# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 Y a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_109_47# B a_193_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VGND C a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_193_47# A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
X0 a_277_47# C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_277_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_27_47# B a_277_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VGND C a_277_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
X0 a_445_47# A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_27_47# B a_445_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_27_47# B a_445_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_445_47# A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VGND C a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_445_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_27_47# C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VGND C a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_27_47# C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 Y A a_445_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 a_445_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 Y A a_445_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
X0 a_53_93# A_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_232_47# B a_316_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_53_93# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_316_47# a_53_93# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VPWR a_53_93# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VGND C a_232_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
X0 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_408_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_218_47# B a_408_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_218_47# C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_27_47# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_408_47# B a_218_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_27_47# A_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 VGND C a_218_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 Y a_27_47# a_408_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
X0 a_633_47# B a_215_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_215_47# B a_633_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_215_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_215_47# B a_633_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VGND C a_633_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_633_47# B a_215_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_633_47# C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 Y a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_633_47# C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 a_215_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 VGND C a_633_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 a_27_47# A_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 a_27_47# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 Y a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
X0 a_277_47# A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_193_47# B a_277_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_109_47# C a_193_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VGND D a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
X0 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_277_47# C a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_27_47# C a_277_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_277_47# B a_471_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VGND D a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_27_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 Y A a_471_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_471_47# A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_471_47# B a_277_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_803_47# B a_445_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_27_47# C a_445_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_27_47# C a_445_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_803_47# B a_445_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 Y A a_803_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND D a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_445_47# C a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_27_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 Y A a_803_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 VGND D a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_27_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_803_47# A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X24 a_803_47# A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X28 a_445_47# B a_803_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 a_445_47# C a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X31 a_445_47# B a_803_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
X0 Y a_41_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_232_47# C a_316_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_423_47# a_41_93# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_41_93# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_316_47# B a_423_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_41_93# A_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VGND D a_232_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
X0 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_215_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_465_47# B a_215_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_27_47# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_215_47# B a_465_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_655_47# C a_465_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VGND D a_655_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_27_47# A_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_465_47# C a_655_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 Y a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_655_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
X0 a_633_47# B a_215_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VGND D a_991_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_215_47# B a_633_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_215_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_215_47# B a_633_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_991_47# C a_633_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_991_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 a_633_47# B a_215_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_633_47# C a_991_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 VGND D a_991_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 Y a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 a_633_47# C a_991_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 a_215_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 a_991_47# C a_633_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 a_27_47# A_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X29 a_27_47# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X30 Y a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X32 a_991_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X33 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nand4bb_1 A_N B_N C D VGND VNB VPB VPWR Y
X0 Y a_496_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_426_47# a_496_21# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VPWR A_N a_496_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 VGND A_N a_496_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_27_93# B_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_326_47# a_27_93# a_426_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_27_93# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VPWR a_27_93# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VGND D a_218_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_218_47# C a_326_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nand4bb_2 A_N B_N C D VGND VNB VPB VPWR Y
X0 a_341_47# a_27_47# a_591_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_781_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 Y a_193_47# a_341_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VGND D a_781_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_341_47# a_193_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 Y a_193_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_27_47# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 VPWR a_193_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VPWR A_N a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X13 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 VGND A_N a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_27_47# B_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_591_47# a_27_47# a_341_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 a_591_47# C a_781_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_781_47# C a_591_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nand4bb_4 A_N B_N C D VGND VNB VPB VPWR Y
X0 a_1266_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_432_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_432_47# a_193_47# a_850_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 Y a_193_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VGND D a_1266_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VPWR a_193_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_432_47# a_193_47# a_850_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_1266_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 Y a_193_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 Y a_27_47# a_432_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_850_47# a_193_47# a_432_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 VPWR a_193_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 a_432_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 a_850_47# C a_1266_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 VGND D a_1266_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 a_850_47# C a_1266_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 VGND B_N a_193_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 a_27_47# A_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 a_1266_47# C a_850_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X29 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X30 a_1266_47# C a_850_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 a_27_47# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X32 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X33 VPWR B_N a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X34 Y a_27_47# a_432_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X35 a_850_47# a_193_47# a_432_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
X0 a_109_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 Y B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
X0 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
X0 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
X0 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X24 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X28 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X29 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
X0 a_74_47# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 Y a_74_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_74_47# B_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VPWR A a_265_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_265_297# a_74_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
X0 Y a_251_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 Y a_251_21# a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VGND a_251_21# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_27_297# a_251_21# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_251_21# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_251_21# B_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
X0 a_27_297# a_419_21# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 Y a_419_21# a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 Y a_419_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_27_297# a_419_21# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 Y a_419_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_419_21# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 Y a_419_21# a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_419_21# B_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VGND a_419_21# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 VGND a_419_21# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_193_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 Y C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 Y C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_109_297# B a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
X0 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 Y C a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_281_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_27_297# B a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 Y C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_281_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 VGND C Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
X0 a_27_297# B a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_449_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_449_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 Y C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VGND C Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_449_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 Y C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_27_297# B a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 Y C a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 Y C a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 a_449_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 VGND C Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VPWR C_N a_91_199# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_161_297# B a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VGND C_N a_91_199# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 Y a_91_199# a_161_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_245_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 Y a_91_199# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
X0 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_281_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_27_297# B a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 Y a_531_21# a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_281_297# a_531_21# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 Y a_531_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_531_21# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VGND a_531_21# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_531_21# C_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
X0 a_197_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_197_297# B a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VPWR A a_197_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR A a_197_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_555_297# B a_197_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_555_297# a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_197_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_197_297# B a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 Y a_27_47# a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_27_47# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_27_47# C_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 VGND a_27_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 VGND a_27_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 a_555_297# B a_197_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 Y a_27_47# a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 Y a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 a_555_297# a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 Y a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
X0 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_191_297# B a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_297_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 Y C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VGND D Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_109_297# C a_191_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 Y D a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
X0 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_281_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_27_297# B a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_281_297# C a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_475_297# C a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 Y D VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 Y C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VGND C Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_475_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 VGND D Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 Y D a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
X0 a_27_297# B a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_807_297# C a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_449_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_449_297# C a_807_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 Y D a_807_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 Y D a_807_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 Y D VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_807_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_807_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VGND D Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 Y C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 a_27_297# B a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 Y C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 a_449_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X24 Y D VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 a_807_297# C a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 VGND C Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 VGND D Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 a_449_297# C a_807_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X30 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 VGND C Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
X0 VPWR D_N a_91_199# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 VGND D_N a_91_199# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_161_297# C a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_245_297# B a_341_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 Y a_91_199# a_161_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 Y C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_341_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND a_91_199# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
X0 a_277_297# C a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 Y a_694_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VGND a_694_21# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 Y a_694_21# a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND C Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_474_297# a_694_21# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_694_21# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_27_297# B a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_474_297# C a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 Y C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_277_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 a_694_21# D_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
X0 Y a_1191_21# a_803_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VGND C Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VGND a_1191_21# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_803_297# a_1191_21# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VGND C Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_445_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_445_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_27_297# B a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 Y a_1191_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_445_297# C a_803_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_803_297# C a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_1191_21# D_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 a_1191_21# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 a_445_297# C a_803_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 a_803_297# C a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 VGND a_1191_21# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 a_27_297# B a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 a_803_297# a_1191_21# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X28 Y C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 Y a_1191_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X32 Y a_1191_21# a_803_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X33 Y C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nor4bb_1 A B C_N D_N VGND VNB VPB VPWR Y
X0 VGND a_205_93# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_573_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_27_410# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_393_297# a_27_410# a_477_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_477_297# B a_573_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 Y a_205_93# a_393_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VGND D_N a_205_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VPWR D_N a_205_93# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 Y a_27_410# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_27_410# C_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nor4bb_2 A B C_N D_N VGND VNB VPB VPWR Y
X0 a_776_297# B a_418_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_336_297# a_201_93# a_418_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_336_297# a_27_410# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_27_410# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 VGND a_201_93# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR A a_776_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_418_297# a_201_93# a_336_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 Y a_27_410# a_336_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 Y a_27_410# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VGND a_27_410# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VPWR C_N a_201_93# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 a_776_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 Y a_201_93# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 VGND C_N a_201_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_27_410# D_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_418_297# B a_776_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nor4bb_4 A B C_N D_N VGND VNB VPB VPWR Y
X0 a_729_297# B a_1087_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VGND a_197_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VPWR D_N a_197_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 Y a_197_47# a_311_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 Y a_197_47# a_311_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VGND a_27_297# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VPWR A a_1087_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_27_297# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VPWR A a_1087_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_311_297# a_197_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_27_297# C_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_311_297# a_197_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 Y a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 a_1087_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 Y a_197_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 a_1087_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 a_729_297# B a_1087_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 VGND D_N a_197_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 VGND a_197_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 a_311_297# a_27_297# a_729_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 a_311_297# a_27_297# a_729_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 VGND a_27_297# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 a_729_297# a_27_297# a_311_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X30 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 a_729_297# a_27_297# a_311_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X32 a_1087_297# B a_729_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X33 a_1087_297# B a_729_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X34 Y a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X35 Y a_197_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 a_76_199# a_206_369# a_489_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VPWR a_206_369# a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 VPWR A1_N a_206_369# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_206_369# A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 VGND B1 a_489_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 X a_76_199# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_489_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 X a_76_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_205_47# A2_N a_206_369# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_76_199# B2 a_585_369# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_585_369# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 VGND A1_N a_205_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 VPWR A1_N a_295_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X1 a_295_369# A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 a_581_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VGND a_84_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_294_47# A2_N a_295_369# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VGND A1_N a_294_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 X a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_84_21# a_295_369# a_581_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 X a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VPWR a_295_369# a_84_21# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X10 VPWR a_84_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_665_369# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X12 a_84_21# B2 a_665_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X13 VGND B1 a_581_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 a_415_21# A2_N a_717_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VGND a_193_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_27_47# a_415_21# a_193_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR a_193_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VGND a_193_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_193_297# a_415_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_717_47# A2_N a_415_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VGND B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_193_297# a_415_21# a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 X a_193_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VGND A1_N a_717_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VPWR a_193_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_415_21# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 VPWR A1_N a_415_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 a_27_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 VPWR A2_N a_415_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 VPWR a_415_21# a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 VPWR B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 a_109_297# B2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 a_717_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 a_415_21# A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X24 X a_193_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 a_109_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 X a_193_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 X a_193_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
X0 a_112_297# A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 Y B2 a_478_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VGND B1 a_394_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR A1_N a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VPWR a_112_297# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_478_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_112_47# A2_N a_112_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_394_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VGND A1_N a_112_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 Y a_112_297# a_394_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
X0 a_113_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VGND B2 a_471_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_113_297# A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_113_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_113_297# A2_N a_113_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VPWR A2_N a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VPWR A1_N a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VGND A1_N a_113_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 Y a_113_297# a_471_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VPWR B1 a_730_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_113_47# A2_N a_113_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_471_47# a_113_297# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VGND B1 a_471_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 Y a_113_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 Y B2 a_730_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_471_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VPWR a_113_297# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 a_730_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 a_730_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_471_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
X0 VPWR A1_N a_113_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VGND B2 a_807_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VGND B1 a_807_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_113_47# A2_N a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_113_47# A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_113_47# A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_807_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_113_47# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_27_47# A2_N a_113_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_1241_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VPWR A2_N a_113_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 Y B2 a_1241_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VPWR A2_N a_113_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 Y a_113_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 Y B2 a_1241_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_807_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_27_47# A2_N a_113_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 a_807_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 VPWR B1 a_1241_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_1241_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 VPWR a_113_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 a_1241_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 VGND A1_N a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 Y a_113_47# a_807_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 VGND B2 a_807_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 VPWR A1_N a_113_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 a_113_47# A2_N a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 VGND A1_N a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 Y a_113_47# a_807_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 Y a_113_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X30 a_807_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 a_113_47# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X32 VPWR a_113_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X33 a_1241_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X34 a_27_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X35 a_807_47# a_113_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X36 VPWR B1 a_1241_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X37 a_27_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X38 a_807_47# a_113_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X39 VGND B1 a_807_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
X0 a_382_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VGND A1 a_297_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_79_21# B1 a_297_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_297_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_79_21# A2 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
X0 a_384_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_470_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VGND A1 a_384_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_79_21# A2 a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_79_21# B1 a_384_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
X0 a_80_21# A2 a_934_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 X a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VGND A1 a_475_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 X a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_475_47# B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_80_21# B1 a_475_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_80_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 X a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_475_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VPWR B1 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_762_297# A2 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 X a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 VPWR A1 a_762_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 a_934_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 VGND A2 a_475_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 a_475_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o21ai_0 A1 A2 B1 VGND VNB VPB VPWR Y
X0 VGND A2 a_32_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 a_32_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_32_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VPWR A1 a_120_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 a_120_369# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
X0 a_109_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=700000u l=150000u
X2 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VPWR A1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
X0 a_112_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VGND A2 a_29_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VPWR A1 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_29_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VGND A1 a_29_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 Y A2 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_112_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_29_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_29_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 Y B1 a_29_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
X0 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VGND A1 a_32_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 Y B1 a_32_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 Y B1 a_32_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_32_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_32_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND A2 a_32_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_32_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 a_32_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 VGND A2 a_32_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 a_32_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 VGND A1 a_32_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 a_32_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
X0 a_448_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VPWR B1_N a_222_93# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_79_199# a_222_93# a_448_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VGND B1_N a_222_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VGND A1 a_448_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_544_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 X a_79_199# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 X a_79_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VPWR a_222_93# a_79_199# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_79_199# A2 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
X0 X a_174_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VGND a_174_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VPWR a_27_93# a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_174_21# A2 a_574_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_574_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_27_93# B1_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_174_21# a_27_93# a_478_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VGND A1 a_478_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_478_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VPWR a_174_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_27_93# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 X a_174_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
X0 a_575_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VGND a_187_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_27_297# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VPWR A1 a_743_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_187_21# a_27_297# a_575_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VGND A2 a_575_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 X a_187_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_187_21# A2 a_743_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 X a_187_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VGND A1 a_575_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_187_21# a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_575_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VPWR a_187_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VPWR a_187_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_743_297# A2 a_187_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 VGND a_187_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_575_47# a_27_297# a_187_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 a_743_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 VPWR a_27_297# a_187_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 X a_187_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 X a_187_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 a_27_297# B1_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 VGND A1 a_297_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 Y a_105_352# a_297_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VPWR a_105_352# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_297_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_388_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND B1_N a_105_352# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_105_352# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 Y A2 a_388_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 Y a_28_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VGND B1_N a_28_297# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_28_297# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_397_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_397_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_229_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 Y A2 a_397_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 Y a_28_297# a_229_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VGND A1 a_229_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VPWR A1 a_397_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_229_47# a_28_297# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VPWR a_28_297# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_229_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VGND A2 a_229_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 a_225_47# a_33_297# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_225_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_561_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_561_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VPWR A1 a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND A2 a_225_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR A1 a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 Y a_33_297# a_225_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VGND A1 a_225_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_561_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_225_47# a_33_297# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 Y a_33_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 Y A2 a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 Y a_33_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 Y A2 a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 VGND B1_N a_33_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_33_297# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 VPWR a_33_297# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 Y a_33_297# a_225_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 VPWR a_33_297# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 a_561_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 a_225_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 a_225_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 VGND A2 a_225_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 VGND A1 a_225_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 a_225_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 VPWR B1 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_215_47# B1 a_78_199# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 X a_78_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_292_297# B2 a_78_199# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VGND A1 a_215_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_215_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_78_199# A2 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_493_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 X a_78_199# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_78_199# B2 a_215_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 X a_81_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_81_21# B2 a_301_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 X a_81_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_301_47# B1 a_81_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_81_21# A2 a_579_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VPWR B1 a_383_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_383_297# B2 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND A1 a_301_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_301_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_579_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 a_96_21# A2 a_918_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 X a_96_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_566_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_484_47# B1 a_96_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VGND a_96_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VPWR a_96_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_918_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VGND A2 a_484_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 X a_96_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VPWR a_96_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VPWR A1 a_918_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 X a_96_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VGND a_96_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VGND A1 a_484_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_918_297# A2 a_96_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_484_47# B2 a_96_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_484_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 VPWR B1 a_566_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 a_484_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 a_96_21# B2 a_566_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 a_96_21# B2 a_484_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 a_566_297# B2 a_96_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 a_96_21# B1 a_484_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 X a_96_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
X0 Y A2 a_307_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_307_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_109_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 Y B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
X0 Y B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 Y A2 a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_475_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_475_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 VPWR A1 a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
X0 a_797_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_33_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_33_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_33_47# B2 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_33_47# B2 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 Y B1 a_33_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 Y B2 a_797_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_33_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 VPWR B1 a_797_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 VGND A2 a_33_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VPWR B1 a_797_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 Y B2 a_33_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 Y B2 a_33_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 a_33_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_33_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 a_797_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 a_797_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X24 a_797_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 Y B2 a_797_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 a_33_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X28 VGND A1 a_33_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 VGND A1 a_33_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 VGND A2 a_33_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 Y B1 a_33_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 a_253_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VPWR A1 a_253_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 X a_103_199# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 X a_103_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VGND A1 a_253_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_103_199# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_253_47# B1 a_103_199# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VGND A3 a_253_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_253_297# A2 a_337_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_337_297# A3 a_103_199# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 a_430_297# A3 a_108_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 X a_108_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_108_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VGND A1 a_346_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_346_47# B1 a_108_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VGND A3 a_346_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VGND a_108_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VPWR a_108_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VPWR A1 a_346_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 X a_108_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_346_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_346_297# A2 a_430_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 VPWR a_102_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_496_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_496_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR B1 a_102_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_926_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND a_102_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 X a_102_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VPWR a_102_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND a_102_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_672_297# A3 a_102_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_102_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 X a_102_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 X a_102_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_102_21# A3 a_672_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_926_297# A2 a_672_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 VGND A1 a_496_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VGND A3 a_496_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 VPWR A1 a_926_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 a_102_21# B1 a_496_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 a_496_47# B1 a_102_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 VGND A2 a_496_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 a_672_297# A2 a_926_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 X a_102_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 a_496_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
X0 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VGND A3 a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_109_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_109_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_193_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND A1 a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR A1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_109_297# A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
X0 a_281_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_281_297# A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_27_297# A2 a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 Y A3 a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
X0 a_27_297# A2 a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VGND A1 a_31_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_449_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 Y B1 a_31_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VGND A3 a_31_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_449_297# A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_31_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 Y A3 a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_449_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_31_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_31_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 Y A3 a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 VGND A2 a_31_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 a_31_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_27_297# A2 a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 VGND A1 a_31_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 VGND A2 a_31_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X24 a_31_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 Y B1 a_31_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 VGND A3 a_31_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 a_449_297# A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X29 a_31_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 a_31_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 a_31_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 X a_77_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VPWR A1 a_227_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_77_199# B1 a_227_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_227_297# A2 a_323_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_77_199# B2 a_539_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND A3 a_227_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 X a_77_199# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_227_47# B2 a_77_199# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_227_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_323_297# A3 a_77_199# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_539_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 VGND A1 a_227_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 a_429_297# A3 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_345_47# B2 a_79_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_79_21# B1 a_345_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_79_21# B2 a_629_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VGND A1 a_345_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VPWR A1 a_345_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_629_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_345_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VGND A3 a_345_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_345_297# A2 a_429_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 VPWR a_549_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VGND a_549_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 X a_549_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_277_297# A3 a_549_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_739_297# B2 a_549_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR B1 a_739_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_549_297# A3 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_549_297# B2 a_739_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 X a_549_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_739_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_549_297# B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VGND a_549_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_27_47# B1 a_549_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 X a_549_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 a_27_297# A2 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_549_297# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 X a_549_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 a_277_297# A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 a_27_47# B2 a_549_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 VPWR a_549_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
X0 a_109_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_461_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_333_297# A2 a_461_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 Y B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 Y A3 a_333_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VPWR B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o32ai_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
X0 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_729_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 Y A3 a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_475_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VPWR A1 a_729_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_475_297# A2 a_729_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 Y B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_729_297# A2 a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
X0 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 Y A3 a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_1224_297# A2 a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_1224_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_1224_297# A2 a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_806_297# A2 a_1224_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 Y B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_806_297# A2 a_1224_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_1224_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 a_806_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 VPWR A1 a_1224_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 Y B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X29 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 VPWR A1 a_1224_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X31 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X32 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X33 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X34 Y A3 a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X35 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X36 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X37 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X38 a_806_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X39 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
X0 a_393_297# A3 a_511_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_321_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_321_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR B1 a_103_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VGND A1 a_321_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_103_21# A4 a_393_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_103_21# B1 a_321_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 X a_103_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_619_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_511_297# A2 a_619_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 X a_103_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VGND A3 a_321_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
X0 a_496_297# A3 a_597_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_79_21# B1 a_393_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_597_297# A2 a_697_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VGND A3 a_393_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_697_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VGND A1 a_393_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_79_21# A4 a_496_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_393_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_393_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
X0 a_639_297# A3 a_889_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_889_297# A2 a_1083_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_467_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_79_21# A4 a_639_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_889_297# A3 a_639_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_79_21# B1 a_467_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_639_297# A4 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_467_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VGND A1 a_467_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VGND A3 a_467_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_467_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VPWR A1 a_1083_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_467_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VGND A2 a_467_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 a_1083_297# A2 a_889_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 a_467_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 a_1083_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 VGND A4 a_467_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o41ai_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
X0 a_432_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_109_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VGND A3 a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_109_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_193_297# A3 a_348_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 Y B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VGND A1 a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 Y A4 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_348_297# A2 a_432_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o41ai_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
X0 a_549_297# A2 a_743_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_299_297# A3 a_549_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 Y A4 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_549_297# A3 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_299_297# A4 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_27_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VPWR A1 a_743_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_743_297# A2 a_549_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 VGND A4 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 a_743_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
X0 VPWR A1 a_1243_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VGND A4 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VGND A4 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_467_297# A4 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 Y A4 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_885_297# A2 a_1243_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_885_297# A2 a_1243_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_885_297# A3 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 VPWR A1 a_1243_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 a_1243_297# A2 a_885_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 a_27_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 a_467_297# A3 a_885_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_1243_297# A2 a_885_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 a_27_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 a_1243_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 a_885_297# A3 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X29 a_467_297# A4 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X30 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 a_467_297# A3 a_885_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X32 a_1243_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X33 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X34 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X35 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X36 Y A4 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X37 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X38 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X39 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 VPWR C1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_215_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_215_47# B1 a_510_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_297_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VPWR A1 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND A2 a_215_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_510_47# C1 a_79_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 VPWR B1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_27_47# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_110_47# B1 a_182_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_27_47# C1 a_110_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_27_47# A2 a_373_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_373_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VGND A2 a_182_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_182_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_557_47# C1 a_79_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_474_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_950_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_79_21# C1 a_748_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_748_47# B1 a_474_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND A1 a_474_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_474_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VPWR A1 a_950_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 VGND A2 a_474_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VPWR C1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 a_79_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 a_1122_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 a_79_21# A2 a_1122_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 a_474_47# B1 a_557_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
X0 a_110_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VPWR A1 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_326_47# C1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_27_47# B1 a_326_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
X0 Y A2 a_487_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_27_47# C1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_487_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_487_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 Y C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND A2 a_286_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_27_47# B1 a_286_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_286_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_286_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VPWR A1 a_487_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_286_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 VGND A1 a_286_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
X0 a_27_47# B1 a_978_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 Y C1 a_1314_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_110_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 Y C1 a_806_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VPWR A1 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_978_47# C1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_110_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 Y A2 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 VPWR A1 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 a_110_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 Y A2 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 a_27_47# B1 a_806_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 a_806_47# C1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 a_1314_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 a_806_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 a_110_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X29 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 a_51_297# A2 a_512_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_512_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VPWR a_51_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VGND a_51_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_149_47# B1 a_240_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_51_297# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VPWR B1 a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_240_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_240_47# B2 a_149_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VGND A2 a_240_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_245_297# B2 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_51_297# C1 a_149_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 VGND a_38_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_225_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_38_47# C1 a_141_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_225_47# B2 a_141_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VGND A2 a_225_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_141_47# B1 a_225_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_237_297# B2 a_38_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VPWR B1 a_237_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 X a_38_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_38_47# A2 a_497_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_497_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 VPWR a_38_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 X a_38_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_38_47# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 VGND A2 a_277_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_27_47# B2 a_277_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_277_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_277_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_277_47# B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_277_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VGND A1 a_277_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_27_47# B1 a_277_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_717_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_109_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 VPWR B1 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 VPWR A1 a_717_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 a_27_47# C1 a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 a_109_47# A2 a_717_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_109_47# B2 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 VPWR C1 a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 a_109_47# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 a_277_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 a_717_297# A2 a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X24 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 a_277_297# B2 a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
X0 VPWR B1 a_295_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VGND A1 a_213_123# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_213_123# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 Y A2 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_493_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_109_47# B2 a_213_123# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 Y C1 a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_295_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_213_123# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
X0 a_734_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_300_47# B2 a_28_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_734_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 Y A2 a_734_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_28_47# C1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_382_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 Y C1 a_28_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_28_47# B2 a_300_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VGND A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_382_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 VPWR B1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_300_47# B1 a_28_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 Y B2 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_300_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VPWR A1 a_734_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 a_28_47# B1 a_300_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 VGND A2 a_300_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
X0 Y B2 a_553_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 Y C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_27_47# B1 a_471_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VGND A2 a_471_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_471_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_553_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VPWR A1 a_1241_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_553_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_27_47# C1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_471_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_471_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 VPWR B1 a_553_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 a_27_47# C1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 Y A2 a_1241_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 Y A2 a_1241_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_471_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_471_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 VPWR A1 a_1241_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 a_27_47# B2 a_471_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 a_1241_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X24 a_1241_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 Y C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 a_27_47# B1 a_471_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 VGND A2 a_471_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 VGND A1 a_471_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 a_553_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X30 a_1241_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X31 VPWR B1 a_553_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X32 VGND A1 a_471_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X33 Y B2 a_553_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X34 a_1241_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X35 a_471_47# B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X36 a_553_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X37 a_471_47# B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X38 a_471_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X39 a_27_47# B2 a_471_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 a_266_47# B1 a_585_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VGND A1 a_266_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VPWR C1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_266_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 X a_81_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND A3 a_266_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_266_297# A2 a_368_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_81_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_585_47# C1 a_81_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_368_297# A3 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VPWR A1 a_266_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 X a_81_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 VPWR a_91_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_360_297# A2 a_460_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_360_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_91_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_460_297# A3 a_91_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_360_47# B1 a_677_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VGND A3 a_360_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VGND A1 a_360_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VPWR C1 a_91_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 X a_91_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VGND a_91_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VPWR A1 a_360_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_677_47# C1 a_91_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 X a_91_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 a_79_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VPWR C1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_717_47# B1 a_467_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_79_21# C1 a_467_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_717_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VGND A2 a_717_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VGND A3 a_717_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_1147_297# A2 a_875_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_1147_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_467_47# B1 a_717_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_467_47# C1 a_79_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_875_297# A2 a_1147_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 VPWR A1 a_1147_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 a_79_21# A3 a_875_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 a_717_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 a_717_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 a_875_297# A3 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X24 VGND A1 a_717_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o311ai_0 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
X0 a_138_47# B1 a_458_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VPWR A1 a_138_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 VGND A3 a_138_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VGND A1 a_138_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_458_47# C1 Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_138_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 a_222_369# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X8 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 a_138_369# A2 a_222_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
X0 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_138_47# B1 a_458_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_222_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_138_297# A2 a_222_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VGND A3 a_138_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VGND A1 a_138_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_458_47# C1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_138_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VPWR A1 a_138_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
X0 a_55_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_301_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 Y C1 a_729_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_51_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 Y A3 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_729_47# C1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_729_47# B1 a_55_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VGND A3 a_55_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 VGND A2 a_55_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_55_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VPWR A1 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_301_297# A2 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 a_55_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 VGND A1 a_55_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 a_55_47# B1 a_729_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 a_51_297# A2 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
X0 VPWR A1 a_39_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_125_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_461_297# A2 a_39_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_461_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VGND A2 a_125_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_125_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_39_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_39_297# A2 a_461_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 Y A3 a_461_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VGND A3 a_125_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 Y C1 a_1163_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_39_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_125_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_1163_47# C1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 VGND A1 a_125_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 a_39_297# A2 a_461_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_125_47# B1 a_1163_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 a_125_47# B1 a_1163_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X24 a_461_297# A2 a_39_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 VGND A1 a_125_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 Y A3 a_461_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X28 Y C1 a_1163_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 a_125_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 a_125_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 a_125_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X32 a_461_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X33 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X34 a_1163_47# B1 a_125_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X35 a_1163_47# C1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X36 a_1163_47# B1 a_125_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X37 VGND A2 a_125_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X38 VGND A3 a_125_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X39 VPWR A1 a_39_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
X0 VPWR D1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_306_47# C1 a_409_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VGND A1 a_512_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_79_21# D1 a_306_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_512_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_79_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_79_21# A2 a_676_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_676_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_409_47# B1 a_512_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
X0 a_386_47# C1 a_458_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 X a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_458_47# B1 a_566_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_566_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VGND A1 a_566_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_80_21# D1 a_386_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_674_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_80_21# A2 a_674_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VPWR B1 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_80_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VPWR D1 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 X a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
X0 VGND A2 a_361_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_681_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_361_47# B1 a_445_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_361_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VPWR C1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_27_297# A2 a_681_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_445_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_277_47# B1 a_361_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VPWR A1 a_852_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_27_47# C1 a_277_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_852_297# A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 a_27_297# D1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 a_27_297# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_27_47# D1 a_27_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 a_27_297# D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 VGND A1 a_361_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 VPWR D1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 a_361_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
X0 a_235_47# B1 a_343_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_343_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VGND A1 a_343_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 Y D1 a_163_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_454_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 Y A2 a_454_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_163_47# C1 a_235_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
X0 Y A2 a_664_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_664_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VPWR A1 a_664_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_497_47# B1 a_298_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_497_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_27_47# D1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VGND A1 a_497_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_298_47# B1 a_497_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_497_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 Y D1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VGND A2 a_497_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 a_664_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 a_27_47# C1 a_298_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 a_298_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
X0 a_803_47# B1 a_445_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_27_47# C1 a_445_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_27_47# C1 a_445_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_803_47# B1 a_445_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VPWR A1 a_1163_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VGND A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 Y D1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_1163_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_1163_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_445_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_1163_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 a_803_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 VPWR A1 a_1163_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 VGND A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 VGND A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 Y A2 a_1163_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 VGND A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X24 a_27_47# D1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 a_803_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 Y A2 a_1163_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 a_803_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 Y D1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X30 a_27_47# D1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X32 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X33 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X34 a_445_47# B1 a_803_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X35 a_803_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X36 a_445_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X37 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X38 a_1163_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X39 a_445_47# B1 a_803_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__or2_0 A B VGND VNB VPB VPWR X
X0 VGND a_68_355# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_150_355# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 VGND B a_68_355# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_68_355# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_68_355# B a_150_355# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 VPWR a_68_355# X VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
X0 a_150_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 VGND a_68_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VGND B a_68_297# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_68_297# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_68_297# B a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 VPWR a_68_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
X0 a_39_297# B a_121_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 X a_39_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VGND a_39_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR a_39_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_39_297# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VGND B a_39_297# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_121_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 X a_39_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
X0 a_35_297# B a_121_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 X a_35_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 X a_35_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VPWR a_35_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VPWR a_35_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 X a_35_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_35_297# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VGND B a_35_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_121_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 X a_35_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
X0 a_219_297# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_27_53# B_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VGND a_27_53# a_219_297# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VGND a_219_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_219_297# a_27_53# a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_301_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 VPWR B_N a_27_53# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VPWR a_219_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
X0 VGND a_218_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_218_297# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_27_53# B_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_218_297# a_27_53# a_300_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_300_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 X a_218_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VPWR B_N a_27_53# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 X a_218_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VPWR a_218_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VGND a_27_53# a_218_297# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
X0 X a_219_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_219_297# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VGND a_219_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 X a_219_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_27_53# B_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 X a_219_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR B_N a_27_53# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VPWR a_219_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND a_219_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_219_297# a_27_53# a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_301_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 VGND a_27_53# a_219_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 X a_219_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VPWR a_219_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
X0 VPWR a_29_53# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_111_297# B a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_29_53# C a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 VGND a_29_53# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_29_53# C VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_29_53# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_183_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VGND B a_29_53# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
X0 VPWR a_30_53# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_112_297# B a_184_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_184_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 X a_30_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_30_53# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_30_53# C a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_30_53# C VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 X a_30_53# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VGND B a_30_53# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VGND a_30_53# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
X0 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_193_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_27_47# C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_27_47# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_109_297# B a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
X0 a_215_53# a_109_93# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VGND a_215_53# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_215_53# a_109_93# a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_297_297# B a_369_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_369_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 VPWR a_215_53# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_215_53# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VGND C_N a_109_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VGND B a_215_53# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VPWR C_N a_109_93# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
X0 VGND a_27_47# a_176_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_176_21# B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_27_47# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 VGND A a_176_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_27_47# C_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VPWR A a_388_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 a_472_297# a_27_47# a_176_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_388_297# B a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
X0 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_542_297# B a_626_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_626_297# a_27_47# a_176_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_27_47# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VGND A a_176_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_27_47# C_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 VGND a_27_47# a_176_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VPWR A a_542_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_176_21# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
X0 a_27_297# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VGND D a_27_297# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VGND B a_27_297# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_109_297# C a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_205_297# B a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_27_297# C VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_277_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_27_297# D a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
X0 a_27_297# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VGND D a_27_297# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VGND B a_27_297# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_109_297# C a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_205_297# B a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_27_297# C VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_277_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_27_297# D a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
X0 a_32_297# C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_114_297# C a_220_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VGND D a_32_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 X a_32_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_32_297# D a_114_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND a_32_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 X a_32_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 X a_32_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VPWR a_32_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VPWR a_32_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_32_297# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_304_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 X a_32_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VGND B a_32_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_220_297# B a_304_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 VGND a_32_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
X0 VGND a_109_53# a_215_297# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_215_297# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VGND B a_215_297# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_297_297# C a_392_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_215_297# a_109_53# a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_392_297# B a_465_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 VGND a_215_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VGND D_N a_109_53# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_215_297# C VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VPWR D_N a_109_53# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_465_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 VPWR a_215_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
X0 a_176_21# a_27_53# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_27_53# D_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VGND C a_176_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_176_21# B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VPWR A a_387_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_387_297# B a_483_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_483_297# C a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_27_53# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 a_555_297# a_27_53# a_176_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X12 VGND A a_176_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
X0 a_403_297# B a_487_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_297_297# C a_403_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_487_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND a_109_93# a_215_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VGND a_215_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_215_297# a_109_93# a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_215_297# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VGND D_N a_109_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VPWR D_N a_109_93# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 VPWR a_215_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VPWR a_215_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VGND B a_215_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VGND a_215_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 a_215_297# C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
X0 VGND a_205_93# a_311_413# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_393_413# a_27_410# a_489_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_311_413# a_205_93# a_393_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_27_410# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_27_410# C_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_489_297# B a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_561_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VPWR a_311_413# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_311_413# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VGND B a_311_413# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VGND D_N a_205_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VPWR D_N a_205_93# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X12 a_311_413# a_27_410# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 VGND a_311_413# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
X0 VPWR a_316_413# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VGND a_316_413# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_27_410# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 VGND B a_316_413# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_316_413# a_27_410# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_316_413# a_206_93# a_398_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 VGND D_N a_206_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_398_413# a_27_410# a_494_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_494_297# B a_566_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 VGND a_206_93# a_316_413# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VPWR D_N a_206_93# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 a_316_413# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_566_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X13 X a_316_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_27_410# C_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 X a_316_413# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
X0 X a_315_380# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_499_297# B a_583_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VGND a_205_93# a_315_380# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 X a_315_380# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VGND a_315_380# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_27_410# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_27_410# C_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_315_380# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_315_380# a_205_93# a_397_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 X a_315_380# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VGND B a_315_380# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VGND a_315_380# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VPWR a_315_380# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VGND D_N a_205_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 VPWR a_315_380# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 VPWR D_N a_205_93# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X16 a_397_297# a_27_410# a_499_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 a_583_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 X a_315_380# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 a_315_380# a_27_410# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__probe_p_8 A VGND VNB VPB VPWR X
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__probec_p_8 A VGND VNB VPB VPWR X
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__sdfbbn_1 CLK_N D RESET_B SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
X0 VPWR SET_B a_1102_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_1800_413# a_1887_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 VGND a_1102_21# a_1614_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X3 a_2596_47# a_1887_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X4 a_1351_329# a_1396_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X5 a_1887_21# a_1714_47# a_2122_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X6 a_2122_329# a_1396_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X7 VGND a_1887_21# Q_N VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_1822_47# a_1887_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_917_47# a_193_47# a_1017_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_1017_413# a_1102_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 VGND SET_B a_1241_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_1102_21# a_917_47# a_1351_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X13 VGND a_423_315# a_735_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 VPWR a_1102_21# a_1572_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X15 a_917_47# a_27_47# a_1030_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X16 VPWR SCD a_381_363# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X17 a_381_363# a_423_315# a_453_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 a_1030_47# a_1102_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_1887_21# a_1396_21# a_2004_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X20 a_381_47# SCE a_453_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 a_735_47# D a_453_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_1572_329# a_193_47# a_1714_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X23 VPWR a_1887_21# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X24 a_2596_47# a_1887_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 a_423_315# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 a_2004_47# a_1714_47# a_1887_21# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X27 a_1396_21# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 a_1241_47# a_917_47# a_1102_21# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X29 a_1714_47# a_27_47# a_1800_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X30 VGND a_2596_47# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 a_1396_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X32 a_423_315# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X33 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 a_1614_47# a_27_47# a_1714_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X35 a_27_47# CLK_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X36 a_27_47# CLK_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X37 a_752_413# D a_453_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X38 a_1714_47# a_193_47# a_1822_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X39 VPWR a_2596_47# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X40 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X41 a_453_47# a_27_47# a_917_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X42 VGND SCD a_381_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X43 a_453_47# a_193_47# a_917_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X44 VPWR SCE a_752_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X45 VPWR SET_B a_1887_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X46 a_1102_21# a_1396_21# a_1241_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X47 VGND SET_B a_2004_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__sdfbbn_2 CLK_N D RESET_B SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
X0 VGND a_423_315# a_764_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VPWR a_2696_47# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VPWR SET_B a_1107_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_423_315# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_1800_413# a_1888_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 VGND SET_B a_1251_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_1351_329# a_1401_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X7 a_1251_47# a_931_47# a_1107_21# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X8 a_1888_21# a_1714_47# a_2122_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X9 a_2122_329# a_1401_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X10 a_1888_21# a_1401_21# a_2004_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X11 VGND a_1888_21# Q_N VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_2696_47# a_1888_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 Q a_2696_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_931_47# a_193_47# a_1017_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 a_1017_413# a_1107_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X16 a_1107_21# a_931_47# a_1351_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X17 a_2696_47# a_1888_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 a_2004_47# a_1714_47# a_1888_21# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X19 VPWR a_1107_21# a_1572_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X20 VGND a_2696_47# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 VPWR SCD a_381_363# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X22 a_381_363# a_423_315# a_453_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X23 a_381_47# SCE a_453_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 a_1572_329# a_193_47# a_1714_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X25 a_1714_47# a_193_47# a_1823_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X26 VGND a_1107_21# a_1619_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X27 VPWR a_1888_21# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X28 a_1401_21# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 a_1714_47# a_27_47# a_1800_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X30 a_764_47# D a_453_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 a_423_315# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X32 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X33 Q_N a_1888_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X34 a_1619_47# a_27_47# a_1714_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X35 a_27_47# CLK_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X36 a_1107_21# a_1401_21# a_1251_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X37 a_1401_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X38 a_27_47# CLK_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X39 a_752_413# D a_453_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X40 a_453_47# a_193_47# a_931_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X41 Q_N a_1888_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X42 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X43 a_453_47# a_27_47# a_931_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X44 VGND SCD a_381_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X45 a_931_47# a_27_47# a_1041_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X46 a_1823_47# a_1888_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X47 Q a_2696_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X48 VPWR SCE a_752_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X49 VPWR SET_B a_1888_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X50 VGND SET_B a_2004_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X51 a_1041_47# a_1107_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__sdfbbp_1 CLK D RESET_B SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
X0 VGND a_423_315# a_764_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VPWR SET_B a_1107_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_423_315# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_1800_413# a_1887_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 VGND SET_B a_1251_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_1107_21# a_1400_21# a_1251_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X6 a_2596_47# a_1887_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 a_1351_329# a_1400_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X8 a_1887_21# a_1714_47# a_2122_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X9 a_2122_329# a_1400_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X10 VGND a_1887_21# Q_N VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_1822_47# a_1887_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_931_47# a_27_47# a_1017_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X13 a_1017_413# a_1107_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X14 a_1107_21# a_931_47# a_1351_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X15 VPWR a_1107_21# a_1572_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X16 VPWR SCD a_381_363# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X17 a_381_363# a_423_315# a_453_363# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 a_1251_47# a_931_47# a_1107_21# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X19 a_1887_21# a_1400_21# a_2026_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X20 a_1572_329# a_27_47# a_1714_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X21 VPWR a_1887_21# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 a_2596_47# a_1887_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_2026_47# a_1714_47# a_1887_21# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X24 a_1400_21# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 a_1714_47# a_193_47# a_1800_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X26 VGND a_2596_47# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 a_764_47# D a_453_363# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 a_1400_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X29 a_423_315# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X30 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 a_381_47# SCE a_453_363# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X32 a_1618_47# a_193_47# a_1714_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X33 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X35 a_752_413# D a_453_363# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X36 a_1714_47# a_27_47# a_1822_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X37 VPWR a_2596_47# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X38 a_453_363# a_27_47# a_931_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X39 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X40 a_453_363# a_193_47# a_931_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X41 VGND SCD a_381_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X42 VGND a_1107_21# a_1618_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X43 a_931_47# a_193_47# a_1041_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X44 VPWR SCE a_752_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X45 VPWR SET_B a_1887_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X46 VGND SET_B a_2026_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X47 a_1041_47# a_1107_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__sdfrbp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q Q_N
X0 a_1245_303# a_193_47# a_1592_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X1 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_1079_413# a_193_47# a_1187_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X3 VGND a_299_66# a_569_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_538_389# D a_620_389# VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=150000u
X5 a_2324_47# a_1767_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
X6 a_620_389# a_193_47# a_1079_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_1592_47# a_193_47# a_1758_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_1245_303# a_27_47# a_1592_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 a_1758_413# a_1767_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_1946_47# a_1592_47# a_1767_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_620_389# a_27_47# a_1079_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X12 a_1293_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 VGND a_1767_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_1191_413# a_1245_303# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 VGND RESET_B a_1946_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_780_389# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=150000u
X17 a_569_119# D a_620_389# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_620_389# a_299_66# a_780_389# VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=150000u
X19 a_620_389# SCE a_817_66# VNB sky130_fd_pr__nfet_01v8 w=420000u l=500000u
X20 VPWR a_2324_47# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
X21 a_2324_47# a_1767_21# VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X22 VPWR a_1079_413# a_1245_303# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X23 VPWR SCE a_538_389# VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=150000u
X24 a_1079_413# a_27_47# a_1191_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X25 VPWR RESET_B a_1191_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X26 a_299_66# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=150000u
X27 a_1187_47# a_1245_303# a_1293_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 VPWR RESET_B a_1767_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X31 a_1767_21# a_1592_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X32 VPWR a_1767_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X33 a_1592_47# a_27_47# a_1701_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X34 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X35 a_299_66# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X36 a_817_66# SCD VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=180000u
X37 VGND a_1079_413# a_1245_303# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X38 a_1701_47# a_1767_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X39 VGND a_2324_47# Q_N VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__sdfrbp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q Q_N
X0 a_1245_303# a_193_47# a_1592_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X1 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_1079_413# a_193_47# a_1187_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X3 a_2135_47# a_1767_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X4 VGND a_299_66# a_569_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_538_389# D a_620_389# VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=150000u
X6 a_620_389# a_193_47# a_1079_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_1592_47# a_193_47# a_1758_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_1245_303# a_27_47# a_1592_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 a_1758_413# a_1767_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_1946_47# a_1592_47# a_1767_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 Q a_1767_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_620_389# a_27_47# a_1079_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X13 a_1293_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_1191_413# a_1245_303# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 VGND RESET_B a_1946_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_780_389# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=150000u
X17 a_569_119# D a_620_389# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_620_389# a_299_66# a_780_389# VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=150000u
X19 a_620_389# SCE a_817_66# VNB sky130_fd_pr__nfet_01v8 w=420000u l=500000u
X20 VPWR a_1079_413# a_1245_303# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X21 VGND a_1767_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 Q_N a_2135_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 VPWR SCE a_538_389# VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=150000u
X24 a_1079_413# a_27_47# a_1191_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X25 VPWR RESET_B a_1191_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X26 Q_N a_2135_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 a_2135_47# a_1767_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 VGND a_2135_47# Q_N VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 a_299_66# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=150000u
X30 a_1187_47# a_1245_303# a_1293_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X32 VPWR a_1767_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X33 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X34 VPWR RESET_B a_1767_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X35 a_1767_21# a_1592_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X36 VPWR a_2135_47# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X37 a_1592_47# a_27_47# a_1701_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X38 Q a_1767_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X39 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X40 a_299_66# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X41 a_817_66# SCD VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=180000u
X42 VGND a_1079_413# a_1245_303# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X43 a_1701_47# a_1767_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__sdfrtn_1 CLK_N D RESET_B SCD SCE VGND VNB VPB VPWR Q
X0 a_1245_303# a_27_47# a_1592_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X1 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_1079_413# a_27_47# a_1187_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X3 VGND a_299_66# a_569_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_538_389# D a_620_389# VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=150000u
X5 a_620_389# a_27_47# a_1079_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_1592_47# a_27_47# a_1758_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_1245_303# a_193_47# a_1592_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_1758_413# a_1767_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 a_1946_47# a_1592_47# a_1767_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_620_389# a_193_47# a_1079_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X11 a_1293_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VGND a_1767_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_1191_413# a_1245_303# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X14 VGND RESET_B a_1946_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_780_389# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=150000u
X16 a_569_119# D a_620_389# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_620_389# a_299_66# a_780_389# VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=150000u
X18 a_620_389# SCE a_817_66# VNB sky130_fd_pr__nfet_01v8 w=420000u l=500000u
X19 VPWR a_1079_413# a_1245_303# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X20 VPWR SCE a_538_389# VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=150000u
X21 a_1079_413# a_193_47# a_1191_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X22 VPWR RESET_B a_1191_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X23 a_299_66# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=150000u
X24 a_1187_47# a_1245_303# a_1293_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 a_27_47# CLK_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 VPWR RESET_B a_1767_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X28 a_1767_21# a_1592_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X29 VPWR a_1767_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X30 a_1592_47# a_193_47# a_1701_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X31 a_27_47# CLK_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X32 a_299_66# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X33 a_817_66# SCD VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=180000u
X34 VGND a_1079_413# a_1245_303# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X35 a_1701_47# a_1767_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__sdfrtp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
X0 a_1245_303# a_193_47# a_1592_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X1 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_1079_413# a_193_47# a_1187_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X3 VGND a_299_66# a_569_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_538_389# D a_620_389# VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=150000u
X5 a_620_389# a_193_47# a_1079_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_1592_47# a_193_47# a_1758_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_1245_303# a_27_47# a_1592_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_1758_413# a_1767_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 a_1946_47# a_1592_47# a_1767_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_620_389# a_27_47# a_1079_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X11 a_1293_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VGND a_1767_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_1191_413# a_1245_303# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X14 VGND RESET_B a_1946_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_780_389# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=150000u
X16 a_569_119# D a_620_389# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_620_389# a_299_66# a_780_389# VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=150000u
X18 a_620_389# SCE a_817_66# VNB sky130_fd_pr__nfet_01v8 w=420000u l=500000u
X19 VPWR a_1079_413# a_1245_303# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X20 VPWR SCE a_538_389# VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=150000u
X21 a_1079_413# a_27_47# a_1191_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X22 VPWR RESET_B a_1191_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X23 a_299_66# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=150000u
X24 a_1187_47# a_1245_303# a_1293_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 VPWR RESET_B a_1767_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X28 a_1767_21# a_1592_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X29 VPWR a_1767_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X30 a_1592_47# a_27_47# a_1701_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X31 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X32 a_299_66# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X33 a_817_66# SCD VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=180000u
X34 VGND a_1079_413# a_1245_303# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X35 a_1701_47# a_1767_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__sdfrtp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
X0 a_1245_303# a_193_47# a_1592_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X1 Q a_1767_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_1079_413# a_193_47# a_1187_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X4 VGND a_299_66# a_569_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_538_389# D a_620_389# VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=150000u
X6 a_620_389# a_193_47# a_1079_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_1592_47# a_193_47# a_1758_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_1245_303# a_27_47# a_1592_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 a_1758_413# a_1767_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_1946_47# a_1592_47# a_1767_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_620_389# a_27_47# a_1079_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X12 a_1293_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 VGND a_1767_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_1191_413# a_1245_303# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 VGND RESET_B a_1946_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_780_389# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=150000u
X17 a_569_119# D a_620_389# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_620_389# a_299_66# a_780_389# VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=150000u
X19 a_620_389# SCE a_817_66# VNB sky130_fd_pr__nfet_01v8 w=420000u l=500000u
X20 VPWR a_1079_413# a_1245_303# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X21 VPWR SCE a_538_389# VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=150000u
X22 a_1079_413# a_27_47# a_1191_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X23 VPWR RESET_B a_1191_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X24 a_299_66# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=150000u
X25 a_1187_47# a_1245_303# a_1293_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 VPWR RESET_B a_1767_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X29 a_1767_21# a_1592_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X30 VPWR a_1767_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X31 a_1592_47# a_27_47# a_1701_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X32 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X33 a_299_66# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 a_817_66# SCD VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=180000u
X35 VGND a_1079_413# a_1245_303# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X36 a_1701_47# a_1767_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X37 Q a_1767_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__sdfrtp_4 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
X0 a_1245_303# a_193_47# a_1592_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X1 Q a_1767_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_1079_413# a_193_47# a_1187_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X4 Q a_1767_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VGND a_299_66# a_569_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_538_389# D a_620_389# VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=150000u
X7 a_620_389# a_193_47# a_1079_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_1592_47# a_193_47# a_1758_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 a_1245_303# a_27_47# a_1592_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_1758_413# a_1767_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 a_1946_47# a_1592_47# a_1767_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VGND a_1767_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_620_389# a_27_47# a_1079_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X14 a_1293_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 VGND a_1767_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_1191_413# a_1245_303# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X17 VGND RESET_B a_1946_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_780_389# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=150000u
X19 a_569_119# D a_620_389# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_620_389# a_299_66# a_780_389# VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=150000u
X21 a_620_389# SCE a_817_66# VNB sky130_fd_pr__nfet_01v8 w=420000u l=500000u
X22 VPWR a_1079_413# a_1245_303# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X23 VPWR SCE a_538_389# VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=150000u
X24 a_1079_413# a_27_47# a_1191_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X25 VPWR RESET_B a_1191_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X26 a_299_66# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=540000u l=150000u
X27 a_1187_47# a_1245_303# a_1293_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 VPWR RESET_B a_1767_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X31 a_1767_21# a_1592_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X32 VPWR a_1767_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X33 a_1592_47# a_27_47# a_1701_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X34 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X35 a_299_66# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X36 a_817_66# SCD VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=180000u
X37 VGND a_1079_413# a_1245_303# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X38 VPWR a_1767_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X39 a_1701_47# a_1767_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X40 Q a_1767_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X41 Q a_1767_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__sdfsbp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
X0 a_1087_47# a_1129_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_1879_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VPWR a_1587_329# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VPWR a_643_369# a_809_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X4 a_1129_21# a_997_413# a_1347_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_319_21# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X6 a_265_47# a_319_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_1347_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_643_369# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 VPWR a_997_413# a_1514_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X10 VPWR a_1587_329# a_1770_295# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 a_1587_329# a_809_369# a_1712_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X12 a_1514_329# a_643_369# a_1587_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X13 a_1807_47# a_1770_295# a_1879_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_1129_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 a_181_47# D a_265_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_319_21# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_997_413# a_809_369# a_1087_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 VGND a_997_413# a_1514_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X19 VGND a_2412_47# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 VPWR a_2412_47# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 a_109_47# SCE a_181_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_643_369# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_997_413# a_643_369# a_1081_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X24 VPWR a_997_413# a_1129_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X25 a_1514_47# a_809_369# a_1587_329# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X26 a_181_47# a_319_21# a_27_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X27 a_2412_47# a_1587_329# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X28 a_1712_413# a_1770_295# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X29 a_27_369# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X30 VPWR SCE a_193_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X31 a_181_47# a_809_369# a_997_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X32 a_1587_329# a_643_369# a_1807_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X33 VGND a_1587_329# a_1770_295# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 a_193_369# D a_181_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X35 VGND SCD a_109_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X36 VGND a_643_369# a_809_369# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X37 VGND a_1587_329# Q_N VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X38 VPWR SET_B a_1587_329# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X39 a_1081_413# a_1129_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X40 a_181_47# a_643_369# a_997_413# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X41 a_2412_47# a_1587_329# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__sdfsbp_2 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
X0 a_1132_21# a_1006_47# a_1350_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_1885_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_181_47# a_652_47# a_1006_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VGND a_1597_329# a_1781_295# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VPWR a_1006_47# a_1525_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X5 Q_N a_1597_329# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_1525_329# a_652_47# a_1597_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X7 a_1597_329# a_818_47# a_1723_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_1350_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_2501_47# a_1597_329# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 Q a_2501_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_1006_47# a_652_47# a_1102_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X12 a_1132_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X13 a_1006_47# a_818_47# a_1090_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 VPWR a_1006_47# a_1132_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 a_1813_47# a_1781_295# a_1885_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_181_47# D a_265_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_265_47# a_328_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_1517_47# a_818_47# a_1597_329# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X19 VGND a_1597_329# Q_N VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_181_47# a_818_47# a_1006_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X21 VPWR a_1597_329# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 a_1723_413# a_1781_295# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X23 a_109_47# SCE a_181_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 a_328_21# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 VGND a_1006_47# a_1517_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X26 VPWR SET_B a_1597_329# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X27 VGND a_2501_47# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 a_652_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X29 a_652_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X30 a_1102_413# a_1132_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X31 Q_N a_1597_329# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X32 a_27_369# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X33 VPWR SCE a_193_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X34 a_1597_329# a_652_47# a_1813_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 a_193_369# D a_181_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X36 a_181_47# a_328_21# a_27_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X37 VGND SCD a_109_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X38 VPWR a_2501_47# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X39 a_2501_47# a_1597_329# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X40 a_1090_47# a_1132_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X41 VPWR a_652_47# a_818_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X42 VPWR a_1597_329# a_1781_295# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X43 VGND a_652_47# a_818_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X44 a_328_21# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X45 Q a_2501_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__sdfstp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
X0 a_1087_47# a_1129_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VPWR a_997_413# a_1525_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X2 a_1525_329# a_643_369# a_1597_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X3 a_1597_329# a_809_369# a_1723_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_1597_329# a_643_369# a_1815_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VPWR a_643_369# a_809_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X6 a_1129_21# a_997_413# a_1347_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_319_21# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X8 a_1129_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 a_265_47# a_319_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_1347_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_643_369# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X12 VPWR a_2227_47# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VPWR a_997_413# a_1129_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X14 a_181_47# D a_265_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_319_21# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_997_413# a_809_369# a_1087_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 VGND a_997_413# a_1514_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X18 a_1514_47# a_809_369# a_1597_329# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X19 VGND a_1597_329# a_1781_295# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_1723_413# a_1781_295# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X21 a_109_47# SCE a_181_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_643_369# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_997_413# a_643_369# a_1081_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X24 a_181_47# a_319_21# a_27_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X25 a_1887_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 a_27_369# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X27 VPWR SCE a_193_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X28 a_181_47# a_809_369# a_997_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X29 a_193_369# D a_181_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X30 a_1815_47# a_1781_295# a_1887_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 VPWR a_1597_329# a_1781_295# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X32 VGND SCD a_109_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X33 a_2227_47# a_1597_329# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X34 VGND a_643_369# a_809_369# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 VGND a_2227_47# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X36 VPWR SET_B a_1597_329# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X37 a_1081_413# a_1129_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X38 a_181_47# a_643_369# a_997_413# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X39 a_2227_47# a_1597_329# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__sdfstp_2 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
X0 a_1087_47# a_1129_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VPWR a_997_413# a_1525_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X2 Q a_2227_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_1525_329# a_643_369# a_1597_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X4 a_1597_329# a_809_369# a_1723_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_1597_329# a_643_369# a_1815_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VGND a_2227_47# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VPWR a_643_369# a_809_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X8 a_1129_21# a_997_413# a_1347_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_319_21# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X10 a_1129_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 a_265_47# a_319_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_1347_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_643_369# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X14 VPWR a_2227_47# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 VPWR a_997_413# a_1129_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X16 a_181_47# D a_265_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_319_21# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_997_413# a_809_369# a_1087_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 VGND a_997_413# a_1514_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X20 a_1514_47# a_809_369# a_1597_329# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X21 VGND a_1597_329# a_1781_295# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_1723_413# a_1781_295# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X23 a_109_47# SCE a_181_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 a_643_369# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 a_997_413# a_643_369# a_1081_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X26 a_181_47# a_319_21# a_27_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X27 a_1887_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 a_27_369# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X29 VPWR SCE a_193_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X30 a_181_47# a_809_369# a_997_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X31 a_193_369# D a_181_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X32 a_1815_47# a_1781_295# a_1887_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X33 VPWR a_1597_329# a_1781_295# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X34 VGND SCD a_109_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 a_2227_47# a_1597_329# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X36 VGND a_643_369# a_809_369# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X37 VPWR SET_B a_1597_329# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X38 Q a_2227_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X39 a_1081_413# a_1129_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X40 a_181_47# a_643_369# a_997_413# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X41 a_2227_47# a_1597_329# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__sdfstp_4 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
X0 a_1087_47# a_1129_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VPWR a_997_413# a_1525_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X2 VPWR a_2227_47# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_1525_329# a_643_369# a_1597_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X4 a_1597_329# a_809_369# a_1723_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_1597_329# a_643_369# a_1815_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VGND a_2227_47# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VPWR a_643_369# a_809_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X8 a_1129_21# a_997_413# a_1347_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 Q a_2227_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_319_21# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X11 a_1129_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X12 a_265_47# a_319_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_1347_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_643_369# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X15 a_2227_47# a_1597_329# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 VPWR a_2227_47# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 Q a_2227_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 VPWR a_997_413# a_1129_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X19 a_181_47# D a_265_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_319_21# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 a_997_413# a_809_369# a_1087_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 VGND a_997_413# a_1514_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X23 a_1514_47# a_809_369# a_1597_329# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X24 VGND a_1597_329# a_1781_295# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 VGND a_2227_47# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 a_1723_413# a_1781_295# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X27 a_109_47# SCE a_181_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 a_643_369# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 a_997_413# a_643_369# a_1081_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X30 a_181_47# a_319_21# a_27_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X31 a_1887_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X32 a_27_369# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X33 VPWR SCE a_193_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X34 a_181_47# a_809_369# a_997_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X35 a_193_369# D a_181_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X36 a_1815_47# a_1781_295# a_1887_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X37 VPWR a_1597_329# a_1781_295# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X38 VGND SCD a_109_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X39 VGND a_643_369# a_809_369# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X40 VPWR SET_B a_1597_329# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X41 a_1081_413# a_1129_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X42 a_181_47# a_643_369# a_997_413# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X43 Q a_2227_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X44 a_2227_47# a_1597_329# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X45 Q a_2227_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__sdfxbp_1 CLK D SCD SCE VGND VNB VPB VPWR Q Q_N
X0 a_1089_183# a_193_47# a_1346_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X1 VPWR SCE a_465_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 a_1027_47# a_1089_183# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_1023_413# a_1089_183# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 VPWR a_1948_47# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_299_47# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X6 a_1517_315# a_1346_413# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_930_413# a_193_47# a_1027_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X8 a_1089_183# a_27_47# a_1346_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 a_1517_315# a_1346_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_640_369# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X11 VPWR a_1517_315# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_483_47# D a_556_369# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_1346_413# a_193_47# a_1430_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X14 a_1948_47# a_1517_315# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_465_369# D a_556_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X16 a_556_369# SCE a_657_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 VGND a_930_413# a_1089_183# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X18 a_556_369# a_193_47# a_930_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X19 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 VPWR a_930_413# a_1089_183# VPB sky130_fd_pr__pfet_01v8_hvt w=750000u l=150000u
X22 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X23 a_1948_47# a_1517_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X24 a_930_413# a_27_47# a_1023_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X25 a_556_369# a_27_47# a_930_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X26 a_1346_413# a_27_47# a_1475_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X27 VGND a_1948_47# Q_N VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X29 a_556_369# a_299_47# a_640_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X30 a_299_47# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 a_657_47# SCD VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X32 a_1430_413# a_1517_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X33 VGND a_299_47# a_483_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 a_1475_47# a_1517_315# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 VGND a_1517_315# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__sdfxbp_2 CLK D SCD SCE VGND VNB VPB VPWR Q Q_N
X0 a_560_369# a_299_47# a_644_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X1 a_1097_183# a_27_47# a_1354_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_2049_47# a_1525_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X3 a_560_369# a_193_47# a_938_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 VPWR a_938_413# a_1097_183# VPB sky130_fd_pr__pfet_01v8_hvt w=750000u l=150000u
X6 a_1035_47# a_1097_183# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_466_369# D a_560_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X8 a_1525_315# a_1354_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VGND a_2049_47# Q_N VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VPWR SCE a_466_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X11 a_560_369# SCE a_661_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_1354_413# a_27_47# a_1483_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X13 VGND a_938_413# a_1097_183# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X14 VGND a_1525_315# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_299_47# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X16 a_487_47# D a_560_369# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_560_369# a_27_47# a_938_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X18 a_1097_183# a_193_47# a_1354_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X19 VPWR a_2049_47# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 a_1438_413# a_1525_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X21 VPWR a_1525_315# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 a_1483_47# a_1525_315# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_644_369# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X24 a_299_47# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 a_938_413# a_27_47# a_1031_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X26 a_661_47# SCD VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 Q_N a_2049_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X28 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 VGND a_299_47# a_487_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X30 Q a_1525_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X31 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X32 Q_N a_2049_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X33 a_1525_315# a_1354_413# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X34 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X35 a_938_413# a_193_47# a_1035_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X36 a_1031_413# a_1097_183# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X37 a_1354_413# a_193_47# a_1438_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X38 Q a_1525_315# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X39 a_2049_47# a_1525_315# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__sdfxtp_1 CLK D SCD SCE VGND VNB VPB VPWR Q
X0 a_1478_47# a_1520_315# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 a_1092_183# a_193_47# a_1349_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X3 a_1520_315# a_1349_413# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VPWR SCE a_467_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 a_1433_413# a_1520_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_1030_47# a_1092_183# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VPWR a_1520_315# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_299_47# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 a_933_413# a_193_47# a_1030_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X10 a_640_369# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X11 a_1092_183# a_27_47# a_1349_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X12 a_483_47# D a_556_369# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_467_369# D a_556_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X14 a_299_47# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_556_369# SCE a_657_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_1026_413# a_1092_183# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X17 a_1349_413# a_193_47# a_1433_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X18 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 VGND a_933_413# a_1092_183# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X21 VGND a_1520_315# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 a_1520_315# a_1349_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X23 a_556_369# a_299_47# a_640_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X24 a_556_369# a_193_47# a_933_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X25 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X26 a_657_47# SCD VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 VGND a_299_47# a_483_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 VPWR a_933_413# a_1092_183# VPB sky130_fd_pr__pfet_01v8_hvt w=750000u l=150000u
X29 a_933_413# a_27_47# a_1026_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X30 a_556_369# a_27_47# a_933_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X31 a_1349_413# a_27_47# a_1478_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__sdfxtp_2 CLK D SCD SCE VGND VNB VPB VPWR Q
X0 a_660_47# SCD VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_1355_413# a_193_47# a_1439_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 VGND a_1526_315# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VGND a_299_47# a_486_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_1526_315# a_1355_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X6 a_1098_183# a_27_47# a_1355_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_1098_183# a_193_47# a_1355_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X8 a_559_369# a_193_47# a_939_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 VPWR SCE a_467_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X10 a_1484_47# a_1526_315# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_299_47# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X12 a_1526_315# a_1355_413# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VPWR a_939_413# a_1098_183# VPB sky130_fd_pr__pfet_01v8_hvt w=750000u l=150000u
X14 a_559_369# SCE a_660_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_643_369# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X16 a_939_413# a_193_47# a_1036_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X17 VPWR a_1526_315# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 a_1439_413# a_1526_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X19 Q a_1526_315# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_299_47# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 a_486_47# D a_559_369# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_939_413# a_27_47# a_1032_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X24 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 VGND a_939_413# a_1098_183# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X26 Q a_1526_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 a_467_369# D a_559_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X28 a_1036_47# a_1098_183# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X30 a_559_369# a_27_47# a_939_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X31 a_1355_413# a_27_47# a_1484_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X32 a_559_369# a_299_47# a_643_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X33 a_1032_413# a_1098_183# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__sdfxtp_4 CLK D SCD SCE VGND VNB VPB VPWR Q
X0 Q a_1527_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 Q a_1527_315# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_560_369# a_299_47# a_644_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X3 a_1033_413# a_1099_183# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 VPWR a_1527_315# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X6 VPWR a_1527_315# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_1527_315# a_1356_413# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_466_369# D a_560_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 a_1099_183# a_27_47# a_1356_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_1527_315# a_1356_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 Q a_1527_315# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VPWR SCE a_466_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X13 a_560_369# SCE a_661_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_940_413# a_193_47# a_1037_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X15 VGND a_1527_315# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_1356_413# a_193_47# a_1440_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X17 a_299_47# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 a_487_47# D a_560_369# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_560_369# a_193_47# a_940_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X20 VGND a_940_413# a_1099_183# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X21 Q a_1527_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 VPWR a_940_413# a_1099_183# VPB sky130_fd_pr__pfet_01v8_hvt w=750000u l=150000u
X23 a_1037_47# a_1099_183# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 a_644_369# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X25 a_560_369# a_27_47# a_940_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X26 a_1356_413# a_27_47# a_1485_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X27 a_299_47# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 a_1440_413# a_1527_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X29 a_661_47# SCD VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X30 VGND a_1527_315# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X32 VGND a_299_47# a_487_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X33 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 a_940_413# a_27_47# a_1033_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X35 a_1485_47# a_1527_315# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X36 a_1099_183# a_193_47# a_1356_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X37 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__sdlclkp_1 CLK GATE SCE VGND VNB VPB VPWR GCLK
X0 a_1012_47# a_464_315# a_1094_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VGND a_1012_47# GCLK VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_27_47# a_256_243# a_286_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_286_413# a_256_147# a_382_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 VGND CLK a_256_147# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_256_243# a_256_147# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X6 a_394_47# a_464_315# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_256_243# a_256_147# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VPWR a_286_413# a_464_315# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_1012_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X10 VPWR SCE a_109_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X11 VGND GATE a_27_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VPWR a_464_315# a_1012_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X13 a_27_47# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_286_413# a_256_243# a_394_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X15 VPWR a_1012_47# GCLK VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 a_27_47# a_256_147# a_286_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X17 a_109_369# GATE a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 VGND a_286_413# a_464_315# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 VPWR CLK a_256_147# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X20 a_1094_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 a_382_413# a_464_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__sdlclkp_2 CLK GATE SCE VGND VNB VPB VPWR GCLK
X0 a_383_413# a_465_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 VGND a_287_413# a_465_315# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_1102_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_395_47# a_465_315# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VPWR a_1020_47# GCLK VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_27_47# a_257_147# a_287_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X6 a_1020_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 a_27_47# a_257_243# a_287_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 GCLK a_1020_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_287_413# a_257_147# a_383_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 GCLK a_1020_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_1020_47# a_465_315# a_1102_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_287_413# a_257_243# a_395_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X13 VGND CLK a_257_147# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 VPWR a_287_413# a_465_315# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_257_243# a_257_147# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 VPWR SCE a_109_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X17 a_257_243# a_257_147# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 VPWR CLK a_257_147# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X19 VGND GATE a_27_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 VGND a_1020_47# GCLK VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 a_27_47# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_109_369# GATE a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X23 VPWR a_465_315# a_1020_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__sdlclkp_4 CLK GATE SCE VGND VNB VPB VPWR GCLK
X0 VPWR a_1045_47# GCLK VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_383_413# a_465_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 VPWR a_1045_47# GCLK VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 VGND a_287_413# a_465_315# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VPWR CLK a_257_147# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 VGND a_1045_47# GCLK VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR a_465_315# a_1045_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 GCLK a_1045_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_395_47# a_465_315# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_27_47# a_257_147# a_287_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X10 a_1127_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 GCLK a_1045_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_27_47# a_257_243# a_287_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X13 a_1045_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_287_413# a_257_147# a_383_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 a_287_413# a_257_243# a_395_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X16 VGND CLK a_257_147# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_257_243# a_257_147# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 VPWR a_287_413# a_465_315# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_257_243# a_257_147# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_1045_47# a_465_315# a_1127_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 VGND a_1045_47# GCLK VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 VPWR SCE a_109_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X23 VGND GATE a_27_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 a_27_47# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 a_109_369# GATE a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X26 GCLK a_1045_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 GCLK a_1045_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__sedfxbp_1 CLK D DE SCD SCE VGND VNB VPB VPWR Q Q_N
X0 VPWR a_1610_159# a_1960_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_1446_413# a_27_47# a_1537_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_729_47# a_791_264# a_299_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VPWR a_2051_413# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VPWR SCD a_1231_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 a_791_264# a_2051_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X6 a_2051_413# a_193_47# a_2135_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_299_47# D a_381_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X8 a_381_369# a_423_343# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 a_1226_119# SCE a_915_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_1960_413# a_27_47# a_2051_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 VGND a_1446_413# a_1610_159# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X12 VGND a_791_264# Q_N VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_1231_369# a_885_21# a_915_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X14 a_2135_413# a_791_264# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 a_915_47# a_27_47# a_1446_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X16 a_2051_413# a_27_47# a_2177_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X17 VPWR DE a_729_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 a_299_47# a_885_21# a_915_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_381_47# DE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 VPWR a_1446_413# a_1610_159# VPB sky130_fd_pr__pfet_01v8_hvt w=750000u l=150000u
X21 VGND a_1610_159# a_1974_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_1974_47# a_193_47# a_2051_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X23 VGND SCD a_1226_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 a_729_369# a_791_264# a_299_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X25 a_2177_47# a_791_264# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 a_299_47# SCE a_915_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X27 a_423_343# DE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 a_915_47# a_193_47# a_1446_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X29 VGND a_2051_413# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 VPWR a_791_264# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X31 a_885_21# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X32 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X33 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 VGND a_423_343# a_729_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 a_1561_47# a_1610_159# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X36 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X37 a_1537_413# a_1610_159# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X38 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X39 a_299_47# D a_381_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X40 a_1446_413# a_193_47# a_1561_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X41 a_791_264# a_2051_413# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X42 a_423_343# DE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X43 a_885_21# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__sedfxbp_2 CLK D DE SCD SCE VGND VNB VPB VPWR Q Q_N
X0 VPWR a_1610_159# a_1960_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 Q_N a_791_264# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_791_264# a_2051_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X3 a_1446_413# a_27_47# a_1537_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_729_47# a_791_264# a_299_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 Q a_2051_413# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR SCD a_1231_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 Q a_2051_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_2051_413# a_193_47# a_2135_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 VGND a_2051_413# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_299_47# D a_381_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X11 a_381_369# a_423_343# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X12 VPWR a_2051_413# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_1226_119# SCE a_915_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_1960_413# a_27_47# a_2051_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 VGND a_1446_413# a_1610_159# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X16 VGND a_791_264# Q_N VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 a_1231_369# a_885_21# a_915_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 a_2135_413# a_791_264# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X19 a_915_47# a_27_47# a_1446_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X20 a_2051_413# a_27_47# a_2177_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X21 VPWR DE a_729_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X22 a_299_47# a_885_21# a_915_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_381_47# DE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 VPWR a_1446_413# a_1610_159# VPB sky130_fd_pr__pfet_01v8_hvt w=750000u l=150000u
X25 VGND a_1610_159# a_1974_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 a_1974_47# a_193_47# a_2051_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X27 VGND SCD a_1226_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 a_729_369# a_791_264# a_299_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X29 a_2177_47# a_791_264# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X30 a_299_47# SCE a_915_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X31 a_423_343# DE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X32 a_915_47# a_193_47# a_1446_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X33 VPWR a_791_264# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X34 a_791_264# a_2051_413# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 a_885_21# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X36 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X37 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X38 VGND a_423_343# a_729_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X39 a_1561_47# a_1610_159# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X40 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X41 a_1537_413# a_1610_159# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X42 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X43 a_299_47# D a_381_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X44 a_1446_413# a_193_47# a_1561_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X45 a_423_343# DE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X46 a_885_21# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X47 Q_N a_791_264# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__sedfxtp_1 CLK D DE SCD SCE VGND VNB VPB VPWR Q
X0 VPWR a_1610_159# a_1960_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_791_264# a_2051_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 a_1446_413# a_27_47# a_1537_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_729_47# a_791_264# a_299_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VPWR SCD a_1231_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 a_2051_413# a_193_47# a_2135_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_299_47# D a_381_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 a_381_369# a_423_343# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X8 a_1226_119# SCE a_915_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_1960_413# a_27_47# a_2051_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 VGND a_1446_413# a_1610_159# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X11 a_1231_369# a_885_21# a_915_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X12 a_2135_413# a_791_264# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X13 a_915_47# a_27_47# a_1446_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X14 a_2051_413# a_27_47# a_2177_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X15 VPWR DE a_729_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X16 a_299_47# a_885_21# a_915_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_381_47# DE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 VPWR a_1446_413# a_1610_159# VPB sky130_fd_pr__pfet_01v8_hvt w=750000u l=150000u
X19 VGND a_1610_159# a_1974_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_1974_47# a_193_47# a_2051_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X21 VGND a_2051_413# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 VGND SCD a_1226_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_729_369# a_791_264# a_299_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X24 a_2177_47# a_791_264# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 a_299_47# SCE a_915_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X26 a_423_343# DE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 a_915_47# a_193_47# a_1446_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X28 a_791_264# a_2051_413# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 a_885_21# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X30 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X32 VGND a_423_343# a_729_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X33 a_1561_47# a_1610_159# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X35 a_1537_413# a_1610_159# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X36 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X37 a_299_47# D a_381_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X38 a_1446_413# a_193_47# a_1561_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X39 a_423_343# DE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X40 a_885_21# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X41 VPWR a_2051_413# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__sedfxtp_2 CLK D DE SCD SCE VGND VNB VPB VPWR Q
X0 VPWR a_1610_159# a_1960_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_791_264# a_2051_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 a_1446_413# a_27_47# a_1537_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_729_47# a_791_264# a_299_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 Q a_2051_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 Q a_2051_413# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR SCD a_1231_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 a_2051_413# a_193_47# a_2135_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_299_47# D a_381_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 a_381_369# a_423_343# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X10 a_1226_119# SCE a_915_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_1960_413# a_27_47# a_2051_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X12 VGND a_1446_413# a_1610_159# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X13 a_1231_369# a_885_21# a_915_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X14 a_2135_413# a_791_264# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 a_915_47# a_27_47# a_1446_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X16 a_2051_413# a_27_47# a_2177_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X17 VPWR DE a_729_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 a_299_47# a_885_21# a_915_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_381_47# DE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 VPWR a_1446_413# a_1610_159# VPB sky130_fd_pr__pfet_01v8_hvt w=750000u l=150000u
X21 VGND a_1610_159# a_1974_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_1974_47# a_193_47# a_2051_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X23 VGND a_2051_413# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 VGND SCD a_1226_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 a_729_369# a_791_264# a_299_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X26 a_2177_47# a_791_264# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 a_299_47# SCE a_915_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X28 a_423_343# DE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 a_915_47# a_193_47# a_1446_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X30 a_791_264# a_2051_413# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 a_885_21# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X32 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X33 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 VGND a_423_343# a_729_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 a_1561_47# a_1610_159# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X36 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X37 a_1537_413# a_1610_159# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X38 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X39 a_299_47# D a_381_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X40 a_1446_413# a_193_47# a_1561_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X41 a_423_343# DE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X42 a_885_21# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X43 VPWR a_2051_413# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__sedfxtp_4 CLK D DE SCD SCE VGND VNB VPB VPWR Q
X0 VPWR a_1610_159# a_1960_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_791_264# a_2051_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 a_1446_413# a_27_47# a_1537_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_729_47# a_791_264# a_299_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 Q a_2051_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 Q a_2051_413# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR SCD a_1231_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 a_2051_413# a_193_47# a_2135_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_299_47# D a_381_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 a_381_369# a_423_343# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X10 Q a_2051_413# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_1226_119# SCE a_915_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_1960_413# a_27_47# a_2051_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X13 VGND a_1446_413# a_1610_159# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X14 Q a_2051_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_1231_369# a_885_21# a_915_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X16 a_2135_413# a_791_264# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X17 a_915_47# a_27_47# a_1446_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X18 a_2051_413# a_27_47# a_2177_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X19 VPWR DE a_729_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X20 a_299_47# a_885_21# a_915_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 VGND a_2051_413# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 a_381_47# DE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 VPWR a_1446_413# a_1610_159# VPB sky130_fd_pr__pfet_01v8_hvt w=750000u l=150000u
X24 VGND a_1610_159# a_1974_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 VPWR a_2051_413# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 a_1974_47# a_193_47# a_2051_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X27 VGND a_2051_413# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 VGND SCD a_1226_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 a_729_369# a_791_264# a_299_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X30 a_2177_47# a_791_264# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 a_299_47# SCE a_915_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X32 a_423_343# DE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X33 a_915_47# a_193_47# a_1446_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X34 a_791_264# a_2051_413# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 a_885_21# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X36 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X37 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X38 VGND a_423_343# a_729_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X39 a_1561_47# a_1610_159# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X40 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X41 a_1537_413# a_1610_159# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X42 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X43 a_299_47# D a_381_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X44 a_1446_413# a_193_47# a_1561_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X45 a_423_343# DE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X46 a_885_21# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X47 VPWR a_2051_413# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__tap_1 VGND VNB VPB VPWR
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__tap_2 VGND VNB VPB VPWR
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__tapvgnd2_1 VGND VPB VPWR
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__tapvgnd_1 VGND VPB VPWR
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
X0 VPWR A a_377_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_377_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 Y a_47_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_129_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VGND B a_285_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_47_47# B a_129_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR B a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_47_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND A a_285_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_285_47# a_47_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
X0 VPWR B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VGND B a_560_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 Y B a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VPWR A a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_27_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_474_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 Y a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_474_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_560_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VPWR a_27_297# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_27_47# B a_27_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_560_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 Y a_27_297# a_560_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 a_27_297# B a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 VGND A a_560_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 a_560_47# a_27_297# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
X0 VGND A a_38_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_38_297# B a_38_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VGND A a_38_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_38_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VPWR A a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 VPWR a_38_297# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_38_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VPWR a_38_297# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_38_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_820_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 Y a_38_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_38_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_820_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 Y a_38_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 Y a_38_297# a_902_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 VGND B a_902_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_38_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X17 Y B a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 a_38_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 VGND B a_902_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_902_47# a_38_297# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 Y B a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 a_902_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 a_902_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 a_902_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 VPWR A a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 a_38_297# B a_38_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 VGND A a_902_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 VGND A a_902_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 a_820_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X30 a_38_47# B a_38_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 Y a_38_297# a_902_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X32 VPWR A a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X33 a_902_47# a_38_297# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X34 a_38_47# B a_38_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X35 VPWR B a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X36 a_902_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X37 VPWR B a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X38 a_820_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X39 VPWR A a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__xnor3_1 A B C VGND VNB VPB VPWR X
X0 a_355_49# C a_78_199# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X1 VGND C a_216_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_841_297# B a_331_325# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X3 a_331_325# a_735_297# a_1106_49# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 X a_78_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_1106_49# B a_331_325# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X6 VGND a_841_297# a_1106_49# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X7 VGND B a_735_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VPWR C a_216_93# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 a_355_49# a_735_297# a_1106_49# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X10 a_1106_49# B a_355_49# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X11 a_841_297# A VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X12 a_331_325# C a_78_199# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X13 VPWR B a_735_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_841_297# B a_355_49# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X15 a_331_325# a_735_297# a_841_297# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X16 X a_78_199# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 VPWR a_841_297# a_1106_49# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 a_78_199# a_216_93# a_355_49# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X19 a_841_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 a_78_199# a_216_93# a_331_325# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X21 a_355_49# a_735_297# a_841_297# VNB sky130_fd_pr__nfet_01v8 w=600000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__xnor3_2 A B C VGND VNB VPB VPWR X
X0 VPWR a_87_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_933_297# B a_423_325# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X2 a_447_49# a_827_297# a_1198_49# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X3 X a_87_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_447_49# C a_87_21# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X5 VPWR C a_308_93# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X6 VGND a_87_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_423_325# C a_87_21# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X8 a_87_21# a_308_93# a_423_325# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X9 a_447_49# a_827_297# a_933_297# VNB sky130_fd_pr__nfet_01v8 w=600000u l=150000u
X10 a_423_325# a_827_297# a_933_297# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X11 a_933_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 a_87_21# a_308_93# a_447_49# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X13 VGND C a_308_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_423_325# a_827_297# a_1198_49# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 VGND a_933_297# a_1198_49# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X16 VGND B a_827_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 VPWR a_933_297# a_1198_49# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 X a_87_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 VPWR B a_827_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X20 a_1198_49# B a_423_325# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X21 a_1198_49# B a_447_49# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X22 a_933_297# A VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X23 a_933_297# B a_447_49# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__xnor3_4 A B C VGND VNB VPB VPWR X
X0 a_1382_49# B a_607_325# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X1 a_631_49# C a_101_21# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X2 VGND a_1117_297# a_1382_49# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X3 VPWR a_101_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VPWR B a_1011_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_1382_49# B a_631_49# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X6 a_1117_297# A VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X7 a_1117_297# B a_631_49# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X8 a_1117_297# B a_607_325# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X9 VGND a_101_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_631_49# a_1011_297# a_1382_49# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X11 X a_101_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VPWR C a_492_93# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X13 a_101_21# a_492_93# a_631_49# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X14 a_101_21# a_492_93# a_607_325# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X15 a_631_49# a_1011_297# a_1117_297# VNB sky130_fd_pr__nfet_01v8 w=600000u l=150000u
X16 a_607_325# C a_101_21# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X17 a_607_325# a_1011_297# a_1117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X18 X a_101_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 VGND B a_1011_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 VPWR a_1117_297# a_1382_49# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 X a_101_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 VGND a_101_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 VGND C a_492_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 a_1117_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 a_607_325# a_1011_297# a_1382_49# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 X a_101_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 VPWR a_101_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
X0 a_35_297# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VGND B a_35_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 X a_35_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_285_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VPWR A a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_35_297# B a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_117_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_285_47# B X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_285_297# a_35_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 VGND A a_285_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_112_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 X a_112_47# a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_27_297# B a_112_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_470_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_112_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VGND A a_470_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 X a_112_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_470_47# B X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VGND B a_112_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_470_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_470_297# a_112_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VPWR A a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_470_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 VGND A a_112_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 X B a_470_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 a_112_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 VPWR B a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 VGND a_112_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
X0 a_806_297# a_112_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 VGND A a_806_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 VGND a_112_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VPWR B a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 VPWR A a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 a_112_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND B a_112_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_806_47# B X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VPWR A a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_806_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VGND B a_112_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_806_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_806_297# a_112_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 a_806_47# B X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 a_806_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_112_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 VGND A a_112_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 a_27_297# B a_112_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 VGND A a_806_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 VGND a_112_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 a_112_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X25 VGND A a_112_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 a_806_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 a_806_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X28 X a_112_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 X B a_806_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 a_112_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 X a_112_47# a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X32 a_112_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X33 a_112_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X34 VPWR B a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X35 X B a_806_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X36 X a_112_47# a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X37 X a_112_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X38 a_27_297# B a_112_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X39 a_806_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__xor3_1 A B C VGND VNB VPB VPWR X
X0 a_112_21# a_266_93# a_404_49# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X1 a_386_325# a_827_297# a_1198_49# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 X a_112_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_386_325# a_827_297# a_931_365# VNB sky130_fd_pr__nfet_01v8 w=600000u l=150000u
X4 a_404_49# a_827_297# a_931_365# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X5 a_931_365# B a_404_49# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X6 a_404_49# C a_112_21# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X7 a_931_365# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 a_404_49# a_827_297# a_1198_49# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_386_325# C a_112_21# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X10 VGND a_931_365# a_1198_49# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X11 VPWR a_931_365# a_1198_49# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 VPWR B a_827_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VGND C a_266_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_112_21# a_266_93# a_386_325# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X15 VGND B a_827_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_931_365# B a_386_325# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X17 a_1198_49# B a_404_49# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 a_1198_49# B a_386_325# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X19 a_931_365# A VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X20 VPWR C a_266_93# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X21 X a_112_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__xor3_2 A B C VGND VNB VPB VPWR X
X0 a_478_325# C a_120_21# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X1 VGND C a_358_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VGND B a_919_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR a_1023_365# a_1290_49# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_1290_49# B a_478_325# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X5 a_1023_365# A VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X6 X a_120_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VPWR B a_919_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X8 VGND a_120_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_1290_49# B a_496_49# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X10 a_496_49# C a_120_21# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X11 a_1023_365# B a_478_325# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X12 VPWR C a_358_93# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X13 a_478_325# a_919_297# a_1023_365# VNB sky130_fd_pr__nfet_01v8 w=600000u l=150000u
X14 a_496_49# a_919_297# a_1290_49# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_120_21# a_358_93# a_496_49# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X16 a_1023_365# B a_496_49# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X17 X a_120_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 a_496_49# a_919_297# a_1023_365# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X19 VGND a_1023_365# a_1290_49# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X20 VPWR a_120_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X21 a_478_325# a_919_297# a_1290_49# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X22 a_120_21# a_358_93# a_478_325# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X23 a_1023_365# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends


******* EOF

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__xor3_4 A B C VGND VNB VPB VPWR X
X0 a_602_325# a_1031_297# a_1402_49# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X1 VGND C a_480_297# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VGND a_1135_365# a_1402_49# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X3 a_602_325# C a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X4 a_602_325# a_1031_297# a_1135_365# VNB sky130_fd_pr__nfet_01v8 w=600000u l=150000u
X5 a_608_49# a_1031_297# a_1135_365# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X6 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_1135_365# B a_608_49# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X8 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_608_49# C a_79_21# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X10 a_1135_365# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X12 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_608_49# a_1031_297# a_1402_49# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 a_1402_49# B a_608_49# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X16 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 VGND B a_1031_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 VPWR C a_480_297# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X19 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 a_79_21# a_480_297# a_602_325# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X22 a_1402_49# B a_602_325# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X23 a_1135_365# A VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X24 a_1135_365# B a_602_325# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X25 VPWR B a_1031_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X26 VPWR a_1135_365# a_1402_49# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X27 a_79_21# a_480_297# a_608_49# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
.ends


******* EOF

** End of included library ./pdk/sky130_fd_sc_hd.spice

.subckt mgmt_protect caravel_clk caravel_clk2 caravel_rstn mprj_ack_i_core mprj_ack_i_user mprj_cyc_o_core mprj_cyc_o_user mprj_iena_wb mprj_stb_o_core mprj_stb_o_user mprj_we_o_core mprj_we_o_user user1_vcc_powergood user1_vdd_powergood user2_vcc_powergood user2_vdd_powergood user_clock user_clock2 user_reset vccd vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd vssd1 vssd2 la_data_in_core[0] la_data_in_core[1] la_data_in_core[2] la_data_in_core[3] la_data_in_core[4] la_data_in_core[5] la_data_in_core[6] la_data_in_core[7] la_data_in_core[8] la_data_in_core[9] la_data_in_core[10] la_data_in_core[11] la_data_in_core[12] la_data_in_core[13] la_data_in_core[14] la_data_in_core[15] la_data_in_core[16] la_data_in_core[17] la_data_in_core[18] la_data_in_core[19] la_data_in_core[20] la_data_in_core[21] la_data_in_core[22] la_data_in_core[23] la_data_in_core[24] la_data_in_core[25] la_data_in_core[26] la_data_in_core[27] la_data_in_core[28] la_data_in_core[29] la_data_in_core[30] la_data_in_core[31] la_data_in_core[32] la_data_in_core[33] la_data_in_core[34] la_data_in_core[35] la_data_in_core[36] la_data_in_core[37] la_data_in_core[38] la_data_in_core[39] la_data_in_core[40] la_data_in_core[41] la_data_in_core[42] la_data_in_core[43] la_data_in_core[44] la_data_in_core[45] la_data_in_core[46] la_data_in_core[47] la_data_in_core[48] la_data_in_core[49] la_data_in_core[50] la_data_in_core[51] la_data_in_core[52] la_data_in_core[53] la_data_in_core[54] la_data_in_core[55] la_data_in_core[56] la_data_in_core[57] la_data_in_core[58] la_data_in_core[59] la_data_in_core[60] la_data_in_core[61] la_data_in_core[62] la_data_in_core[63] la_data_in_core[64] la_data_in_core[65] la_data_in_core[66] la_data_in_core[67] la_data_in_core[68] la_data_in_core[69] la_data_in_core[70] la_data_in_core[71] la_data_in_core[72] la_data_in_core[73] la_data_in_core[74] la_data_in_core[75] la_data_in_core[76] la_data_in_core[77] la_data_in_core[78] la_data_in_core[79] la_data_in_core[80] la_data_in_core[81] la_data_in_core[82] la_data_in_core[83] la_data_in_core[84] la_data_in_core[85] la_data_in_core[86] la_data_in_core[87] la_data_in_core[88] la_data_in_core[89] la_data_in_core[90] la_data_in_core[91] la_data_in_core[92] la_data_in_core[93] la_data_in_core[94] la_data_in_core[95] la_data_in_core[96] la_data_in_core[97] la_data_in_core[98] la_data_in_core[99] la_data_in_core[100] la_data_in_core[101] la_data_in_core[102] la_data_in_core[103] la_data_in_core[104] la_data_in_core[105] la_data_in_core[106] la_data_in_core[107] la_data_in_core[108] la_data_in_core[109] la_data_in_core[110] la_data_in_core[111] la_data_in_core[112] la_data_in_core[113] la_data_in_core[114] la_data_in_core[115] la_data_in_core[116] la_data_in_core[117] la_data_in_core[118] la_data_in_core[119] la_data_in_core[120] la_data_in_core[121] la_data_in_core[122] la_data_in_core[123] la_data_in_core[124] la_data_in_core[125] la_data_in_core[126] la_data_in_core[127] la_data_in_mprj[0] la_data_in_mprj[1] la_data_in_mprj[2] la_data_in_mprj[3] la_data_in_mprj[4] la_data_in_mprj[5] la_data_in_mprj[6] la_data_in_mprj[7] la_data_in_mprj[8] la_data_in_mprj[9] la_data_in_mprj[10] la_data_in_mprj[11] la_data_in_mprj[12] la_data_in_mprj[13] la_data_in_mprj[14] la_data_in_mprj[15] la_data_in_mprj[16] la_data_in_mprj[17] la_data_in_mprj[18] la_data_in_mprj[19] la_data_in_mprj[20] la_data_in_mprj[21] la_data_in_mprj[22] la_data_in_mprj[23] la_data_in_mprj[24] la_data_in_mprj[25] la_data_in_mprj[26] la_data_in_mprj[27] la_data_in_mprj[28] la_data_in_mprj[29] la_data_in_mprj[30] la_data_in_mprj[31] la_data_in_mprj[32] la_data_in_mprj[33] la_data_in_mprj[34] la_data_in_mprj[35] la_data_in_mprj[36] la_data_in_mprj[37] la_data_in_mprj[38] la_data_in_mprj[39] la_data_in_mprj[40] la_data_in_mprj[41] la_data_in_mprj[42] la_data_in_mprj[43] la_data_in_mprj[44] la_data_in_mprj[45] la_data_in_mprj[46] la_data_in_mprj[47] la_data_in_mprj[48] la_data_in_mprj[49] la_data_in_mprj[50] la_data_in_mprj[51] la_data_in_mprj[52] la_data_in_mprj[53] la_data_in_mprj[54] la_data_in_mprj[55] la_data_in_mprj[56] la_data_in_mprj[57] la_data_in_mprj[58] la_data_in_mprj[59] la_data_in_mprj[60] la_data_in_mprj[61] la_data_in_mprj[62] la_data_in_mprj[63] la_data_in_mprj[64] la_data_in_mprj[65] la_data_in_mprj[66] la_data_in_mprj[67] la_data_in_mprj[68] la_data_in_mprj[69] la_data_in_mprj[70] la_data_in_mprj[71] la_data_in_mprj[72] la_data_in_mprj[73] la_data_in_mprj[74] la_data_in_mprj[75] la_data_in_mprj[76] la_data_in_mprj[77] la_data_in_mprj[78] la_data_in_mprj[79] la_data_in_mprj[80] la_data_in_mprj[81] la_data_in_mprj[82] la_data_in_mprj[83] la_data_in_mprj[84] la_data_in_mprj[85] la_data_in_mprj[86] la_data_in_mprj[87] la_data_in_mprj[88] la_data_in_mprj[89] la_data_in_mprj[90] la_data_in_mprj[91] la_data_in_mprj[92] la_data_in_mprj[93] la_data_in_mprj[94] la_data_in_mprj[95] la_data_in_mprj[96] la_data_in_mprj[97] la_data_in_mprj[98] la_data_in_mprj[99] la_data_in_mprj[100] la_data_in_mprj[101] la_data_in_mprj[102] la_data_in_mprj[103] la_data_in_mprj[104] la_data_in_mprj[105] la_data_in_mprj[106] la_data_in_mprj[107] la_data_in_mprj[108] la_data_in_mprj[109] la_data_in_mprj[110] la_data_in_mprj[111] la_data_in_mprj[112] la_data_in_mprj[113] la_data_in_mprj[114] la_data_in_mprj[115] la_data_in_mprj[116] la_data_in_mprj[117] la_data_in_mprj[118] la_data_in_mprj[119] la_data_in_mprj[120] la_data_in_mprj[121] la_data_in_mprj[122] la_data_in_mprj[123] la_data_in_mprj[124] la_data_in_mprj[125] la_data_in_mprj[126] la_data_in_mprj[127] la_data_out_core[0] la_data_out_core[1] la_data_out_core[2] la_data_out_core[3] la_data_out_core[4] la_data_out_core[5] la_data_out_core[6] la_data_out_core[7] la_data_out_core[8] la_data_out_core[9] la_data_out_core[10] la_data_out_core[11] la_data_out_core[12] la_data_out_core[13] la_data_out_core[14] la_data_out_core[15] la_data_out_core[16] la_data_out_core[17] la_data_out_core[18] la_data_out_core[19] la_data_out_core[20] la_data_out_core[21] la_data_out_core[22] la_data_out_core[23] la_data_out_core[24] la_data_out_core[25] la_data_out_core[26] la_data_out_core[27] la_data_out_core[28] la_data_out_core[29] la_data_out_core[30] la_data_out_core[31] la_data_out_core[32] la_data_out_core[33] la_data_out_core[34] la_data_out_core[35] la_data_out_core[36] la_data_out_core[37] la_data_out_core[38] la_data_out_core[39] la_data_out_core[40] la_data_out_core[41] la_data_out_core[42] la_data_out_core[43] la_data_out_core[44] la_data_out_core[45] la_data_out_core[46] la_data_out_core[47] la_data_out_core[48] la_data_out_core[49] la_data_out_core[50] la_data_out_core[51] la_data_out_core[52] la_data_out_core[53] la_data_out_core[54] la_data_out_core[55] la_data_out_core[56] la_data_out_core[57] la_data_out_core[58] la_data_out_core[59] la_data_out_core[60] la_data_out_core[61] la_data_out_core[62] la_data_out_core[63] la_data_out_core[64] la_data_out_core[65] la_data_out_core[66] la_data_out_core[67] la_data_out_core[68] la_data_out_core[69] la_data_out_core[70] la_data_out_core[71] la_data_out_core[72] la_data_out_core[73] la_data_out_core[74] la_data_out_core[75] la_data_out_core[76] la_data_out_core[77] la_data_out_core[78] la_data_out_core[79] la_data_out_core[80] la_data_out_core[81] la_data_out_core[82] la_data_out_core[83] la_data_out_core[84] la_data_out_core[85] la_data_out_core[86] la_data_out_core[87] la_data_out_core[88] la_data_out_core[89] la_data_out_core[90] la_data_out_core[91] la_data_out_core[92] la_data_out_core[93] la_data_out_core[94] la_data_out_core[95] la_data_out_core[96] la_data_out_core[97] la_data_out_core[98] la_data_out_core[99] la_data_out_core[100] la_data_out_core[101] la_data_out_core[102] la_data_out_core[103] la_data_out_core[104] la_data_out_core[105] la_data_out_core[106] la_data_out_core[107] la_data_out_core[108] la_data_out_core[109] la_data_out_core[110] la_data_out_core[111] la_data_out_core[112] la_data_out_core[113] la_data_out_core[114] la_data_out_core[115] la_data_out_core[116] la_data_out_core[117] la_data_out_core[118] la_data_out_core[119] la_data_out_core[120] la_data_out_core[121] la_data_out_core[122] la_data_out_core[123] la_data_out_core[124] la_data_out_core[125] la_data_out_core[126] la_data_out_core[127] la_data_out_mprj[0] la_data_out_mprj[1] la_data_out_mprj[2] la_data_out_mprj[3] la_data_out_mprj[4] la_data_out_mprj[5] la_data_out_mprj[6] la_data_out_mprj[7] la_data_out_mprj[8] la_data_out_mprj[9] la_data_out_mprj[10] la_data_out_mprj[11] la_data_out_mprj[12] la_data_out_mprj[13] la_data_out_mprj[14] la_data_out_mprj[15] la_data_out_mprj[16] la_data_out_mprj[17] la_data_out_mprj[18] la_data_out_mprj[19] la_data_out_mprj[20] la_data_out_mprj[21] la_data_out_mprj[22] la_data_out_mprj[23] la_data_out_mprj[24] la_data_out_mprj[25] la_data_out_mprj[26] la_data_out_mprj[27] la_data_out_mprj[28] la_data_out_mprj[29] la_data_out_mprj[30] la_data_out_mprj[31] la_data_out_mprj[32] la_data_out_mprj[33] la_data_out_mprj[34] la_data_out_mprj[35] la_data_out_mprj[36] la_data_out_mprj[37] la_data_out_mprj[38] la_data_out_mprj[39] la_data_out_mprj[40] la_data_out_mprj[41] la_data_out_mprj[42] la_data_out_mprj[43] la_data_out_mprj[44] la_data_out_mprj[45] la_data_out_mprj[46] la_data_out_mprj[47] la_data_out_mprj[48] la_data_out_mprj[49] la_data_out_mprj[50] la_data_out_mprj[51] la_data_out_mprj[52] la_data_out_mprj[53] la_data_out_mprj[54] la_data_out_mprj[55] la_data_out_mprj[56] la_data_out_mprj[57] la_data_out_mprj[58] la_data_out_mprj[59] la_data_out_mprj[60] la_data_out_mprj[61] la_data_out_mprj[62] la_data_out_mprj[63] la_data_out_mprj[64] la_data_out_mprj[65] la_data_out_mprj[66] la_data_out_mprj[67] la_data_out_mprj[68] la_data_out_mprj[69] la_data_out_mprj[70] la_data_out_mprj[71] la_data_out_mprj[72] la_data_out_mprj[73] la_data_out_mprj[74] la_data_out_mprj[75] la_data_out_mprj[76] la_data_out_mprj[77] la_data_out_mprj[78] la_data_out_mprj[79] la_data_out_mprj[80] la_data_out_mprj[81] la_data_out_mprj[82] la_data_out_mprj[83] la_data_out_mprj[84] la_data_out_mprj[85] la_data_out_mprj[86] la_data_out_mprj[87] la_data_out_mprj[88] la_data_out_mprj[89] la_data_out_mprj[90] la_data_out_mprj[91] la_data_out_mprj[92] la_data_out_mprj[93] la_data_out_mprj[94] la_data_out_mprj[95] la_data_out_mprj[96] la_data_out_mprj[97] la_data_out_mprj[98] la_data_out_mprj[99] la_data_out_mprj[100] la_data_out_mprj[101] la_data_out_mprj[102] la_data_out_mprj[103] la_data_out_mprj[104] la_data_out_mprj[105] la_data_out_mprj[106] la_data_out_mprj[107] la_data_out_mprj[108] la_data_out_mprj[109] la_data_out_mprj[110] la_data_out_mprj[111] la_data_out_mprj[112] la_data_out_mprj[113] la_data_out_mprj[114] la_data_out_mprj[115] la_data_out_mprj[116] la_data_out_mprj[117] la_data_out_mprj[118] la_data_out_mprj[119] la_data_out_mprj[120] la_data_out_mprj[121] la_data_out_mprj[122] la_data_out_mprj[123] la_data_out_mprj[124] la_data_out_mprj[125] la_data_out_mprj[126] la_data_out_mprj[127] la_iena_mprj[0] la_iena_mprj[1] la_iena_mprj[2] la_iena_mprj[3] la_iena_mprj[4] la_iena_mprj[5] la_iena_mprj[6] la_iena_mprj[7] la_iena_mprj[8] la_iena_mprj[9] la_iena_mprj[10] la_iena_mprj[11] la_iena_mprj[12] la_iena_mprj[13] la_iena_mprj[14] la_iena_mprj[15] la_iena_mprj[16] la_iena_mprj[17] la_iena_mprj[18] la_iena_mprj[19] la_iena_mprj[20] la_iena_mprj[21] la_iena_mprj[22] la_iena_mprj[23] la_iena_mprj[24] la_iena_mprj[25] la_iena_mprj[26] la_iena_mprj[27] la_iena_mprj[28] la_iena_mprj[29] la_iena_mprj[30] la_iena_mprj[31] la_iena_mprj[32] la_iena_mprj[33] la_iena_mprj[34] la_iena_mprj[35] la_iena_mprj[36] la_iena_mprj[37] la_iena_mprj[38] la_iena_mprj[39] la_iena_mprj[40] la_iena_mprj[41] la_iena_mprj[42] la_iena_mprj[43] la_iena_mprj[44] la_iena_mprj[45] la_iena_mprj[46] la_iena_mprj[47] la_iena_mprj[48] la_iena_mprj[49] la_iena_mprj[50] la_iena_mprj[51] la_iena_mprj[52] la_iena_mprj[53] la_iena_mprj[54] la_iena_mprj[55] la_iena_mprj[56] la_iena_mprj[57] la_iena_mprj[58] la_iena_mprj[59] la_iena_mprj[60] la_iena_mprj[61] la_iena_mprj[62] la_iena_mprj[63] la_iena_mprj[64] la_iena_mprj[65] la_iena_mprj[66] la_iena_mprj[67] la_iena_mprj[68] la_iena_mprj[69] la_iena_mprj[70] la_iena_mprj[71] la_iena_mprj[72] la_iena_mprj[73] la_iena_mprj[74] la_iena_mprj[75] la_iena_mprj[76] la_iena_mprj[77] la_iena_mprj[78] la_iena_mprj[79] la_iena_mprj[80] la_iena_mprj[81] la_iena_mprj[82] la_iena_mprj[83] la_iena_mprj[84] la_iena_mprj[85] la_iena_mprj[86] la_iena_mprj[87] la_iena_mprj[88] la_iena_mprj[89] la_iena_mprj[90] la_iena_mprj[91] la_iena_mprj[92] la_iena_mprj[93] la_iena_mprj[94] la_iena_mprj[95] la_iena_mprj[96] la_iena_mprj[97] la_iena_mprj[98] la_iena_mprj[99] la_iena_mprj[100] la_iena_mprj[101] la_iena_mprj[102] la_iena_mprj[103] la_iena_mprj[104] la_iena_mprj[105] la_iena_mprj[106] la_iena_mprj[107] la_iena_mprj[108] la_iena_mprj[109] la_iena_mprj[110] la_iena_mprj[111] la_iena_mprj[112] la_iena_mprj[113] la_iena_mprj[114] la_iena_mprj[115] la_iena_mprj[116] la_iena_mprj[117] la_iena_mprj[118] la_iena_mprj[119] la_iena_mprj[120] la_iena_mprj[121] la_iena_mprj[122] la_iena_mprj[123] la_iena_mprj[124] la_iena_mprj[125] la_iena_mprj[126] la_iena_mprj[127] la_oenb_core[0] la_oenb_core[1] la_oenb_core[2] la_oenb_core[3] la_oenb_core[4] la_oenb_core[5] la_oenb_core[6] la_oenb_core[7] la_oenb_core[8] la_oenb_core[9] la_oenb_core[10] la_oenb_core[11] la_oenb_core[12] la_oenb_core[13] la_oenb_core[14] la_oenb_core[15] la_oenb_core[16] la_oenb_core[17] la_oenb_core[18] la_oenb_core[19] la_oenb_core[20] la_oenb_core[21] la_oenb_core[22] la_oenb_core[23] la_oenb_core[24] la_oenb_core[25] la_oenb_core[26] la_oenb_core[27] la_oenb_core[28] la_oenb_core[29] la_oenb_core[30] la_oenb_core[31] la_oenb_core[32] la_oenb_core[33] la_oenb_core[34] la_oenb_core[35] la_oenb_core[36] la_oenb_core[37] la_oenb_core[38] la_oenb_core[39] la_oenb_core[40] la_oenb_core[41] la_oenb_core[42] la_oenb_core[43] la_oenb_core[44] la_oenb_core[45] la_oenb_core[46] la_oenb_core[47] la_oenb_core[48] la_oenb_core[49] la_oenb_core[50] la_oenb_core[51] la_oenb_core[52] la_oenb_core[53] la_oenb_core[54] la_oenb_core[55] la_oenb_core[56] la_oenb_core[57] la_oenb_core[58] la_oenb_core[59] la_oenb_core[60] la_oenb_core[61] la_oenb_core[62] la_oenb_core[63] la_oenb_core[64] la_oenb_core[65] la_oenb_core[66] la_oenb_core[67] la_oenb_core[68] la_oenb_core[69] la_oenb_core[70] la_oenb_core[71] la_oenb_core[72] la_oenb_core[73] la_oenb_core[74] la_oenb_core[75] la_oenb_core[76] la_oenb_core[77] la_oenb_core[78] la_oenb_core[79] la_oenb_core[80] la_oenb_core[81] la_oenb_core[82] la_oenb_core[83] la_oenb_core[84] la_oenb_core[85] la_oenb_core[86] la_oenb_core[87] la_oenb_core[88] la_oenb_core[89] la_oenb_core[90] la_oenb_core[91] la_oenb_core[92] la_oenb_core[93] la_oenb_core[94] la_oenb_core[95] la_oenb_core[96] la_oenb_core[97] la_oenb_core[98] la_oenb_core[99] la_oenb_core[100] la_oenb_core[101] la_oenb_core[102] la_oenb_core[103] la_oenb_core[104] la_oenb_core[105] la_oenb_core[106] la_oenb_core[107] la_oenb_core[108] la_oenb_core[109] la_oenb_core[110] la_oenb_core[111] la_oenb_core[112] la_oenb_core[113] la_oenb_core[114] la_oenb_core[115] la_oenb_core[116] la_oenb_core[117] la_oenb_core[118] la_oenb_core[119] la_oenb_core[120] la_oenb_core[121] la_oenb_core[122] la_oenb_core[123] la_oenb_core[124] la_oenb_core[125] la_oenb_core[126] la_oenb_core[127] la_oenb_mprj[0] la_oenb_mprj[1] la_oenb_mprj[2] la_oenb_mprj[3] la_oenb_mprj[4] la_oenb_mprj[5] la_oenb_mprj[6] la_oenb_mprj[7] la_oenb_mprj[8] la_oenb_mprj[9] la_oenb_mprj[10] la_oenb_mprj[11] la_oenb_mprj[12] la_oenb_mprj[13] la_oenb_mprj[14] la_oenb_mprj[15] la_oenb_mprj[16] la_oenb_mprj[17] la_oenb_mprj[18] la_oenb_mprj[19] la_oenb_mprj[20] la_oenb_mprj[21] la_oenb_mprj[22] la_oenb_mprj[23] la_oenb_mprj[24] la_oenb_mprj[25] la_oenb_mprj[26] la_oenb_mprj[27] la_oenb_mprj[28] la_oenb_mprj[29] la_oenb_mprj[30] la_oenb_mprj[31] la_oenb_mprj[32] la_oenb_mprj[33] la_oenb_mprj[34] la_oenb_mprj[35] la_oenb_mprj[36] la_oenb_mprj[37] la_oenb_mprj[38] la_oenb_mprj[39] la_oenb_mprj[40] la_oenb_mprj[41] la_oenb_mprj[42] la_oenb_mprj[43] la_oenb_mprj[44] la_oenb_mprj[45] la_oenb_mprj[46] la_oenb_mprj[47] la_oenb_mprj[48] la_oenb_mprj[49] la_oenb_mprj[50] la_oenb_mprj[51] la_oenb_mprj[52] la_oenb_mprj[53] la_oenb_mprj[54] la_oenb_mprj[55] la_oenb_mprj[56] la_oenb_mprj[57] la_oenb_mprj[58] la_oenb_mprj[59] la_oenb_mprj[60] la_oenb_mprj[61] la_oenb_mprj[62] la_oenb_mprj[63] la_oenb_mprj[64] la_oenb_mprj[65] la_oenb_mprj[66] la_oenb_mprj[67] la_oenb_mprj[68] la_oenb_mprj[69] la_oenb_mprj[70] la_oenb_mprj[71] la_oenb_mprj[72] la_oenb_mprj[73] la_oenb_mprj[74] la_oenb_mprj[75] la_oenb_mprj[76] la_oenb_mprj[77] la_oenb_mprj[78] la_oenb_mprj[79] la_oenb_mprj[80] la_oenb_mprj[81] la_oenb_mprj[82] la_oenb_mprj[83] la_oenb_mprj[84] la_oenb_mprj[85] la_oenb_mprj[86] la_oenb_mprj[87] la_oenb_mprj[88] la_oenb_mprj[89] la_oenb_mprj[90] la_oenb_mprj[91] la_oenb_mprj[92] la_oenb_mprj[93] la_oenb_mprj[94] la_oenb_mprj[95] la_oenb_mprj[96] la_oenb_mprj[97] la_oenb_mprj[98] la_oenb_mprj[99] la_oenb_mprj[100] la_oenb_mprj[101] la_oenb_mprj[102] la_oenb_mprj[103] la_oenb_mprj[104] la_oenb_mprj[105] la_oenb_mprj[106] la_oenb_mprj[107] la_oenb_mprj[108] la_oenb_mprj[109] la_oenb_mprj[110] la_oenb_mprj[111] la_oenb_mprj[112] la_oenb_mprj[113] la_oenb_mprj[114] la_oenb_mprj[115] la_oenb_mprj[116] la_oenb_mprj[117] la_oenb_mprj[118] la_oenb_mprj[119] la_oenb_mprj[120] la_oenb_mprj[121] la_oenb_mprj[122] la_oenb_mprj[123] la_oenb_mprj[124] la_oenb_mprj[125] la_oenb_mprj[126] la_oenb_mprj[127] mprj_adr_o_core[0] mprj_adr_o_core[1] mprj_adr_o_core[2] mprj_adr_o_core[3] mprj_adr_o_core[4] mprj_adr_o_core[5] mprj_adr_o_core[6] mprj_adr_o_core[7] mprj_adr_o_core[8] mprj_adr_o_core[9] mprj_adr_o_core[10] mprj_adr_o_core[11] mprj_adr_o_core[12] mprj_adr_o_core[13] mprj_adr_o_core[14] mprj_adr_o_core[15] mprj_adr_o_core[16] mprj_adr_o_core[17] mprj_adr_o_core[18] mprj_adr_o_core[19] mprj_adr_o_core[20] mprj_adr_o_core[21] mprj_adr_o_core[22] mprj_adr_o_core[23] mprj_adr_o_core[24] mprj_adr_o_core[25] mprj_adr_o_core[26] mprj_adr_o_core[27] mprj_adr_o_core[28] mprj_adr_o_core[29] mprj_adr_o_core[30] mprj_adr_o_core[31] mprj_adr_o_user[0] mprj_adr_o_user[1] mprj_adr_o_user[2] mprj_adr_o_user[3] mprj_adr_o_user[4] mprj_adr_o_user[5] mprj_adr_o_user[6] mprj_adr_o_user[7] mprj_adr_o_user[8] mprj_adr_o_user[9] mprj_adr_o_user[10] mprj_adr_o_user[11] mprj_adr_o_user[12] mprj_adr_o_user[13] mprj_adr_o_user[14] mprj_adr_o_user[15] mprj_adr_o_user[16] mprj_adr_o_user[17] mprj_adr_o_user[18] mprj_adr_o_user[19] mprj_adr_o_user[20] mprj_adr_o_user[21] mprj_adr_o_user[22] mprj_adr_o_user[23] mprj_adr_o_user[24] mprj_adr_o_user[25] mprj_adr_o_user[26] mprj_adr_o_user[27] mprj_adr_o_user[28] mprj_adr_o_user[29] mprj_adr_o_user[30] mprj_adr_o_user[31] mprj_dat_i_core[0] mprj_dat_i_core[1] mprj_dat_i_core[2] mprj_dat_i_core[3] mprj_dat_i_core[4] mprj_dat_i_core[5] mprj_dat_i_core[6] mprj_dat_i_core[7] mprj_dat_i_core[8] mprj_dat_i_core[9] mprj_dat_i_core[10] mprj_dat_i_core[11] mprj_dat_i_core[12] mprj_dat_i_core[13] mprj_dat_i_core[14] mprj_dat_i_core[15] mprj_dat_i_core[16] mprj_dat_i_core[17] mprj_dat_i_core[18] mprj_dat_i_core[19] mprj_dat_i_core[20] mprj_dat_i_core[21] mprj_dat_i_core[22] mprj_dat_i_core[23] mprj_dat_i_core[24] mprj_dat_i_core[25] mprj_dat_i_core[26] mprj_dat_i_core[27] mprj_dat_i_core[28] mprj_dat_i_core[29] mprj_dat_i_core[30] mprj_dat_i_core[31] mprj_dat_i_user[0] mprj_dat_i_user[1] mprj_dat_i_user[2] mprj_dat_i_user[3] mprj_dat_i_user[4] mprj_dat_i_user[5] mprj_dat_i_user[6] mprj_dat_i_user[7] mprj_dat_i_user[8] mprj_dat_i_user[9] mprj_dat_i_user[10] mprj_dat_i_user[11] mprj_dat_i_user[12] mprj_dat_i_user[13] mprj_dat_i_user[14] mprj_dat_i_user[15] mprj_dat_i_user[16] mprj_dat_i_user[17] mprj_dat_i_user[18] mprj_dat_i_user[19] mprj_dat_i_user[20] mprj_dat_i_user[21] mprj_dat_i_user[22] mprj_dat_i_user[23] mprj_dat_i_user[24] mprj_dat_i_user[25] mprj_dat_i_user[26] mprj_dat_i_user[27] mprj_dat_i_user[28] mprj_dat_i_user[29] mprj_dat_i_user[30] mprj_dat_i_user[31] mprj_dat_o_core[0] mprj_dat_o_core[1] mprj_dat_o_core[2] mprj_dat_o_core[3] mprj_dat_o_core[4] mprj_dat_o_core[5] mprj_dat_o_core[6] mprj_dat_o_core[7] mprj_dat_o_core[8] mprj_dat_o_core[9] mprj_dat_o_core[10] mprj_dat_o_core[11] mprj_dat_o_core[12] mprj_dat_o_core[13] mprj_dat_o_core[14] mprj_dat_o_core[15] mprj_dat_o_core[16] mprj_dat_o_core[17] mprj_dat_o_core[18] mprj_dat_o_core[19] mprj_dat_o_core[20] mprj_dat_o_core[21] mprj_dat_o_core[22] mprj_dat_o_core[23] mprj_dat_o_core[24] mprj_dat_o_core[25] mprj_dat_o_core[26] mprj_dat_o_core[27] mprj_dat_o_core[28] mprj_dat_o_core[29] mprj_dat_o_core[30] mprj_dat_o_core[31] mprj_dat_o_user[0] mprj_dat_o_user[1] mprj_dat_o_user[2] mprj_dat_o_user[3] mprj_dat_o_user[4] mprj_dat_o_user[5] mprj_dat_o_user[6] mprj_dat_o_user[7] mprj_dat_o_user[8] mprj_dat_o_user[9] mprj_dat_o_user[10] mprj_dat_o_user[11] mprj_dat_o_user[12] mprj_dat_o_user[13] mprj_dat_o_user[14] mprj_dat_o_user[15] mprj_dat_o_user[16] mprj_dat_o_user[17] mprj_dat_o_user[18] mprj_dat_o_user[19] mprj_dat_o_user[20] mprj_dat_o_user[21] mprj_dat_o_user[22] mprj_dat_o_user[23] mprj_dat_o_user[24] mprj_dat_o_user[25] mprj_dat_o_user[26] mprj_dat_o_user[27] mprj_dat_o_user[28] mprj_dat_o_user[29] mprj_dat_o_user[30] mprj_dat_o_user[31] mprj_sel_o_core[0] mprj_sel_o_core[1] mprj_sel_o_core[2] mprj_sel_o_core[3] mprj_sel_o_user[0] mprj_sel_o_user[1] mprj_sel_o_user[2] mprj_sel_o_user[3] user_irq[0] user_irq[1] user_irq[2] user_irq_core[0] user_irq_core[1] user_irq_core[2] user_irq_ena[0] user_irq_ena[1] user_irq_ena[2] 

XANTENNA__329__A net478 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__330__A net479 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__331__A net480 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__332__A net481 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__333__A net483 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__334__A net484 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__335__A net485 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__336__A net486 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__337__A net487 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__338__A net488 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__339__A net489 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__340__A net490 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__341__A net491 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__342__A net492 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__343__A net494 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__344__A net495 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__345__A net496 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__346__A net497 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__347__A net498 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__348__A net499 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__349__A net500 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__350__A net501 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__351__A net502 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__352__A net503 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__353__A net505 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__354__A net506 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__355__A net507 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__356__A net508 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__357__A net509 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__358__A net510 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__359__A net511 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__360__A net512 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__361__A net513 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__362__A net514 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__363__A net389 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__364__A net390 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__365__A net391 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__366__A net392 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__367__A net393 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__368__A net394 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__369__A net395 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__370__A net396 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__371__A net397 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__372__A net398 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__373__A net400 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__374__A net401 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__375__A net402 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__376__A net403 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__377__A net404 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__378__A net405 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__379__A net406 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__380__A net407 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__381__A net408 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__382__A net409 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__383__A net411 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__384__A net412 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__385__A net413 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__386__A net414 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__387__A net415 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__388__A net416 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__389__A net417 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__390__A net418 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__391__A net1 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__392__A net2 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__393__A net549 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__394__A net619 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__395__A net620 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__396__A net615 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__397__A net616 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__398__A net617 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__399__A net618 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__400__A net517 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__401__A net528 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__402__A net539 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__403__A net542 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__404__A net543 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__405__A net544 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__406__A net545 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__407__A net546 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__408__A net547 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__409__A net548 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__410__A net518 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__411__A net519 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__412__A net520 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__413__A net521 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__414__A net522 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__415__A net523 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__416__A net524 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__417__A net525 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__418__A net526 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__419__A net527 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__420__A net529 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__421__A net530 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__422__A net531 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__423__A net532 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__424__A net533 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__425__A net534 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__426__A net535 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__427__A net536 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__428__A net537 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__429__A net538 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__430__A net540 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__431__A net541 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__432__A net582 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__433__A net593 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__434__A net604 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__435__A net607 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__436__A net608 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__437__A net609 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__438__A net610 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__439__A net611 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__440__A net612 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__441__A net613 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__442__A net583 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__443__A net584 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__444__A net585 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__445__A net586 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__446__A net587 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__447__A net588 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__448__A net589 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__449__A net590 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__450__A net591 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__451__A net592 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__452__A net594 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__453__A net595 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__454__A net596 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__455__A net597 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__456__A net598 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__457__A net599 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__458__A net600 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__459__A net601 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__460__A net602 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__461__A net603 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__462__A net605 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__463__A net606 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__464__A net132 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__465__A net171 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__466__A net182 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__467__A net193 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__468__A net204 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__469__A net215 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__470__A net226 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__471__A net237 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__472__A net248 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__473__A net259 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__474__A net143 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__475__A net154 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__476__A net163 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__477__A net164 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__478__A net165 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__479__A net166 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__480__A net167 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__481__A net168 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__482__A net169 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__483__A net170 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__484__A net172 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__485__A net173 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__486__A net174 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__487__A net175 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__488__A net176 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__489__A net177 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__490__A net178 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__491__A net179 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__492__A net180 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__493__A net181 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__494__A net183 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__495__A net184 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__496__A net185 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__497__A net186 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__498__A net187 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__499__A net188 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__500__A net189 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__501__A net190 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__502__A net191 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__503__A net192 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__504__A net194 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__505__A net195 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__506__A net196 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__507__A net197 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__508__A net198 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__509__A net199 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__510__A net200 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__511__A net201 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__512__A net202 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__513__A net203 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__514__A net205 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__515__A net206 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__516__A net207 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__517__A net208 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__518__A net209 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__519__A net210 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__520__A net211 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__521__A net212 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__522__A net213 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__523__A net214 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__524__A net216 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__525__A net217 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__526__A net218 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__527__A net219 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__528__A net220 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__529__A net221 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__530__A net222 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__531__A net223 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__532__A net224 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__533__A net225 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__534__A net227 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__535__A net228 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__536__A net229 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__537__A net230 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__538__A net231 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__539__A net232 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__540__A net233 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__541__A net234 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__542__A net235 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__543__A net236 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__544__A net238 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__545__A net239 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__546__A net240 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__547__A net241 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__548__A net242 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__549__A net243 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__550__A net244 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__551__A net245 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__552__A net246 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__553__A net247 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__554__A net249 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__555__A net250 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__556__A net251 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__557__A net252 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__558__A net253 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__559__A net254 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__560__A net255 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__561__A net256 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__562__A net257 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__563__A net258 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__564__A net133 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__565__A net134 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__566__A net135 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__567__A net136 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__568__A net137 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__569__A net138 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__570__A net139 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__571__A net140 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__572__A net141 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__573__A net142 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__574__A net144 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__575__A net145 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__576__A net146 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__577__A net147 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__578__A net148 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__579__A net149 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__580__A net150 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__581__A net151 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__582__A net152 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__583__A net153 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__584__A net155 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__585__A net156 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__586__A net157 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__587__A net158 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__588__A net159 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__589__A net160 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__590__A net161 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__591__A net162 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__592__A net388 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__593__A net427 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__594__A net438 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__595__A net449 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__596__A net460 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__597__A net471 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__598__A net482 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__599__A net493 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__600__A net504 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__601__A net515 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__602__A net399 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__603__A net410 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__604__A net419 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__605__A net420 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__606__A net421 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__607__A net422 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__608__A net423 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__609__A net424 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__610__A net425 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__611__A net426 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__612__A net428 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__613__A net429 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__614__A net430 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__615__A net431 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__616__A net432 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__617__A net433 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__618__A net434 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__619__A net435 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__620__A net436 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__621__A net437 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__622__A net439 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__623__A net440 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__624__A net441 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__625__A net442 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__626__A net443 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__627__A net444 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__628__A net445 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__629__A net446 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__630__A net447 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__631__A net448 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__632__A net450 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__633__A net451 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__634__A net452 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__635__A net453 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__636__A net454 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__637__A net455 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__638__A net456 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__639__A net457 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__640__A net458 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__641__A net459 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__642__A net461 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__643__A net462 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__644__A net463 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__645__A net464 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__646__A net465 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__647__A net466 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__648__A net467 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__649__A net468 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__650__A net469 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__651__A net470 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__652__A net472 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__653__A net473 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__654__A net474 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__655__A net475 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__656__A net476 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__657__A net477 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input100_A la_data_out_core[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input101_A la_data_out_core[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input102_A la_data_out_core[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input103_A la_data_out_core[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input104_A la_data_out_core[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input105_A la_data_out_core[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input106_A la_data_out_core[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input107_A la_data_out_core[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input108_A la_data_out_core[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input109_A la_data_out_core[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input10_A la_data_out_core[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input110_A la_data_out_core[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input111_A la_data_out_core[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input112_A la_data_out_core[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input113_A la_data_out_core[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input114_A la_data_out_core[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input115_A la_data_out_core[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input116_A la_data_out_core[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input117_A la_data_out_core[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input118_A la_data_out_core[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input119_A la_data_out_core[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input11_A la_data_out_core[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input120_A la_data_out_core[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input121_A la_data_out_core[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input122_A la_data_out_core[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input123_A la_data_out_core[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input124_A la_data_out_core[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input125_A la_data_out_core[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input126_A la_data_out_core[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input127_A la_data_out_core[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input128_A la_data_out_core[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input129_A la_data_out_core[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input12_A la_data_out_core[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input130_A la_data_out_core[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input131_A la_data_out_core[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input132_A la_data_out_mprj[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input133_A la_data_out_mprj[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input134_A la_data_out_mprj[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input135_A la_data_out_mprj[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input136_A la_data_out_mprj[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input137_A la_data_out_mprj[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input138_A la_data_out_mprj[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input139_A la_data_out_mprj[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input13_A la_data_out_core[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input140_A la_data_out_mprj[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input141_A la_data_out_mprj[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input142_A la_data_out_mprj[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input143_A la_data_out_mprj[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input144_A la_data_out_mprj[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input145_A la_data_out_mprj[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input146_A la_data_out_mprj[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input147_A la_data_out_mprj[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input148_A la_data_out_mprj[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input149_A la_data_out_mprj[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input14_A la_data_out_core[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input150_A la_data_out_mprj[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input151_A la_data_out_mprj[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input152_A la_data_out_mprj[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input153_A la_data_out_mprj[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input154_A la_data_out_mprj[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input155_A la_data_out_mprj[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input156_A la_data_out_mprj[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input157_A la_data_out_mprj[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input158_A la_data_out_mprj[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input159_A la_data_out_mprj[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input15_A la_data_out_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input160_A la_data_out_mprj[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input161_A la_data_out_mprj[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input162_A la_data_out_mprj[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input163_A la_data_out_mprj[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input164_A la_data_out_mprj[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input165_A la_data_out_mprj[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input166_A la_data_out_mprj[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input167_A la_data_out_mprj[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input168_A la_data_out_mprj[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input169_A la_data_out_mprj[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input16_A la_data_out_core[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input170_A la_data_out_mprj[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input171_A la_data_out_mprj[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input172_A la_data_out_mprj[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input173_A la_data_out_mprj[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input174_A la_data_out_mprj[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input175_A la_data_out_mprj[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input176_A la_data_out_mprj[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input177_A la_data_out_mprj[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input178_A la_data_out_mprj[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input179_A la_data_out_mprj[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input17_A la_data_out_core[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input180_A la_data_out_mprj[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input181_A la_data_out_mprj[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input182_A la_data_out_mprj[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input183_A la_data_out_mprj[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input184_A la_data_out_mprj[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input185_A la_data_out_mprj[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input186_A la_data_out_mprj[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input187_A la_data_out_mprj[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input188_A la_data_out_mprj[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input189_A la_data_out_mprj[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input18_A la_data_out_core[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input190_A la_data_out_mprj[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input191_A la_data_out_mprj[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input192_A la_data_out_mprj[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input193_A la_data_out_mprj[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input194_A la_data_out_mprj[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input195_A la_data_out_mprj[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input196_A la_data_out_mprj[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input197_A la_data_out_mprj[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input198_A la_data_out_mprj[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input199_A la_data_out_mprj[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input19_A la_data_out_core[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input1_A caravel_clk vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input200_A la_data_out_mprj[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input201_A la_data_out_mprj[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input202_A la_data_out_mprj[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input203_A la_data_out_mprj[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input204_A la_data_out_mprj[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input205_A la_data_out_mprj[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input206_A la_data_out_mprj[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input207_A la_data_out_mprj[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input208_A la_data_out_mprj[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input209_A la_data_out_mprj[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input20_A la_data_out_core[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input210_A la_data_out_mprj[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input211_A la_data_out_mprj[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input212_A la_data_out_mprj[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input213_A la_data_out_mprj[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input214_A la_data_out_mprj[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input215_A la_data_out_mprj[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input216_A la_data_out_mprj[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input217_A la_data_out_mprj[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input218_A la_data_out_mprj[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input219_A la_data_out_mprj[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input21_A la_data_out_core[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input220_A la_data_out_mprj[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input221_A la_data_out_mprj[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input222_A la_data_out_mprj[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input223_A la_data_out_mprj[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input224_A la_data_out_mprj[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input225_A la_data_out_mprj[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input226_A la_data_out_mprj[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input227_A la_data_out_mprj[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input228_A la_data_out_mprj[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input229_A la_data_out_mprj[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input22_A la_data_out_core[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input230_A la_data_out_mprj[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input231_A la_data_out_mprj[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input232_A la_data_out_mprj[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input233_A la_data_out_mprj[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input234_A la_data_out_mprj[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input235_A la_data_out_mprj[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input236_A la_data_out_mprj[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input237_A la_data_out_mprj[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input238_A la_data_out_mprj[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input239_A la_data_out_mprj[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input23_A la_data_out_core[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input240_A la_data_out_mprj[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input241_A la_data_out_mprj[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input242_A la_data_out_mprj[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input243_A la_data_out_mprj[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input244_A la_data_out_mprj[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input245_A la_data_out_mprj[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input246_A la_data_out_mprj[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input247_A la_data_out_mprj[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input248_A la_data_out_mprj[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input249_A la_data_out_mprj[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input24_A la_data_out_core[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input250_A la_data_out_mprj[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input251_A la_data_out_mprj[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input252_A la_data_out_mprj[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input253_A la_data_out_mprj[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input254_A la_data_out_mprj[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input255_A la_data_out_mprj[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input256_A la_data_out_mprj[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input257_A la_data_out_mprj[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input258_A la_data_out_mprj[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input259_A la_data_out_mprj[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input25_A la_data_out_core[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input260_A la_iena_mprj[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input261_A la_iena_mprj[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input262_A la_iena_mprj[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input263_A la_iena_mprj[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input264_A la_iena_mprj[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input265_A la_iena_mprj[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input266_A la_iena_mprj[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input267_A la_iena_mprj[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input268_A la_iena_mprj[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input269_A la_iena_mprj[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input26_A la_data_out_core[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input270_A la_iena_mprj[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input271_A la_iena_mprj[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input272_A la_iena_mprj[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input273_A la_iena_mprj[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input274_A la_iena_mprj[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input275_A la_iena_mprj[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input276_A la_iena_mprj[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input277_A la_iena_mprj[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input278_A la_iena_mprj[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input279_A la_iena_mprj[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input27_A la_data_out_core[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input280_A la_iena_mprj[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input281_A la_iena_mprj[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input282_A la_iena_mprj[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input283_A la_iena_mprj[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input284_A la_iena_mprj[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input285_A la_iena_mprj[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input286_A la_iena_mprj[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input287_A la_iena_mprj[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input288_A la_iena_mprj[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input289_A la_iena_mprj[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input28_A la_data_out_core[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input290_A la_iena_mprj[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input291_A la_iena_mprj[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input292_A la_iena_mprj[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input293_A la_iena_mprj[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input294_A la_iena_mprj[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input295_A la_iena_mprj[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input296_A la_iena_mprj[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input297_A la_iena_mprj[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input298_A la_iena_mprj[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input299_A la_iena_mprj[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input29_A la_data_out_core[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input2_A caravel_clk2 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input300_A la_iena_mprj[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input301_A la_iena_mprj[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input302_A la_iena_mprj[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input303_A la_iena_mprj[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input304_A la_iena_mprj[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input305_A la_iena_mprj[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input306_A la_iena_mprj[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input307_A la_iena_mprj[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input308_A la_iena_mprj[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input309_A la_iena_mprj[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input30_A la_data_out_core[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input310_A la_iena_mprj[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input311_A la_iena_mprj[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input312_A la_iena_mprj[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input313_A la_iena_mprj[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input314_A la_iena_mprj[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input315_A la_iena_mprj[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input316_A la_iena_mprj[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input317_A la_iena_mprj[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input318_A la_iena_mprj[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input319_A la_iena_mprj[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input31_A la_data_out_core[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input320_A la_iena_mprj[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input321_A la_iena_mprj[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input322_A la_iena_mprj[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input323_A la_iena_mprj[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input324_A la_iena_mprj[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input325_A la_iena_mprj[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input326_A la_iena_mprj[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input327_A la_iena_mprj[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input328_A la_iena_mprj[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input329_A la_iena_mprj[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input32_A la_data_out_core[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input330_A la_iena_mprj[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input331_A la_iena_mprj[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input332_A la_iena_mprj[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input333_A la_iena_mprj[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input334_A la_iena_mprj[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input335_A la_iena_mprj[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input336_A la_iena_mprj[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input337_A la_iena_mprj[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input338_A la_iena_mprj[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input339_A la_iena_mprj[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input33_A la_data_out_core[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input340_A la_iena_mprj[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input341_A la_iena_mprj[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input342_A la_iena_mprj[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input343_A la_iena_mprj[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input344_A la_iena_mprj[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input345_A la_iena_mprj[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input346_A la_iena_mprj[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input347_A la_iena_mprj[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input348_A la_iena_mprj[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input349_A la_iena_mprj[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input34_A la_data_out_core[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input350_A la_iena_mprj[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input351_A la_iena_mprj[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input352_A la_iena_mprj[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input353_A la_iena_mprj[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input354_A la_iena_mprj[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input355_A la_iena_mprj[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input356_A la_iena_mprj[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input357_A la_iena_mprj[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input358_A la_iena_mprj[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input359_A la_iena_mprj[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input35_A la_data_out_core[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input360_A la_iena_mprj[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input361_A la_iena_mprj[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input362_A la_iena_mprj[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input363_A la_iena_mprj[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input364_A la_iena_mprj[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input365_A la_iena_mprj[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input366_A la_iena_mprj[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input367_A la_iena_mprj[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input368_A la_iena_mprj[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input369_A la_iena_mprj[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input36_A la_data_out_core[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input370_A la_iena_mprj[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input371_A la_iena_mprj[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input372_A la_iena_mprj[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input373_A la_iena_mprj[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input374_A la_iena_mprj[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input375_A la_iena_mprj[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input376_A la_iena_mprj[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input377_A la_iena_mprj[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input378_A la_iena_mprj[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input379_A la_iena_mprj[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input37_A la_data_out_core[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input380_A la_iena_mprj[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input381_A la_iena_mprj[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input382_A la_iena_mprj[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input383_A la_iena_mprj[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input384_A la_iena_mprj[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input385_A la_iena_mprj[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input386_A la_iena_mprj[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input387_A la_iena_mprj[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input388_A la_oenb_mprj[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input389_A la_oenb_mprj[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input38_A la_data_out_core[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input390_A la_oenb_mprj[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input391_A la_oenb_mprj[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input392_A la_oenb_mprj[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input393_A la_oenb_mprj[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input394_A la_oenb_mprj[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input395_A la_oenb_mprj[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input396_A la_oenb_mprj[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input397_A la_oenb_mprj[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input398_A la_oenb_mprj[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input399_A la_oenb_mprj[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input39_A la_data_out_core[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input3_A caravel_rstn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input400_A la_oenb_mprj[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input401_A la_oenb_mprj[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input402_A la_oenb_mprj[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input403_A la_oenb_mprj[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input404_A la_oenb_mprj[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input405_A la_oenb_mprj[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input406_A la_oenb_mprj[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input407_A la_oenb_mprj[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input408_A la_oenb_mprj[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input409_A la_oenb_mprj[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input40_A la_data_out_core[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input410_A la_oenb_mprj[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input411_A la_oenb_mprj[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input412_A la_oenb_mprj[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input413_A la_oenb_mprj[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input414_A la_oenb_mprj[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input415_A la_oenb_mprj[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input416_A la_oenb_mprj[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input417_A la_oenb_mprj[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input418_A la_oenb_mprj[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input419_A la_oenb_mprj[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input41_A la_data_out_core[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input420_A la_oenb_mprj[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input421_A la_oenb_mprj[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input422_A la_oenb_mprj[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input423_A la_oenb_mprj[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input424_A la_oenb_mprj[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input425_A la_oenb_mprj[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input426_A la_oenb_mprj[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input427_A la_oenb_mprj[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input428_A la_oenb_mprj[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input429_A la_oenb_mprj[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input42_A la_data_out_core[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input430_A la_oenb_mprj[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input431_A la_oenb_mprj[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input432_A la_oenb_mprj[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input433_A la_oenb_mprj[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input434_A la_oenb_mprj[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input435_A la_oenb_mprj[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input436_A la_oenb_mprj[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input437_A la_oenb_mprj[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input438_A la_oenb_mprj[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input439_A la_oenb_mprj[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input43_A la_data_out_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input440_A la_oenb_mprj[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input441_A la_oenb_mprj[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input442_A la_oenb_mprj[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input443_A la_oenb_mprj[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input444_A la_oenb_mprj[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input445_A la_oenb_mprj[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input446_A la_oenb_mprj[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input447_A la_oenb_mprj[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input448_A la_oenb_mprj[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input449_A la_oenb_mprj[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input44_A la_data_out_core[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input450_A la_oenb_mprj[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input451_A la_oenb_mprj[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input452_A la_oenb_mprj[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input453_A la_oenb_mprj[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input454_A la_oenb_mprj[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input455_A la_oenb_mprj[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input456_A la_oenb_mprj[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input457_A la_oenb_mprj[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input458_A la_oenb_mprj[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input459_A la_oenb_mprj[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input45_A la_data_out_core[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input460_A la_oenb_mprj[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input461_A la_oenb_mprj[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input462_A la_oenb_mprj[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input463_A la_oenb_mprj[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input464_A la_oenb_mprj[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input465_A la_oenb_mprj[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input466_A la_oenb_mprj[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input467_A la_oenb_mprj[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input468_A la_oenb_mprj[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input469_A la_oenb_mprj[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input46_A la_data_out_core[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input470_A la_oenb_mprj[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input471_A la_oenb_mprj[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input472_A la_oenb_mprj[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input473_A la_oenb_mprj[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input474_A la_oenb_mprj[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input475_A la_oenb_mprj[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input476_A la_oenb_mprj[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input477_A la_oenb_mprj[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input478_A la_oenb_mprj[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input479_A la_oenb_mprj[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input47_A la_data_out_core[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input480_A la_oenb_mprj[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input481_A la_oenb_mprj[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input482_A la_oenb_mprj[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input483_A la_oenb_mprj[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input484_A la_oenb_mprj[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input485_A la_oenb_mprj[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input486_A la_oenb_mprj[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input487_A la_oenb_mprj[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input488_A la_oenb_mprj[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input489_A la_oenb_mprj[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input48_A la_data_out_core[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input490_A la_oenb_mprj[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input491_A la_oenb_mprj[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input492_A la_oenb_mprj[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input493_A la_oenb_mprj[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input494_A la_oenb_mprj[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input495_A la_oenb_mprj[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input496_A la_oenb_mprj[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input497_A la_oenb_mprj[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input498_A la_oenb_mprj[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input499_A la_oenb_mprj[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input49_A la_data_out_core[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input4_A la_data_out_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input500_A la_oenb_mprj[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input501_A la_oenb_mprj[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input502_A la_oenb_mprj[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input503_A la_oenb_mprj[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input504_A la_oenb_mprj[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input505_A la_oenb_mprj[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input506_A la_oenb_mprj[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input507_A la_oenb_mprj[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input508_A la_oenb_mprj[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input509_A la_oenb_mprj[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input50_A la_data_out_core[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input510_A la_oenb_mprj[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input511_A la_oenb_mprj[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input512_A la_oenb_mprj[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input513_A la_oenb_mprj[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input514_A la_oenb_mprj[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input515_A la_oenb_mprj[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input516_A mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input517_A mprj_adr_o_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input518_A mprj_adr_o_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input519_A mprj_adr_o_core[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input51_A la_data_out_core[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input520_A mprj_adr_o_core[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input521_A mprj_adr_o_core[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input522_A mprj_adr_o_core[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input523_A mprj_adr_o_core[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input524_A mprj_adr_o_core[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input525_A mprj_adr_o_core[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input526_A mprj_adr_o_core[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input527_A mprj_adr_o_core[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input528_A mprj_adr_o_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input529_A mprj_adr_o_core[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input52_A la_data_out_core[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input530_A mprj_adr_o_core[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input531_A mprj_adr_o_core[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input532_A mprj_adr_o_core[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input533_A mprj_adr_o_core[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input534_A mprj_adr_o_core[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input535_A mprj_adr_o_core[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input536_A mprj_adr_o_core[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input537_A mprj_adr_o_core[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input538_A mprj_adr_o_core[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input539_A mprj_adr_o_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input53_A la_data_out_core[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input540_A mprj_adr_o_core[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input541_A mprj_adr_o_core[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input542_A mprj_adr_o_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input543_A mprj_adr_o_core[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input544_A mprj_adr_o_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input545_A mprj_adr_o_core[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input546_A mprj_adr_o_core[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input547_A mprj_adr_o_core[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input548_A mprj_adr_o_core[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input549_A mprj_cyc_o_core vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input54_A la_data_out_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input550_A mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input551_A mprj_dat_i_user[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input552_A mprj_dat_i_user[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input553_A mprj_dat_i_user[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input554_A mprj_dat_i_user[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input555_A mprj_dat_i_user[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input556_A mprj_dat_i_user[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input557_A mprj_dat_i_user[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input558_A mprj_dat_i_user[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input559_A mprj_dat_i_user[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input55_A la_data_out_core[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input560_A mprj_dat_i_user[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input561_A mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input562_A mprj_dat_i_user[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input563_A mprj_dat_i_user[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input564_A mprj_dat_i_user[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input565_A mprj_dat_i_user[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input566_A mprj_dat_i_user[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input567_A mprj_dat_i_user[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input568_A mprj_dat_i_user[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input569_A mprj_dat_i_user[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input56_A la_data_out_core[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input570_A mprj_dat_i_user[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input571_A mprj_dat_i_user[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input572_A mprj_dat_i_user[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input573_A mprj_dat_i_user[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input574_A mprj_dat_i_user[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input575_A mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input576_A mprj_dat_i_user[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input577_A mprj_dat_i_user[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input578_A mprj_dat_i_user[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input579_A mprj_dat_i_user[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input57_A la_data_out_core[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input580_A mprj_dat_i_user[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input581_A mprj_dat_i_user[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input582_A mprj_dat_o_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input583_A mprj_dat_o_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input584_A mprj_dat_o_core[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input585_A mprj_dat_o_core[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input586_A mprj_dat_o_core[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input587_A mprj_dat_o_core[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input588_A mprj_dat_o_core[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input589_A mprj_dat_o_core[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input58_A la_data_out_core[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input590_A mprj_dat_o_core[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input591_A mprj_dat_o_core[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input592_A mprj_dat_o_core[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input593_A mprj_dat_o_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input594_A mprj_dat_o_core[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input595_A mprj_dat_o_core[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input596_A mprj_dat_o_core[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input597_A mprj_dat_o_core[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input598_A mprj_dat_o_core[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input599_A mprj_dat_o_core[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input59_A la_data_out_core[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input5_A la_data_out_core[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input600_A mprj_dat_o_core[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input601_A mprj_dat_o_core[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input602_A mprj_dat_o_core[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input603_A mprj_dat_o_core[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input604_A mprj_dat_o_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input605_A mprj_dat_o_core[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input606_A mprj_dat_o_core[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input607_A mprj_dat_o_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input608_A mprj_dat_o_core[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input609_A mprj_dat_o_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input60_A la_data_out_core[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input610_A mprj_dat_o_core[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input611_A mprj_dat_o_core[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input612_A mprj_dat_o_core[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input613_A mprj_dat_o_core[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input614_A mprj_iena_wb vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input615_A mprj_sel_o_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input616_A mprj_sel_o_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input617_A mprj_sel_o_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input618_A mprj_sel_o_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input619_A mprj_stb_o_core vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input61_A la_data_out_core[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input620_A mprj_we_o_core vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input621_A user_irq_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input622_A user_irq_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input623_A user_irq_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input624_A user_irq_ena[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input625_A user_irq_ena[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input626_A user_irq_ena[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input62_A la_data_out_core[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input63_A la_data_out_core[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input64_A la_data_out_core[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input65_A la_data_out_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input66_A la_data_out_core[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input67_A la_data_out_core[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input68_A la_data_out_core[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input69_A la_data_out_core[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input6_A la_data_out_core[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input70_A la_data_out_core[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input71_A la_data_out_core[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input72_A la_data_out_core[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input73_A la_data_out_core[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input74_A la_data_out_core[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input75_A la_data_out_core[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input76_A la_data_out_core[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input77_A la_data_out_core[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input78_A la_data_out_core[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input79_A la_data_out_core[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input7_A la_data_out_core[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input80_A la_data_out_core[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input81_A la_data_out_core[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input82_A la_data_out_core[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input83_A la_data_out_core[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input84_A la_data_out_core[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input85_A la_data_out_core[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input86_A la_data_out_core[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input87_A la_data_out_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input88_A la_data_out_core[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input89_A la_data_out_core[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input8_A la_data_out_core[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input90_A la_data_out_core[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input91_A la_data_out_core[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input92_A la_data_out_core[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input93_A la_data_out_core[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input94_A la_data_out_core[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input95_A la_data_out_core[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input96_A la_data_out_core[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input97_A la_data_out_core[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input98_A la_data_out_core[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input99_A la_data_out_core[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input9_A la_data_out_core[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[0]_A  _073_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[0]_TE  \la_data_out_enable[0]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[100]_A  _074_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[100]_TE  \la_data_out_enable[100]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[101]_A  _075_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[101]_TE  \la_data_out_enable[101]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[102]_A  _076_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[102]_TE  \la_data_out_enable[102]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[103]_A  _077_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[103]_TE  \la_data_out_enable[103]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[104]_A  _078_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[104]_TE  \la_data_out_enable[104]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[105]_A  _079_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[105]_TE  \la_data_out_enable[105]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[106]_A  _080_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[106]_TE  \la_data_out_enable[106]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[107]_A  _081_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[107]_TE  \la_data_out_enable[107]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[108]_A  _082_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[108]_TE  \la_data_out_enable[108]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[109]_A  _083_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[109]_TE  \la_data_out_enable[109]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[10]_A  _084_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[10]_TE  \la_data_out_enable[10]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[110]_A  _085_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[110]_TE  \la_data_out_enable[110]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[111]_A  _086_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[111]_TE  \la_data_out_enable[111]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[112]_A  _087_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[112]_TE  \la_data_out_enable[112]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[113]_A  _088_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[113]_TE  \la_data_out_enable[113]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[114]_A  _089_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[114]_TE  \la_data_out_enable[114]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[115]_A  _090_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[115]_TE  \la_data_out_enable[115]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[116]_A  _091_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[116]_TE  \la_data_out_enable[116]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[117]_A  _092_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[117]_TE  \la_data_out_enable[117]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[118]_A  _093_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[118]_TE  \la_data_out_enable[118]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[119]_A  _094_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[119]_TE  \la_data_out_enable[119]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[11]_A  _095_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[11]_TE  \la_data_out_enable[11]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[120]_A  _096_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[120]_TE  \la_data_out_enable[120]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[121]_A  _097_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[121]_TE  \la_data_out_enable[121]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[122]_A  _098_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[122]_TE  \la_data_out_enable[122]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[123]_A  _099_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[123]_TE  \la_data_out_enable[123]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[124]_A  _100_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[124]_TE  \la_data_out_enable[124]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[125]_A  _101_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[125]_TE  \la_data_out_enable[125]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[126]_A  _102_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[126]_TE  \la_data_out_enable[126]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[127]_A  _103_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[127]_TE  \la_data_out_enable[127]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[12]_A  _104_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[12]_TE  \la_data_out_enable[12]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[13]_A  _105_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[13]_TE  \la_data_out_enable[13]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[14]_A  _106_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[14]_TE  \la_data_out_enable[14]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[15]_A  _107_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[15]_TE  \la_data_out_enable[15]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[16]_A  _108_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[16]_TE  \la_data_out_enable[16]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[17]_A  _109_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[17]_TE  \la_data_out_enable[17]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[18]_A  _110_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[18]_TE  \la_data_out_enable[18]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[19]_A  _111_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[19]_TE  \la_data_out_enable[19]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[1]_A  _112_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[1]_TE  \la_data_out_enable[1]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[20]_A  _113_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[20]_TE  \la_data_out_enable[20]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[21]_A  _114_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[21]_TE  \la_data_out_enable[21]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[22]_A  _115_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[22]_TE  \la_data_out_enable[22]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[23]_A  _116_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[23]_TE  \la_data_out_enable[23]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[24]_A  _117_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[24]_TE  \la_data_out_enable[24]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[25]_A  _118_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[25]_TE  \la_data_out_enable[25]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[26]_A  _119_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[26]_TE  \la_data_out_enable[26]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[27]_A  _120_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[27]_TE  \la_data_out_enable[27]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[28]_A  _121_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[28]_TE  \la_data_out_enable[28]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[29]_A  _122_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[29]_TE  \la_data_out_enable[29]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[2]_A  _123_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[2]_TE  \la_data_out_enable[2]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[30]_A  _124_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[30]_TE  \la_data_out_enable[30]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[31]_A  _125_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[31]_TE  \la_data_out_enable[31]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[32]_A  _126_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[32]_TE  \la_data_out_enable[32]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[33]_A  _127_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[33]_TE  \la_data_out_enable[33]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[34]_A  _128_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[34]_TE  \la_data_out_enable[34]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[35]_A  _129_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[35]_TE  \la_data_out_enable[35]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[36]_A  _130_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[36]_TE  \la_data_out_enable[36]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[37]_A  _131_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[37]_TE  \la_data_out_enable[37]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[38]_A  _132_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[38]_TE  \la_data_out_enable[38]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[39]_A  _133_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[39]_TE  \la_data_out_enable[39]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[3]_A  _134_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[3]_TE  \la_data_out_enable[3]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[40]_A  _135_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[40]_TE  \la_data_out_enable[40]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[41]_A  _136_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[41]_TE  \la_data_out_enable[41]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[42]_A  _137_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[42]_TE  \la_data_out_enable[42]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[43]_A  _138_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[43]_TE  \la_data_out_enable[43]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[44]_A  _139_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[44]_TE  \la_data_out_enable[44]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[45]_A  _140_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[45]_TE  \la_data_out_enable[45]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[46]_A  _141_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[46]_TE  \la_data_out_enable[46]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[47]_A  _142_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[47]_TE  \la_data_out_enable[47]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[48]_A  _143_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[48]_TE  \la_data_out_enable[48]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[49]_A  _144_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[49]_TE  \la_data_out_enable[49]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[4]_A  _145_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[4]_TE  \la_data_out_enable[4]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[50]_A  _146_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[50]_TE  \la_data_out_enable[50]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[51]_A  _147_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[51]_TE  \la_data_out_enable[51]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[52]_A  _148_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[52]_TE  \la_data_out_enable[52]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[53]_A  _149_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[53]_TE  \la_data_out_enable[53]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[54]_A  _150_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[54]_TE  \la_data_out_enable[54]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[55]_A  _151_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[55]_TE  \la_data_out_enable[55]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[56]_A  _152_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[56]_TE  \la_data_out_enable[56]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[57]_A  _153_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[57]_TE  \la_data_out_enable[57]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[58]_A  _154_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[58]_TE  \la_data_out_enable[58]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[59]_A  _155_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[59]_TE  \la_data_out_enable[59]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[5]_A  _156_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[5]_TE  \la_data_out_enable[5]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[60]_A  _157_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[60]_TE  \la_data_out_enable[60]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[61]_A  _158_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[61]_TE  \la_data_out_enable[61]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[62]_A  _159_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[62]_TE  \la_data_out_enable[62]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[63]_A  _160_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[63]_TE  \la_data_out_enable[63]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[64]_A  _161_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[64]_TE  \la_data_out_enable[64]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[65]_A  _162_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[65]_TE  \la_data_out_enable[65]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[66]_A  _163_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[66]_TE  \la_data_out_enable[66]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[67]_A  _164_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[67]_TE  \la_data_out_enable[67]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[68]_A  _165_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[68]_TE  \la_data_out_enable[68]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[69]_A  _166_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[69]_TE  \la_data_out_enable[69]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[6]_A  _167_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[6]_TE  \la_data_out_enable[6]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[70]_A  _168_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[70]_TE  \la_data_out_enable[70]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[71]_A  _169_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[71]_TE  \la_data_out_enable[71]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[72]_A  _170_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[72]_TE  \la_data_out_enable[72]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[73]_A  _171_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[73]_TE  \la_data_out_enable[73]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[74]_A  _172_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[74]_TE  \la_data_out_enable[74]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[75]_A  _173_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[75]_TE  \la_data_out_enable[75]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[76]_A  _174_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[76]_TE  \la_data_out_enable[76]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[77]_A  _175_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[77]_TE  \la_data_out_enable[77]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[78]_A  _176_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[78]_TE  \la_data_out_enable[78]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[79]_A  _177_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[79]_TE  \la_data_out_enable[79]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[7]_A  _178_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[7]_TE  \la_data_out_enable[7]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[80]_A  _179_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[80]_TE  \la_data_out_enable[80]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[81]_A  _180_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[81]_TE  \la_data_out_enable[81]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[82]_A  _181_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[82]_TE  \la_data_out_enable[82]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[83]_A  _182_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[83]_TE  \la_data_out_enable[83]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[84]_A  _183_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[84]_TE  \la_data_out_enable[84]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[85]_A  _184_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[85]_TE  \la_data_out_enable[85]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[86]_A  _185_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[86]_TE  \la_data_out_enable[86]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[87]_A  _186_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[87]_TE  \la_data_out_enable[87]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[88]_A  _187_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[88]_TE  \la_data_out_enable[88]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[89]_A  _188_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[89]_TE  \la_data_out_enable[89]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[8]_A  _189_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[8]_TE  \la_data_out_enable[8]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[90]_A  _190_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[90]_TE  \la_data_out_enable[90]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[91]_A  _191_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[91]_TE  \la_data_out_enable[91]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[92]_A  _192_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[92]_TE  \la_data_out_enable[92]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[93]_A  _193_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[93]_TE  \la_data_out_enable[93]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[94]_A  _194_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[94]_TE  \la_data_out_enable[94]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[95]_A  _195_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[95]_TE  \la_data_out_enable[95]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[96]_A  _196_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[96]_TE  \la_data_out_enable[96]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[97]_A  _197_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[97]_TE  \la_data_out_enable[97]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[98]_A  _198_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[98]_TE  \la_data_out_enable[98]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[99]_A  _199_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[99]_TE  \la_data_out_enable[99]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[9]_A  _200_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf[9]_TE  \la_data_out_enable[9]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[0]_A_N  net388 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[0]_B  \mprj_logic1[74]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[100]_A_N  net389 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[100]_B  \mprj_logic1[174]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[101]_A_N  net390 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[101]_B  \mprj_logic1[175]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[102]_A_N  net391 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[102]_B  \mprj_logic1[176]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[103]_A_N  net392 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[103]_B  \mprj_logic1[177]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[104]_A_N  net393 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[104]_B  \mprj_logic1[178]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[105]_A_N  net394 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[105]_B  \mprj_logic1[179]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[106]_A_N  net395 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[106]_B  \mprj_logic1[180]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[107]_A_N  net396 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[107]_B  \mprj_logic1[181]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[108]_A_N  net397 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[108]_B  \mprj_logic1[182]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[109]_A_N  net398 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[109]_B  \mprj_logic1[183]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[10]_A_N  net399 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[10]_B  \mprj_logic1[84]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[110]_A_N  net400 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[110]_B  \mprj_logic1[184]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[111]_A_N  net401 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[111]_B  \mprj_logic1[185]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[112]_A_N  net402 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[112]_B  \mprj_logic1[186]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[113]_A_N  net403 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[113]_B  \mprj_logic1[187]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[114]_A_N  net404 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[114]_B  \mprj_logic1[188]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[115]_A_N  net405 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[115]_B  \mprj_logic1[189]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[116]_A_N  net406 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[116]_B  \mprj_logic1[190]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[117]_A_N  net407 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[117]_B  \mprj_logic1[191]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[118]_A_N  net408 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[118]_B  \mprj_logic1[192]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[119]_A_N  net409 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[119]_B  \mprj_logic1[193]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[11]_A_N  net410 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[11]_B  \mprj_logic1[85]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[120]_A_N  net411 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[120]_B  \mprj_logic1[194]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[121]_A_N  net412 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[121]_B  \mprj_logic1[195]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[122]_A_N  net413 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[122]_B  \mprj_logic1[196]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[123]_A_N  net414 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[123]_B  \mprj_logic1[197]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[124]_A_N  net415 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[124]_B  \mprj_logic1[198]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[125]_A_N  net416 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[125]_B  \mprj_logic1[199]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[126]_A_N  net417 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[126]_B  \mprj_logic1[200]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[127]_A_N  net418 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[127]_B  \mprj_logic1[201]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[12]_A_N  net419 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[12]_B  \mprj_logic1[86]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[13]_A_N  net420 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[13]_B  \mprj_logic1[87]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[14]_A_N  net421 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[14]_B  \mprj_logic1[88]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[15]_A_N  net422 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[15]_B  \mprj_logic1[89]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[16]_A_N  net423 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[16]_B  \mprj_logic1[90]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[17]_A_N  net424 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[17]_B  \mprj_logic1[91]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[18]_A_N  net425 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[18]_B  \mprj_logic1[92]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[19]_A_N  net426 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[19]_B  \mprj_logic1[93]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[1]_A_N  net427 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[1]_B  \mprj_logic1[75]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[20]_A_N  net428 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[20]_B  \mprj_logic1[94]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[21]_A_N  net429 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[21]_B  \mprj_logic1[95]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[22]_A_N  net430 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[22]_B  \mprj_logic1[96]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[23]_A_N  net431 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[23]_B  \mprj_logic1[97]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[24]_A_N  net432 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[24]_B  \mprj_logic1[98]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[25]_A_N  net433 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[25]_B  \mprj_logic1[99]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[26]_A_N  net434 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[26]_B  \mprj_logic1[100]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[27]_A_N  net435 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[27]_B  \mprj_logic1[101]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[28]_A_N  net436 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[28]_B  \mprj_logic1[102]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[29]_A_N  net437 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[29]_B  \mprj_logic1[103]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[2]_A_N  net438 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[2]_B  \mprj_logic1[76]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[30]_A_N  net439 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[30]_B  \mprj_logic1[104]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[31]_A_N  net440 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[31]_B  \mprj_logic1[105]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[32]_A_N  net441 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[32]_B  \mprj_logic1[106]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[33]_A_N  net442 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[33]_B  \mprj_logic1[107]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[34]_A_N  net443 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[34]_B  \mprj_logic1[108]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[35]_A_N  net444 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[35]_B  \mprj_logic1[109]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[36]_A_N  net445 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[36]_B  \mprj_logic1[110]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[37]_A_N  net446 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[37]_B  \mprj_logic1[111]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[38]_A_N  net447 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[38]_B  \mprj_logic1[112]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[39]_A_N  net448 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[39]_B  \mprj_logic1[113]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[3]_A_N  net449 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[3]_B  \mprj_logic1[77]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[40]_A_N  net450 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[40]_B  \mprj_logic1[114]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[41]_A_N  net451 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[41]_B  \mprj_logic1[115]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[42]_A_N  net452 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[42]_B  \mprj_logic1[116]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[43]_A_N  net453 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[43]_B  \mprj_logic1[117]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[44]_A_N  net454 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[44]_B  \mprj_logic1[118]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[45]_A_N  net455 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[45]_B  \mprj_logic1[119]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[46]_A_N  net456 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[46]_B  \mprj_logic1[120]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[47]_A_N  net457 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[47]_B  \mprj_logic1[121]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[48]_A_N  net458 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[48]_B  \mprj_logic1[122]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[49]_A_N  net459 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[49]_B  \mprj_logic1[123]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[4]_A_N  net460 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[4]_B  \mprj_logic1[78]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[50]_A_N  net461 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[50]_B  \mprj_logic1[124]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[51]_A_N  net462 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[51]_B  \mprj_logic1[125]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[52]_A_N  net463 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[52]_B  \mprj_logic1[126]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[53]_A_N  net464 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[53]_B  \mprj_logic1[127]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[54]_A_N  net465 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[54]_B  \mprj_logic1[128]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[55]_A_N  net466 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[55]_B  \mprj_logic1[129]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[56]_A_N  net467 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[56]_B  \mprj_logic1[130]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[57]_A_N  net468 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[57]_B  \mprj_logic1[131]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[58]_A_N  net469 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[58]_B  \mprj_logic1[132]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[59]_A_N  net470 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[59]_B  \mprj_logic1[133]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[5]_A_N  net471 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[5]_B  \mprj_logic1[79]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[60]_A_N  net472 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[60]_B  \mprj_logic1[134]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[61]_A_N  net473 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[61]_B  \mprj_logic1[135]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[62]_A_N  net474 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[62]_B  \mprj_logic1[136]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[63]_A_N  net475 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[63]_B  \mprj_logic1[137]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[64]_A_N  net476 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[64]_B  \mprj_logic1[138]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[65]_A_N  net477 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[65]_B  \mprj_logic1[139]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[66]_A_N  net478 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[66]_B  \mprj_logic1[140]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[67]_A_N  net479 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[67]_B  \mprj_logic1[141]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[68]_A_N  net480 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[68]_B  \mprj_logic1[142]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[69]_A_N  net481 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[69]_B  \mprj_logic1[143]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[6]_A_N  net482 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[6]_B  \mprj_logic1[80]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[70]_A_N  net483 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[70]_B  \mprj_logic1[144]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[71]_A_N  net484 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[71]_B  \mprj_logic1[145]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[72]_A_N  net485 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[72]_B  \mprj_logic1[146]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[73]_A_N  net486 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[73]_B  \mprj_logic1[147]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[74]_A_N  net487 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[74]_B  \mprj_logic1[148]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[75]_A_N  net488 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[75]_B  \mprj_logic1[149]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[76]_A_N  net489 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[76]_B  \mprj_logic1[150]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[77]_A_N  net490 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[77]_B  \mprj_logic1[151]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[78]_A_N  net491 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[78]_B  \mprj_logic1[152]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[79]_A_N  net492 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[79]_B  \mprj_logic1[153]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[7]_A_N  net493 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[7]_B  \mprj_logic1[81]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[80]_A_N  net494 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[80]_B  \mprj_logic1[154]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[81]_A_N  net495 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[81]_B  \mprj_logic1[155]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[82]_A_N  net496 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[82]_B  \mprj_logic1[156]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[83]_A_N  net497 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[83]_B  \mprj_logic1[157]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[84]_A_N  net498 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[84]_B  \mprj_logic1[158]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[85]_A_N  net499 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[85]_B  \mprj_logic1[159]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[86]_A_N  net500 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[86]_B  \mprj_logic1[160]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[87]_A_N  net501 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[87]_B  \mprj_logic1[161]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[88]_A_N  net502 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[88]_B  \mprj_logic1[162]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[89]_A_N  net503 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[89]_B  \mprj_logic1[163]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[8]_A_N  net504 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[8]_B  \mprj_logic1[82]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[90]_A_N  net505 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[90]_B  \mprj_logic1[164]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[91]_A_N  net506 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[91]_B  \mprj_logic1[165]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[92]_A_N  net507 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[92]_B  \mprj_logic1[166]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[93]_A_N  net508 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[93]_B  \mprj_logic1[167]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[94]_A_N  net509 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[94]_B  \mprj_logic1[168]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[95]_A_N  net510 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[95]_B  \mprj_logic1[169]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[96]_A_N  net511 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[96]_B  \mprj_logic1[170]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[97]_A_N  net512 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[97]_B  \mprj_logic1[171]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[98]_A_N  net513 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[98]_B  \mprj_logic1[172]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[99]_A_N  net514 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[99]_B  \mprj_logic1[173]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[9]_A_N  net515 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_la_buf_enable[9]_B  \mprj_logic1[83]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj2_pwrgood_A mprj2_logic1 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj2_vdd_pwrgood_A mprj2_vdd_logic1 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[0]_A  _009_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[0]_TE  \mprj_logic1[10]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[10]_A  _010_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[10]_TE  \mprj_logic1[20]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[11]_A  _011_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[11]_TE  \mprj_logic1[21]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[12]_A  _012_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[12]_TE  \mprj_logic1[22]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[13]_A  _013_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[13]_TE  \mprj_logic1[23]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[14]_A  _014_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[14]_TE  \mprj_logic1[24]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[15]_A  _015_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[15]_TE  \mprj_logic1[25]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[16]_A  _016_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[16]_TE  \mprj_logic1[26]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[17]_A  _017_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[17]_TE  \mprj_logic1[27]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[18]_A  _018_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[18]_TE  \mprj_logic1[28]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[19]_A  _019_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[19]_TE  \mprj_logic1[29]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[1]_A  _020_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[1]_TE  \mprj_logic1[11]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[20]_A  _021_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[20]_TE  \mprj_logic1[30]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[21]_A  _022_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[21]_TE  \mprj_logic1[31]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[22]_A  _023_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[22]_TE  \mprj_logic1[32]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[23]_A  _024_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[23]_TE  \mprj_logic1[33]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[24]_A  _025_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[24]_TE  \mprj_logic1[34]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[25]_A  _026_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[25]_TE  \mprj_logic1[35]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[26]_A  _027_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[26]_TE  \mprj_logic1[36]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[27]_A  _028_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[27]_TE  \mprj_logic1[37]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[28]_A  _029_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[28]_TE  \mprj_logic1[38]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[29]_A  _030_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[29]_TE  \mprj_logic1[39]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[2]_A  _031_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[2]_TE  \mprj_logic1[12]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[30]_A  _032_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[30]_TE  \mprj_logic1[40]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[31]_A  _033_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[31]_TE  \mprj_logic1[41]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[3]_A  _034_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[3]_TE  \mprj_logic1[13]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[4]_A  _035_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[4]_TE  \mprj_logic1[14]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[5]_A  _036_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[5]_TE  \mprj_logic1[15]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[6]_A  _037_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[6]_TE  \mprj_logic1[16]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[7]_A  _038_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[7]_TE  \mprj_logic1[17]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[8]_A  _039_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[8]_TE  \mprj_logic1[18]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[9]_A  _040_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_adr_buf[9]_TE  \mprj_logic1[19]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_clk2_buf_A _001_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_clk2_buf_TE \mprj_logic1[2]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_clk_buf_A _000_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_clk_buf_TE \mprj_logic1[1]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_cyc_buf_A _002_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_cyc_buf_TE \mprj_logic1[3]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[0]_A  _041_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[0]_TE  \mprj_logic1[42]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[10]_A  _042_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[10]_TE  \mprj_logic1[52]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[11]_A  _043_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[11]_TE  \mprj_logic1[53]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[12]_A  _044_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[12]_TE  \mprj_logic1[54]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[13]_A  _045_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[13]_TE  \mprj_logic1[55]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[14]_A  _046_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[14]_TE  \mprj_logic1[56]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[15]_A  _047_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[15]_TE  \mprj_logic1[57]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[16]_A  _048_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[16]_TE  \mprj_logic1[58]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[17]_A  _049_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[17]_TE  \mprj_logic1[59]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[18]_A  _050_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[18]_TE  \mprj_logic1[60]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[19]_A  _051_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[19]_TE  \mprj_logic1[61]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[1]_A  _052_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[1]_TE  \mprj_logic1[43]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[20]_A  _053_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[20]_TE  \mprj_logic1[62]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[21]_A  _054_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[21]_TE  \mprj_logic1[63]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[22]_A  _055_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[22]_TE  \mprj_logic1[64]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[23]_A  _056_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[23]_TE  \mprj_logic1[65]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[24]_A  _057_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[24]_TE  \mprj_logic1[66]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[25]_A  _058_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[25]_TE  \mprj_logic1[67]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[26]_A  _059_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[26]_TE  \mprj_logic1[68]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[27]_A  _060_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[27]_TE  \mprj_logic1[69]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[28]_A  _061_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[28]_TE  \mprj_logic1[70]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[29]_A  _062_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[29]_TE  \mprj_logic1[71]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[2]_A  _063_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[2]_TE  \mprj_logic1[44]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[30]_A  _064_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[30]_TE  \mprj_logic1[72]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[31]_A  _065_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[31]_TE  \mprj_logic1[73]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[3]_A  _066_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[3]_TE  \mprj_logic1[45]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[4]_A  _067_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[4]_TE  \mprj_logic1[46]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[5]_A  _068_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[5]_TE  \mprj_logic1[47]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[6]_A  _069_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[6]_TE  \mprj_logic1[48]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[7]_A  _070_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[7]_TE  \mprj_logic1[49]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[8]_A  _071_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[8]_TE  \mprj_logic1[50]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[9]_A  _072_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_dat_buf[9]_TE  \mprj_logic1[51]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_pwrgood_A \mprj_logic1[461]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_rstn_buf_A net3 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_rstn_buf_TE \mprj_logic1[0]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_sel_buf[0]_A  _005_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_sel_buf[0]_TE  \mprj_logic1[6]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_sel_buf[1]_A  _006_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_sel_buf[1]_TE  \mprj_logic1[7]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_sel_buf[2]_A  _007_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_sel_buf[2]_TE  \mprj_logic1[8]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_sel_buf[3]_A  _008_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_mprj_sel_buf[3]_TE  \mprj_logic1[9]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_stb_buf_A _003_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_stb_buf_TE \mprj_logic1[4]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_vdd_pwrgood_A mprj_vdd_logic1 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_we_buf_A _004_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_we_buf_TE \mprj_logic1[5]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output627_A net627 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output628_A net628 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output629_A net629 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output630_A net630 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output631_A net631 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output632_A net632 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output633_A net633 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output634_A net634 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output635_A net635 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output636_A net636 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output637_A net637 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output638_A net638 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output639_A net639 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output640_A net640 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output641_A net641 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output642_A net642 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output643_A net643 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output644_A net644 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output645_A net645 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output646_A net646 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output647_A net647 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output648_A net648 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output649_A net649 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output650_A net650 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output651_A net651 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output652_A net652 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output653_A net653 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output654_A net654 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output655_A net655 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output656_A net656 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output657_A net657 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output658_A net658 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output659_A net659 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output660_A net660 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output661_A net661 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output662_A net662 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output663_A net663 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output664_A net664 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output665_A net665 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output666_A net666 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output667_A net667 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output668_A net668 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output669_A net669 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output670_A net670 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output671_A net671 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output672_A net672 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output673_A net673 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output674_A net674 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output675_A net675 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output676_A net676 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output677_A net677 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output678_A net678 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output679_A net679 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output680_A net680 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output681_A net681 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output682_A net682 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output683_A net683 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output684_A net684 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output685_A net685 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output686_A net686 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output687_A net687 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output688_A net688 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output689_A net689 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output690_A net690 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output691_A net691 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output692_A net692 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output693_A net693 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output694_A net694 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output695_A net695 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output696_A net696 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output697_A net697 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output698_A net698 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output699_A net699 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output700_A net700 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output701_A net701 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output702_A net702 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output703_A net703 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output704_A net704 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output705_A net705 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output706_A net706 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output707_A net707 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output708_A net708 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output709_A net709 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output710_A net710 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output711_A net711 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output712_A net712 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output713_A net713 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output714_A net714 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output715_A net715 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output716_A net716 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output717_A net717 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output718_A net718 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output719_A net719 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output720_A net720 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output721_A net721 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output722_A net722 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output723_A net723 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output724_A net724 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output725_A net725 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output726_A net726 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output727_A net727 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output728_A net728 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output729_A net729 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output730_A net730 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output731_A net731 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output732_A net732 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output733_A net733 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output734_A net734 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output735_A net735 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output736_A net736 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output737_A net737 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output738_A net738 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output739_A net739 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output740_A net740 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output741_A net741 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output742_A net742 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output743_A net743 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output744_A net744 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output745_A net745 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output746_A net746 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output747_A net747 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output748_A net748 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output749_A net749 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output750_A net750 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output751_A net751 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output752_A net752 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output753_A net753 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output754_A net754 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output755_A net755 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output756_A net756 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output757_A net757 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output758_A net758 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output759_A net759 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output760_A net760 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output761_A net761 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output762_A net762 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output763_A net763 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output764_A net764 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output765_A net765 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output766_A net766 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output767_A net767 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output768_A net768 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output769_A net769 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output770_A net770 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output771_A net771 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output772_A net772 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output773_A net773 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output774_A net774 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output775_A net775 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output776_A net776 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output777_A net777 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output778_A net778 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output779_A net779 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output780_A net780 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output781_A net781 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output782_A net782 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output783_A net783 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output784_A net784 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output785_A net785 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output786_A net786 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output787_A net787 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output788_A net788 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output789_A net789 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output790_A net790 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output791_A net791 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output792_A net792 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output793_A net793 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output794_A net794 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_irq_buffers[0]_A  \user_irq_bar[0]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_irq_buffers[1]_A  \user_irq_bar[1]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_irq_buffers[2]_A  \user_irq_bar[2]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_irq_ena_buf[0]_A  net624 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_irq_ena_buf[0]_B  \mprj_logic1[458]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_irq_ena_buf[1]_A  net625 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_irq_ena_buf[1]_B  \mprj_logic1[459]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_irq_ena_buf[2]_A  net626 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_irq_ena_buf[2]_B  \mprj_logic1[460]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_irq_gates[0]_A  net621 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_irq_gates[0]_B  \user_irq_enable[0]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_irq_gates[1]_A  net622 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_irq_gates[1]_B  \user_irq_enable[1]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_irq_gates[2]_A  net623 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_irq_gates[2]_B  \user_irq_enable[2]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[0]_A  \la_data_in_mprj_bar[0]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[100]_A  \la_data_in_mprj_bar[100]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[101]_A  \la_data_in_mprj_bar[101]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[102]_A  \la_data_in_mprj_bar[102]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[103]_A  \la_data_in_mprj_bar[103]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[104]_A  \la_data_in_mprj_bar[104]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[105]_A  \la_data_in_mprj_bar[105]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[106]_A  \la_data_in_mprj_bar[106]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[107]_A  \la_data_in_mprj_bar[107]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[108]_A  \la_data_in_mprj_bar[108]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[109]_A  \la_data_in_mprj_bar[109]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[10]_A  \la_data_in_mprj_bar[10]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[110]_A  \la_data_in_mprj_bar[110]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[111]_A  \la_data_in_mprj_bar[111]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[112]_A  \la_data_in_mprj_bar[112]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[113]_A  \la_data_in_mprj_bar[113]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[114]_A  \la_data_in_mprj_bar[114]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[115]_A  \la_data_in_mprj_bar[115]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[116]_A  \la_data_in_mprj_bar[116]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[117]_A  \la_data_in_mprj_bar[117]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[118]_A  \la_data_in_mprj_bar[118]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[119]_A  \la_data_in_mprj_bar[119]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[11]_A  \la_data_in_mprj_bar[11]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[120]_A  \la_data_in_mprj_bar[120]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[121]_A  \la_data_in_mprj_bar[121]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[122]_A  \la_data_in_mprj_bar[122]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[123]_A  \la_data_in_mprj_bar[123]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[124]_A  \la_data_in_mprj_bar[124]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[125]_A  \la_data_in_mprj_bar[125]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[126]_A  \la_data_in_mprj_bar[126]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[127]_A  \la_data_in_mprj_bar[127]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[12]_A  \la_data_in_mprj_bar[12]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[13]_A  \la_data_in_mprj_bar[13]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[14]_A  \la_data_in_mprj_bar[14]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[15]_A  \la_data_in_mprj_bar[15]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[16]_A  \la_data_in_mprj_bar[16]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[17]_A  \la_data_in_mprj_bar[17]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[18]_A  \la_data_in_mprj_bar[18]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[19]_A  \la_data_in_mprj_bar[19]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[1]_A  \la_data_in_mprj_bar[1]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[20]_A  \la_data_in_mprj_bar[20]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[21]_A  \la_data_in_mprj_bar[21]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[22]_A  \la_data_in_mprj_bar[22]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[23]_A  \la_data_in_mprj_bar[23]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[24]_A  \la_data_in_mprj_bar[24]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[25]_A  \la_data_in_mprj_bar[25]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[26]_A  \la_data_in_mprj_bar[26]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[27]_A  \la_data_in_mprj_bar[27]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[28]_A  \la_data_in_mprj_bar[28]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[29]_A  \la_data_in_mprj_bar[29]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[2]_A  \la_data_in_mprj_bar[2]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[30]_A  \la_data_in_mprj_bar[30]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[31]_A  \la_data_in_mprj_bar[31]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[32]_A  \la_data_in_mprj_bar[32]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[33]_A  \la_data_in_mprj_bar[33]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[34]_A  \la_data_in_mprj_bar[34]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[35]_A  \la_data_in_mprj_bar[35]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[36]_A  \la_data_in_mprj_bar[36]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[37]_A  \la_data_in_mprj_bar[37]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[38]_A  \la_data_in_mprj_bar[38]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[39]_A  \la_data_in_mprj_bar[39]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[3]_A  \la_data_in_mprj_bar[3]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[40]_A  \la_data_in_mprj_bar[40]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[41]_A  \la_data_in_mprj_bar[41]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[42]_A  \la_data_in_mprj_bar[42]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[43]_A  \la_data_in_mprj_bar[43]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[44]_A  \la_data_in_mprj_bar[44]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[45]_A  \la_data_in_mprj_bar[45]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[46]_A  \la_data_in_mprj_bar[46]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[47]_A  \la_data_in_mprj_bar[47]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[48]_A  \la_data_in_mprj_bar[48]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[49]_A  \la_data_in_mprj_bar[49]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[4]_A  \la_data_in_mprj_bar[4]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[50]_A  \la_data_in_mprj_bar[50]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[51]_A  \la_data_in_mprj_bar[51]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[52]_A  \la_data_in_mprj_bar[52]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[53]_A  \la_data_in_mprj_bar[53]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[54]_A  \la_data_in_mprj_bar[54]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[55]_A  \la_data_in_mprj_bar[55]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[56]_A  \la_data_in_mprj_bar[56]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[57]_A  \la_data_in_mprj_bar[57]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[58]_A  \la_data_in_mprj_bar[58]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[59]_A  \la_data_in_mprj_bar[59]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[5]_A  \la_data_in_mprj_bar[5]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[60]_A  \la_data_in_mprj_bar[60]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[61]_A  \la_data_in_mprj_bar[61]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[62]_A  \la_data_in_mprj_bar[62]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[63]_A  \la_data_in_mprj_bar[63]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[64]_A  \la_data_in_mprj_bar[64]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[65]_A  \la_data_in_mprj_bar[65]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[66]_A  \la_data_in_mprj_bar[66]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[67]_A  \la_data_in_mprj_bar[67]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[68]_A  \la_data_in_mprj_bar[68]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[69]_A  \la_data_in_mprj_bar[69]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[6]_A  \la_data_in_mprj_bar[6]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[70]_A  \la_data_in_mprj_bar[70]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[71]_A  \la_data_in_mprj_bar[71]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[72]_A  \la_data_in_mprj_bar[72]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[73]_A  \la_data_in_mprj_bar[73]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[74]_A  \la_data_in_mprj_bar[74]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[75]_A  \la_data_in_mprj_bar[75]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[76]_A  \la_data_in_mprj_bar[76]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[77]_A  \la_data_in_mprj_bar[77]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[78]_A  \la_data_in_mprj_bar[78]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[79]_A  \la_data_in_mprj_bar[79]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[7]_A  \la_data_in_mprj_bar[7]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[80]_A  \la_data_in_mprj_bar[80]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[81]_A  \la_data_in_mprj_bar[81]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[82]_A  \la_data_in_mprj_bar[82]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[83]_A  \la_data_in_mprj_bar[83]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[84]_A  \la_data_in_mprj_bar[84]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[85]_A  \la_data_in_mprj_bar[85]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[86]_A  \la_data_in_mprj_bar[86]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[87]_A  \la_data_in_mprj_bar[87]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[88]_A  \la_data_in_mprj_bar[88]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[89]_A  \la_data_in_mprj_bar[89]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[8]_A  \la_data_in_mprj_bar[8]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[90]_A  \la_data_in_mprj_bar[90]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[91]_A  \la_data_in_mprj_bar[91]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[92]_A  \la_data_in_mprj_bar[92]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[93]_A  \la_data_in_mprj_bar[93]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[94]_A  \la_data_in_mprj_bar[94]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[95]_A  \la_data_in_mprj_bar[95]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[96]_A  \la_data_in_mprj_bar[96]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[97]_A  \la_data_in_mprj_bar[97]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[98]_A  \la_data_in_mprj_bar[98]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[99]_A  \la_data_in_mprj_bar[99]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_buffers[9]_A  \la_data_in_mprj_bar[9]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[0]_A  net260 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[0]_B  \mprj_logic1[330]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[100]_A  net261 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[100]_B  \mprj_logic1[430]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[101]_A  net262 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[101]_B  \mprj_logic1[431]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[102]_A  net263 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[102]_B  \mprj_logic1[432]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[103]_A  net264 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[103]_B  \mprj_logic1[433]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[104]_A  net265 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[104]_B  \mprj_logic1[434]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[105]_A  net266 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[105]_B  \mprj_logic1[435]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[106]_A  net267 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[106]_B  \mprj_logic1[436]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[107]_A  net268 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[107]_B  \mprj_logic1[437]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[108]_A  net269 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[108]_B  \mprj_logic1[438]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[109]_A  net270 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[109]_B  \mprj_logic1[439]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[10]_A  net271 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[10]_B  \mprj_logic1[340]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[110]_A  net272 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[110]_B  \mprj_logic1[440]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[111]_A  net273 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[111]_B  \mprj_logic1[441]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[112]_A  net274 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[112]_B  \mprj_logic1[442]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[113]_A  net275 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[113]_B  \mprj_logic1[443]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[114]_A  net276 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[114]_B  \mprj_logic1[444]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[115]_A  net277 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[115]_B  \mprj_logic1[445]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[116]_A  net278 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[116]_B  \mprj_logic1[446]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[117]_A  net279 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[117]_B  \mprj_logic1[447]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[118]_A  net280 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[118]_B  \mprj_logic1[448]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[119]_A  net281 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[119]_B  \mprj_logic1[449]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[11]_A  net282 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[11]_B  \mprj_logic1[341]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[120]_A  net283 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[120]_B  \mprj_logic1[450]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[121]_A  net284 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[121]_B  \mprj_logic1[451]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[122]_A  net285 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[122]_B  \mprj_logic1[452]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[123]_A  net286 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[123]_B  \mprj_logic1[453]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[124]_A  net287 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[124]_B  \mprj_logic1[454]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[125]_A  net288 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[125]_B  \mprj_logic1[455]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[126]_A  net289 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[126]_B  \mprj_logic1[456]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[127]_A  net290 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[127]_B  \mprj_logic1[457]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[12]_A  net291 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[12]_B  \mprj_logic1[342]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[13]_A  net292 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[13]_B  \mprj_logic1[343]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[14]_A  net293 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[14]_B  \mprj_logic1[344]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[15]_A  net294 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[15]_B  \mprj_logic1[345]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[16]_A  net295 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[16]_B  \mprj_logic1[346]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[17]_A  net296 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[17]_B  \mprj_logic1[347]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[18]_A  net297 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[18]_B  \mprj_logic1[348]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[19]_A  net298 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[19]_B  \mprj_logic1[349]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[1]_A  net299 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[1]_B  \mprj_logic1[331]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[20]_A  net300 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[20]_B  \mprj_logic1[350]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[21]_A  net301 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[21]_B  \mprj_logic1[351]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[22]_A  net302 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[22]_B  \mprj_logic1[352]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[23]_A  net303 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[23]_B  \mprj_logic1[353]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[24]_A  net304 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[24]_B  \mprj_logic1[354]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[25]_A  net305 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[25]_B  \mprj_logic1[355]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[26]_A  net306 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[26]_B  \mprj_logic1[356]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[27]_A  net307 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[27]_B  \mprj_logic1[357]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[28]_A  net308 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[28]_B  \mprj_logic1[358]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[29]_A  net309 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[29]_B  \mprj_logic1[359]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[2]_A  net310 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[2]_B  \mprj_logic1[332]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[30]_A  net311 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[30]_B  \mprj_logic1[360]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[31]_A  net312 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[31]_B  \mprj_logic1[361]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[32]_A  net313 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[32]_B  \mprj_logic1[362]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[33]_A  net314 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[33]_B  \mprj_logic1[363]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[34]_A  net315 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[34]_B  \mprj_logic1[364]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[35]_A  net316 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[35]_B  \mprj_logic1[365]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[36]_A  net317 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[36]_B  \mprj_logic1[366]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[37]_A  net318 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[37]_B  \mprj_logic1[367]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[38]_A  net319 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[38]_B  \mprj_logic1[368]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[39]_A  net320 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[39]_B  \mprj_logic1[369]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[3]_A  net321 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[3]_B  \mprj_logic1[333]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[40]_A  net322 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[40]_B  \mprj_logic1[370]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[41]_A  net323 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[41]_B  \mprj_logic1[371]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[42]_A  net324 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[42]_B  \mprj_logic1[372]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[43]_A  net325 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[43]_B  \mprj_logic1[373]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[44]_A  net326 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[44]_B  \mprj_logic1[374]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[45]_A  net327 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[45]_B  \mprj_logic1[375]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[46]_A  net328 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[46]_B  \mprj_logic1[376]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[47]_A  net329 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[47]_B  \mprj_logic1[377]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[48]_A  net330 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[48]_B  \mprj_logic1[378]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[49]_A  net331 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[49]_B  \mprj_logic1[379]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[4]_A  net332 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[4]_B  \mprj_logic1[334]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[50]_A  net333 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[50]_B  \mprj_logic1[380]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[51]_A  net334 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[51]_B  \mprj_logic1[381]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[52]_A  net335 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[52]_B  \mprj_logic1[382]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[53]_A  net336 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[53]_B  \mprj_logic1[383]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[54]_A  net337 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[54]_B  \mprj_logic1[384]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[55]_A  net338 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[55]_B  \mprj_logic1[385]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[56]_A  net339 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[56]_B  \mprj_logic1[386]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[57]_A  net340 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[57]_B  \mprj_logic1[387]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[58]_A  net341 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[58]_B  \mprj_logic1[388]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[59]_A  net342 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[59]_B  \mprj_logic1[389]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[5]_A  net343 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[5]_B  \mprj_logic1[335]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[60]_A  net344 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[60]_B  \mprj_logic1[390]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[61]_A  net345 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[61]_B  \mprj_logic1[391]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[62]_A  net346 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[62]_B  \mprj_logic1[392]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[63]_A  net347 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[63]_B  \mprj_logic1[393]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[64]_A  net348 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[64]_B  \mprj_logic1[394]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[65]_A  net349 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[65]_B  \mprj_logic1[395]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[66]_A  net350 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[66]_B  \mprj_logic1[396]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[67]_A  net351 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[67]_B  \mprj_logic1[397]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[68]_A  net352 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[68]_B  \mprj_logic1[398]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[69]_A  net353 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[69]_B  \mprj_logic1[399]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[6]_A  net354 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[6]_B  \mprj_logic1[336]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[70]_A  net355 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[70]_B  \mprj_logic1[400]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[71]_A  net356 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[71]_B  \mprj_logic1[401]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[72]_A  net357 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[72]_B  \mprj_logic1[402]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[73]_A  net358 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[73]_B  \mprj_logic1[403]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[74]_A  net359 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[74]_B  \mprj_logic1[404]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[75]_A  net360 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[75]_B  \mprj_logic1[405]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[76]_A  net361 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[76]_B  \mprj_logic1[406]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[77]_A  net362 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[77]_B  \mprj_logic1[407]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[78]_A  net363 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[78]_B  \mprj_logic1[408]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[79]_A  net364 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[79]_B  \mprj_logic1[409]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[7]_A  net365 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[7]_B  \mprj_logic1[337]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[80]_A  net366 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[80]_B  \mprj_logic1[410]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[81]_A  net367 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[81]_B  \mprj_logic1[411]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[82]_A  net368 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[82]_B  \mprj_logic1[412]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[83]_A  net369 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[83]_B  \mprj_logic1[413]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[84]_A  net370 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[84]_B  \mprj_logic1[414]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[85]_A  net371 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[85]_B  \mprj_logic1[415]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[86]_A  net372 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[86]_B  \mprj_logic1[416]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[87]_A  net373 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[87]_B  \mprj_logic1[417]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[88]_A  net374 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[88]_B  \mprj_logic1[418]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[89]_A  net375 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[89]_B  \mprj_logic1[419]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[8]_A  net376 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[8]_B  \mprj_logic1[338]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[90]_A  net377 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[90]_B  \mprj_logic1[420]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[91]_A  net378 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[91]_B  \mprj_logic1[421]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[92]_A  net379 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[92]_B  \mprj_logic1[422]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[93]_A  net380 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[93]_B  \mprj_logic1[423]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[94]_A  net381 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[94]_B  \mprj_logic1[424]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[95]_A  net382 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[95]_B  \mprj_logic1[425]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[96]_A  net383 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[96]_B  \mprj_logic1[426]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[97]_A  net384 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[97]_B  \mprj_logic1[427]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[98]_A  net385 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[98]_B  \mprj_logic1[428]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[99]_A  net386 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[99]_B  \mprj_logic1[429]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[9]_A  net387 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_ena_buf[9]_B  \mprj_logic1[339]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[0]_A  net4 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[0]_B  \la_data_in_enable[0]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[100]_A  net5 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[100]_B  \la_data_in_enable[100]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[101]_A  net6 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[101]_B  \la_data_in_enable[101]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[102]_A  net7 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[102]_B  \la_data_in_enable[102]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[103]_A  net8 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[103]_B  \la_data_in_enable[103]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[104]_A  net9 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[104]_B  \la_data_in_enable[104]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[105]_A  net10 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[105]_B  \la_data_in_enable[105]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[106]_A  net11 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[106]_B  \la_data_in_enable[106]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[107]_A  net12 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[107]_B  \la_data_in_enable[107]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[108]_A  net13 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[108]_B  \la_data_in_enable[108]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[109]_A  net14 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[109]_B  \la_data_in_enable[109]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[10]_A  net15 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[10]_B  \la_data_in_enable[10]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[110]_A  net16 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[110]_B  \la_data_in_enable[110]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[111]_A  net17 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[111]_B  \la_data_in_enable[111]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[112]_A  net18 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[112]_B  \la_data_in_enable[112]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[113]_A  net19 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[113]_B  \la_data_in_enable[113]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[114]_A  net20 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[114]_B  \la_data_in_enable[114]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[115]_A  net21 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[115]_B  \la_data_in_enable[115]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[116]_A  net22 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[116]_B  \la_data_in_enable[116]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[117]_A  net23 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[117]_B  \la_data_in_enable[117]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[118]_A  net24 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[118]_B  \la_data_in_enable[118]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[119]_A  net25 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[119]_B  \la_data_in_enable[119]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[11]_A  net26 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[11]_B  \la_data_in_enable[11]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[120]_A  net27 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[120]_B  \la_data_in_enable[120]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[121]_A  net28 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[121]_B  \la_data_in_enable[121]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[122]_A  net29 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[122]_B  \la_data_in_enable[122]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[123]_A  net30 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[123]_B  \la_data_in_enable[123]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[124]_A  net31 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[124]_B  \la_data_in_enable[124]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[125]_A  net32 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[125]_B  \la_data_in_enable[125]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[126]_A  net33 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[126]_B  \la_data_in_enable[126]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[127]_A  net34 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[127]_B  \la_data_in_enable[127]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[12]_A  net35 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[12]_B  \la_data_in_enable[12]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[13]_A  net36 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[13]_B  \la_data_in_enable[13]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[14]_A  net37 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[14]_B  \la_data_in_enable[14]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[15]_A  net38 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[15]_B  \la_data_in_enable[15]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[16]_A  net39 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[16]_B  \la_data_in_enable[16]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[17]_A  net40 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[17]_B  \la_data_in_enable[17]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[18]_A  net41 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[18]_B  \la_data_in_enable[18]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[19]_A  net42 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[19]_B  \la_data_in_enable[19]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[1]_A  net43 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[1]_B  \la_data_in_enable[1]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[20]_A  net44 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[20]_B  \la_data_in_enable[20]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[21]_A  net45 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[21]_B  \la_data_in_enable[21]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[22]_A  net46 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[22]_B  \la_data_in_enable[22]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[23]_A  net47 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[23]_B  \la_data_in_enable[23]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[24]_A  net48 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[24]_B  \la_data_in_enable[24]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[25]_A  net49 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[25]_B  \la_data_in_enable[25]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[26]_A  net50 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[26]_B  \la_data_in_enable[26]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[27]_A  net51 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[27]_B  \la_data_in_enable[27]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[28]_A  net52 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[28]_B  \la_data_in_enable[28]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[29]_A  net53 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[29]_B  \la_data_in_enable[29]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[2]_A  net54 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[2]_B  \la_data_in_enable[2]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[30]_A  net55 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[30]_B  \la_data_in_enable[30]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[31]_A  net56 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[31]_B  \la_data_in_enable[31]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[32]_A  net57 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[32]_B  \la_data_in_enable[32]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[33]_A  net58 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[33]_B  \la_data_in_enable[33]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[34]_A  net59 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[34]_B  \la_data_in_enable[34]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[35]_A  net60 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[35]_B  \la_data_in_enable[35]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[36]_A  net61 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[36]_B  \la_data_in_enable[36]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[37]_A  net62 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[37]_B  \la_data_in_enable[37]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[38]_A  net63 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[38]_B  \la_data_in_enable[38]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[39]_A  net64 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[39]_B  \la_data_in_enable[39]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[3]_A  net65 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[3]_B  \la_data_in_enable[3]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[40]_A  net66 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[40]_B  \la_data_in_enable[40]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[41]_A  net67 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[41]_B  \la_data_in_enable[41]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[42]_A  net68 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[42]_B  \la_data_in_enable[42]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[43]_A  net69 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[43]_B  \la_data_in_enable[43]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[44]_A  net70 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[44]_B  \la_data_in_enable[44]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[45]_A  net71 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[45]_B  \la_data_in_enable[45]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[46]_A  net72 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[46]_B  \la_data_in_enable[46]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[47]_A  net73 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[47]_B  \la_data_in_enable[47]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[48]_A  net74 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[48]_B  \la_data_in_enable[48]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[49]_A  net75 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[49]_B  \la_data_in_enable[49]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[4]_A  net76 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[4]_B  \la_data_in_enable[4]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[50]_A  net77 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[50]_B  \la_data_in_enable[50]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[51]_A  net78 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[51]_B  \la_data_in_enable[51]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[52]_A  net79 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[52]_B  \la_data_in_enable[52]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[53]_A  net80 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[53]_B  \la_data_in_enable[53]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[54]_A  net81 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[54]_B  \la_data_in_enable[54]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[55]_A  net82 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[55]_B  \la_data_in_enable[55]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[56]_A  net83 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[56]_B  \la_data_in_enable[56]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[57]_A  net84 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[57]_B  \la_data_in_enable[57]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[58]_A  net85 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[58]_B  \la_data_in_enable[58]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[59]_A  net86 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[59]_B  \la_data_in_enable[59]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[5]_A  net87 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[5]_B  \la_data_in_enable[5]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[60]_A  net88 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[60]_B  \la_data_in_enable[60]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[61]_A  net89 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[61]_B  \la_data_in_enable[61]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[62]_A  net90 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[62]_B  \la_data_in_enable[62]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[63]_A  net91 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[63]_B  \la_data_in_enable[63]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[64]_A  net92 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[64]_B  \la_data_in_enable[64]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[65]_A  net93 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[65]_B  \la_data_in_enable[65]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[66]_A  net94 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[66]_B  \la_data_in_enable[66]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[67]_A  net95 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[67]_B  \la_data_in_enable[67]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[68]_A  net96 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[68]_B  \la_data_in_enable[68]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[69]_A  net97 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[69]_B  \la_data_in_enable[69]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[6]_A  net98 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[6]_B  \la_data_in_enable[6]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[70]_A  net99 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[70]_B  \la_data_in_enable[70]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[71]_A  net100 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[71]_B  \la_data_in_enable[71]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[72]_A  net101 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[72]_B  \la_data_in_enable[72]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[73]_A  net102 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[73]_B  \la_data_in_enable[73]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[74]_A  net103 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[74]_B  \la_data_in_enable[74]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[75]_A  net104 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[75]_B  \la_data_in_enable[75]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[76]_A  net105 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[76]_B  \la_data_in_enable[76]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[77]_A  net106 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[77]_B  \la_data_in_enable[77]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[78]_A  net107 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[78]_B  \la_data_in_enable[78]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[79]_A  net108 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[79]_B  \la_data_in_enable[79]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[7]_A  net109 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[7]_B  \la_data_in_enable[7]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[80]_A  net110 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[80]_B  \la_data_in_enable[80]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[81]_A  net111 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[81]_B  \la_data_in_enable[81]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[82]_A  net112 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[82]_B  \la_data_in_enable[82]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[83]_A  net113 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[83]_B  \la_data_in_enable[83]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[84]_A  net114 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[84]_B  \la_data_in_enable[84]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[85]_A  net115 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[85]_B  \la_data_in_enable[85]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[86]_A  net116 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[86]_B  \la_data_in_enable[86]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[87]_A  net117 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[87]_B  \la_data_in_enable[87]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[88]_A  net118 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[88]_B  \la_data_in_enable[88]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[89]_A  net119 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[89]_B  \la_data_in_enable[89]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[8]_A  net120 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[8]_B  \la_data_in_enable[8]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[90]_A  net121 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[90]_B  \la_data_in_enable[90]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[91]_A  net122 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[91]_B  \la_data_in_enable[91]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[92]_A  net123 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[92]_B  \la_data_in_enable[92]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[93]_A  net124 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[93]_B  \la_data_in_enable[93]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[94]_A  net125 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[94]_B  \la_data_in_enable[94]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[95]_A  net126 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[95]_B  \la_data_in_enable[95]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[96]_A  net127 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[96]_B  \la_data_in_enable[96]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[97]_A  net128 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[97]_B  \la_data_in_enable[97]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[98]_A  net129 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[98]_B  \la_data_in_enable[98]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[99]_A  net130 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[99]_B  \la_data_in_enable[99]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[9]_A  net131 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_in_gates[9]_B  \la_data_in_enable[9]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[0]_A  _201_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[0]_TE  \mprj_logic1[202]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[100]_A  _202_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[100]_TE  \mprj_logic1[302]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[101]_A  _203_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[101]_TE  \mprj_logic1[303]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[102]_A  _204_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[102]_TE  \mprj_logic1[304]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[103]_A  _205_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[103]_TE  \mprj_logic1[305]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[104]_A  _206_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[104]_TE  \mprj_logic1[306]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[105]_A  _207_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[105]_TE  \mprj_logic1[307]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[106]_A  _208_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[106]_TE  \mprj_logic1[308]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[107]_A  _209_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[107]_TE  \mprj_logic1[309]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[108]_A  _210_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[108]_TE  \mprj_logic1[310]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[109]_A  _211_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[109]_TE  \mprj_logic1[311]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[10]_A  _212_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[10]_TE  \mprj_logic1[212]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[110]_A  _213_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[110]_TE  \mprj_logic1[312]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[111]_A  _214_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[111]_TE  \mprj_logic1[313]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[112]_A  _215_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[112]_TE  \mprj_logic1[314]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[113]_A  _216_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[113]_TE  \mprj_logic1[315]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[114]_A  _217_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[114]_TE  \mprj_logic1[316]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[115]_A  _218_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[115]_TE  \mprj_logic1[317]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[116]_A  _219_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[116]_TE  \mprj_logic1[318]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[117]_A  _220_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[117]_TE  \mprj_logic1[319]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[118]_A  _221_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[118]_TE  \mprj_logic1[320]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[119]_A  _222_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[119]_TE  \mprj_logic1[321]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[11]_A  _223_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[11]_TE  \mprj_logic1[213]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[120]_A  _224_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[120]_TE  \mprj_logic1[322]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[121]_A  _225_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[121]_TE  \mprj_logic1[323]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[122]_A  _226_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[122]_TE  \mprj_logic1[324]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[123]_A  _227_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[123]_TE  \mprj_logic1[325]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[124]_A  _228_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[124]_TE  \mprj_logic1[326]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[125]_A  _229_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[125]_TE  \mprj_logic1[327]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[126]_A  _230_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[126]_TE  \mprj_logic1[328]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[127]_A  _231_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[127]_TE  \mprj_logic1[329]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[12]_A  _232_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[12]_TE  \mprj_logic1[214]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[13]_A  _233_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[13]_TE  \mprj_logic1[215]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[14]_A  _234_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[14]_TE  \mprj_logic1[216]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[15]_A  _235_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[15]_TE  \mprj_logic1[217]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[16]_A  _236_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[16]_TE  \mprj_logic1[218]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[17]_A  _237_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[17]_TE  \mprj_logic1[219]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[18]_A  _238_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[18]_TE  \mprj_logic1[220]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[19]_A  _239_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[19]_TE  \mprj_logic1[221]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[1]_A  _240_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[1]_TE  \mprj_logic1[203]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[20]_A  _241_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[20]_TE  \mprj_logic1[222]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[21]_A  _242_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[21]_TE  \mprj_logic1[223]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[22]_A  _243_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[22]_TE  \mprj_logic1[224]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[23]_A  _244_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[23]_TE  \mprj_logic1[225]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[24]_A  _245_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[24]_TE  \mprj_logic1[226]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[25]_A  _246_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[25]_TE  \mprj_logic1[227]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[26]_A  _247_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[26]_TE  \mprj_logic1[228]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[27]_A  _248_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[27]_TE  \mprj_logic1[229]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[28]_A  _249_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[28]_TE  \mprj_logic1[230]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[29]_A  _250_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[29]_TE  \mprj_logic1[231]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[2]_A  _251_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[2]_TE  \mprj_logic1[204]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[30]_A  _252_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[30]_TE  \mprj_logic1[232]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[31]_A  _253_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[31]_TE  \mprj_logic1[233]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[32]_A  _254_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[32]_TE  \mprj_logic1[234]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[33]_A  _255_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[33]_TE  \mprj_logic1[235]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[34]_A  _256_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[34]_TE  \mprj_logic1[236]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[35]_A  _257_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[35]_TE  \mprj_logic1[237]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[36]_A  _258_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[36]_TE  \mprj_logic1[238]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[37]_A  _259_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[37]_TE  \mprj_logic1[239]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[38]_A  _260_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[38]_TE  \mprj_logic1[240]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[39]_A  _261_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[39]_TE  \mprj_logic1[241]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[3]_A  _262_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[3]_TE  \mprj_logic1[205]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[40]_A  _263_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[40]_TE  \mprj_logic1[242]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[41]_A  _264_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[41]_TE  \mprj_logic1[243]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[42]_A  _265_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[42]_TE  \mprj_logic1[244]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[43]_A  _266_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[43]_TE  \mprj_logic1[245]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[44]_A  _267_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[44]_TE  \mprj_logic1[246]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[45]_A  _268_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[45]_TE  \mprj_logic1[247]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[46]_A  _269_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[46]_TE  \mprj_logic1[248]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[47]_A  _270_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[47]_TE  \mprj_logic1[249]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[48]_A  _271_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[48]_TE  \mprj_logic1[250]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[49]_A  _272_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[49]_TE  \mprj_logic1[251]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[4]_A  _273_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[4]_TE  \mprj_logic1[206]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[50]_A  _274_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[50]_TE  \mprj_logic1[252]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[51]_A  _275_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[51]_TE  \mprj_logic1[253]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[52]_A  _276_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[52]_TE  \mprj_logic1[254]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[53]_A  _277_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[53]_TE  \mprj_logic1[255]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[54]_A  _278_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[54]_TE  \mprj_logic1[256]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[55]_A  _279_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[55]_TE  \mprj_logic1[257]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[56]_A  _280_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[56]_TE  \mprj_logic1[258]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[57]_A  _281_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[57]_TE  \mprj_logic1[259]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[58]_A  _282_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[58]_TE  \mprj_logic1[260]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[59]_A  _283_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[59]_TE  \mprj_logic1[261]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[5]_A  _284_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[5]_TE  \mprj_logic1[207]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[60]_A  _285_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[60]_TE  \mprj_logic1[262]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[61]_A  _286_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[61]_TE  \mprj_logic1[263]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[62]_A  _287_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[62]_TE  \mprj_logic1[264]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[63]_A  _288_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[63]_TE  \mprj_logic1[265]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[64]_A  _289_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[64]_TE  \mprj_logic1[266]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[65]_A  _290_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[65]_TE  \mprj_logic1[267]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[66]_A  _291_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[66]_TE  \mprj_logic1[268]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[67]_A  _292_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[67]_TE  \mprj_logic1[269]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[68]_A  _293_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[68]_TE  \mprj_logic1[270]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[69]_A  _294_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[69]_TE  \mprj_logic1[271]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[6]_A  _295_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[6]_TE  \mprj_logic1[208]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[70]_A  _296_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[70]_TE  \mprj_logic1[272]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[71]_A  _297_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[71]_TE  \mprj_logic1[273]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[72]_A  _298_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[72]_TE  \mprj_logic1[274]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[73]_A  _299_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[73]_TE  \mprj_logic1[275]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[74]_A  _300_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[74]_TE  \mprj_logic1[276]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[75]_A  _301_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[75]_TE  \mprj_logic1[277]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[76]_A  _302_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[76]_TE  \mprj_logic1[278]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[77]_A  _303_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[77]_TE  \mprj_logic1[279]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[78]_A  _304_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[78]_TE  \mprj_logic1[280]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[79]_A  _305_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[79]_TE  \mprj_logic1[281]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[7]_A  _306_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[7]_TE  \mprj_logic1[209]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[80]_A  _307_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[80]_TE  \mprj_logic1[282]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[81]_A  _308_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[81]_TE  \mprj_logic1[283]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[82]_A  _309_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[82]_TE  \mprj_logic1[284]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[83]_A  _310_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[83]_TE  \mprj_logic1[285]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[84]_A  _311_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[84]_TE  \mprj_logic1[286]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[85]_A  _312_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[85]_TE  \mprj_logic1[287]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[86]_A  _313_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[86]_TE  \mprj_logic1[288]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[87]_A  _314_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[87]_TE  \mprj_logic1[289]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[88]_A  _315_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[88]_TE  \mprj_logic1[290]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[89]_A  _316_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[89]_TE  \mprj_logic1[291]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[8]_A  _317_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[8]_TE  \mprj_logic1[210]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[90]_A  _318_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[90]_TE  \mprj_logic1[292]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[91]_A  _319_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[91]_TE  \mprj_logic1[293]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[92]_A  _320_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[92]_TE  \mprj_logic1[294]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[93]_A  _321_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[93]_TE  \mprj_logic1[295]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[94]_A  _322_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[94]_TE  \mprj_logic1[296]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[95]_A  _323_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[95]_TE  \mprj_logic1[297]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[96]_A  _324_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[96]_TE  \mprj_logic1[298]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[97]_A  _325_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[97]_TE  \mprj_logic1[299]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[98]_A  _326_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[98]_TE  \mprj_logic1[300]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[99]_A  _327_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[99]_TE  \mprj_logic1[301]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[9]_A  _328_ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_to_mprj_oen_buffers[9]_TE  \mprj_logic1[211]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_wb_ena_buf_A net614 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_wb_ena_buf_B \mprj_logic1[462]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_ack_buffer_A mprj_ack_i_core_bar vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_ack_gate_A net516 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_ack_gate_B wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_buffers[0]_A  \mprj_dat_i_core_bar[0]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_buffers[10]_A  \mprj_dat_i_core_bar[10]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_buffers[11]_A  \mprj_dat_i_core_bar[11]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_buffers[12]_A  \mprj_dat_i_core_bar[12]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_buffers[13]_A  \mprj_dat_i_core_bar[13]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_buffers[14]_A  \mprj_dat_i_core_bar[14]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_buffers[15]_A  \mprj_dat_i_core_bar[15]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_buffers[16]_A  \mprj_dat_i_core_bar[16]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_buffers[17]_A  \mprj_dat_i_core_bar[17]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_buffers[18]_A  \mprj_dat_i_core_bar[18]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_buffers[19]_A  \mprj_dat_i_core_bar[19]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_buffers[1]_A  \mprj_dat_i_core_bar[1]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_buffers[20]_A  \mprj_dat_i_core_bar[20]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_buffers[21]_A  \mprj_dat_i_core_bar[21]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_buffers[22]_A  \mprj_dat_i_core_bar[22]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_buffers[23]_A  \mprj_dat_i_core_bar[23]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_buffers[24]_A  \mprj_dat_i_core_bar[24]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_buffers[25]_A  \mprj_dat_i_core_bar[25]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_buffers[26]_A  \mprj_dat_i_core_bar[26]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_buffers[27]_A  \mprj_dat_i_core_bar[27]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_buffers[28]_A  \mprj_dat_i_core_bar[28]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_buffers[29]_A  \mprj_dat_i_core_bar[29]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_buffers[2]_A  \mprj_dat_i_core_bar[2]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_buffers[30]_A  \mprj_dat_i_core_bar[30]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_buffers[31]_A  \mprj_dat_i_core_bar[31]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_buffers[3]_A  \mprj_dat_i_core_bar[3]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_buffers[4]_A  \mprj_dat_i_core_bar[4]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_buffers[5]_A  \mprj_dat_i_core_bar[5]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_buffers[6]_A  \mprj_dat_i_core_bar[6]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_buffers[7]_A  \mprj_dat_i_core_bar[7]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_buffers[8]_A  \mprj_dat_i_core_bar[8]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_buffers[9]_A  \mprj_dat_i_core_bar[9]\ vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[0]_A  net550 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[0]_B  wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[10]_A  net551 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[10]_B  wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[11]_A  net552 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[11]_B  wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[12]_A  net553 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[12]_B  wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[13]_A  net554 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[13]_B  wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[14]_A  net555 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[14]_B  wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[15]_A  net556 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[15]_B  wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[16]_A  net557 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[16]_B  wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[17]_A  net558 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[17]_B  wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[18]_A  net559 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[18]_B  wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[19]_A  net560 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[19]_B  wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[1]_A  net561 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[1]_B  wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[20]_A  net562 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[20]_B  wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[21]_A  net563 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[21]_B  wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[22]_A  net564 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[22]_B  wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[23]_A  net565 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[23]_B  wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[24]_A  net566 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[24]_B  wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[25]_A  net567 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[25]_B  wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[26]_A  net568 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[26]_B  wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[27]_A  net569 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[27]_B  wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[28]_A  net570 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[28]_B  wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[29]_A  net571 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[29]_B  wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[2]_A  net572 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[2]_B  wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[30]_A  net573 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[30]_B  wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[31]_A  net574 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[31]_B  wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[3]_A  net575 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[3]_B  wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[4]_A  net576 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[4]_B  wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[5]_A  net577 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[5]_B  wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[6]_A  net578 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[6]_B  wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[7]_A  net579 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[7]_B  wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[8]_A  net580 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[8]_B  wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[9]_A  net581 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X\ANTENNA_user_wb_dat_gates[9]_B  wb_in_enable vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1030 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1046 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1172 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1209 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1216 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1224 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1271 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1356 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1411 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1454 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1464 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1532 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1588 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1604 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1628 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1635 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1720 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1728 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1774 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1797 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1805 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1836 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1859 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1898 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1914 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1937 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1945 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1976 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_201 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2049 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2123 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2290 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2346 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_240 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_488 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_54 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_601 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_627 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_69 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_7 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_705 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_736 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_767 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_845 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_85 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_884 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_915 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_929 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1095 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1122 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1186 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1263 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1299 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1326 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1336 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1340 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1347 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1397 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1453 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1487 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1509 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1621 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1688 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1789 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1845 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1899 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1908 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1912 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1916 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1920 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1952 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1956 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_2007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_262 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_383 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_484 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_593 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_626 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_630 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_646 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_688 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_696 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_700 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_712 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_724 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_836 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_893 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_920 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_928 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_943 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_963 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1013 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1084 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1088 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1095 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1153 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1362 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1534 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1856 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1872 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_2007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_374 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_402 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_406 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_484 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_488 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_524 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_604 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_624 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_628 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_675 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_686 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_690 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_915 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_935 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1680 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1784 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1800 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_2007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_400 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_509 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_619 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1686 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1716 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1786 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1796 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1800 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1804 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1828 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1927 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1935 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1955 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_2007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_375 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_396 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_655 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1686 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1698 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1710 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1719 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_1743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_1767 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1775 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_1794 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1798 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_1923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1990 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_2002 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2008 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_604 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1578 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_1633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_2007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_271 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_568 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_584 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_612 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_620 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_630 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_657 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_731 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1619 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1635 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1646 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1686 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1775 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1796 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1800 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1871 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1898 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1999 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_402 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_584 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1749 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1772 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_2004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2008 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_618 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_634 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1556 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_1755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1759 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_1771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1786 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_1803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1888 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_1912 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_1935 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1938 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1968 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1971 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1993 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_354 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_370 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_591 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_713 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1663 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1747 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1822 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1859 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1884 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1887 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1906 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1910 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_2003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_243 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_35 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_542 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_564 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_568 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_576 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_61 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_65 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_738 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1004 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1019 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1027 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1032 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1036 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1040 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1050 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1054 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1068 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1072 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1076 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1080 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1089 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_11 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1103 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1124 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1128 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1132 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1140 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1168 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1172 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1181 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1187 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1243 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1256 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1260 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1360 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1364 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1368 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1380 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1384 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1405 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1488 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1492 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1496 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_15 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1504 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1508 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_153 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1550 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1590 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1598 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1608 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1612 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1616 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1629 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1663 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1678 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1685 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1690 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1705 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1712 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1748 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1752 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1756 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1760 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1767 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1776 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1787 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_180 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1826 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1830 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1834 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_184 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1860 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1864 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1868 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1872 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1876 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1880 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_19 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1900 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1926 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1938 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1965 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1991 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_200 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_204 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2094 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_2105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_2117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2152 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2156 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_2223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_2228 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_2245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2263 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2271 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2284 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2291 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_2326 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2350 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_244 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_25 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_260 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_264 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_288 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_29 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_299 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_319 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_326 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_33 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_368 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_37 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_372 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_376 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_403 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_43 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_434 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_438 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_452 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_461 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_47 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_492 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_496 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_509 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_536 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_543 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_551 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_57 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_574 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_578 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_61 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_620 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_624 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_628 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_649 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_65 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_660 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_668 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_686 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_691 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_702 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_71 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_732 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_736 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_749 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_75 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_760 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_768 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_775 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_789 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_79 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_802 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_815 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_833 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_845 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_87 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_870 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_880 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_884 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_888 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_901 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_91 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_915 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_935 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_940 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_944 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_948 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_95 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_957 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_965 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_984 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_988 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_99 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_1674 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1678 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1682 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_1728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1747 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1767 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_181 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1879 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_188 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1901 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_240 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_244 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_248 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_264 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_268 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_293 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_346 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_350 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_372 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_382 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_490 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_494 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1586 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1598 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_1655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_1753 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1820 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1824 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1912 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1920 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1924 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1928 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1940 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_2002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_2006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_232 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_236 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_240 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_318 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_396 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_403 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_537 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_570 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_680 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_696 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_708 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_89 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_1573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_1579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1590 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_1718 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1722 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1734 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_186 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1900 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1904 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1915 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1980 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_2008 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_624 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_674 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_686 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_1571 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1578 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1582 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_1717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_1727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1831 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_1848 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_1884 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_1941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_1997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_2004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2008 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_312 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_316 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_327 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_374 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_456 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_460 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_466 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_537 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_546 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_576 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_592 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_62 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_74 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_86 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_98 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1591 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1599 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_1663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_1727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1747 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_1803 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1850 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1870 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1887 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1915 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_1935 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1999 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2027 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2050 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2055 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_206 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_2079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2150 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2327 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_461 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_516 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_540 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_57 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_630 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_685 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_691 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_77 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1627 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1649 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1702 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1772 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_1804 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1828 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1873 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2011 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2041 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2100 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2187 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2248 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2322 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_264 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_438 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_656 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_660 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_1614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_1801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1843 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1850 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1942 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2090 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_2195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2299 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_2307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_466 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_551 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_560 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_592 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_596 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_628 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_632 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_705 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_738 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_74 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_78 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_10 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1764 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1843 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1934 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1938 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1991 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_2053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_2133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_22 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2290 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2324 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_299 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_34 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_433 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_46 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_512 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_516 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_54 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_57 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_590 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_6 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_61 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_67 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_705 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_82 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_94 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1027 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_148 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1508 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_156 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1772 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1780 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1788 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1956 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_215 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2300 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_523 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_724 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_75 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_79 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1089 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1460 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1492 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_160 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1621 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1691 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1712 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1942 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2004 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_2185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2246 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2316 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_236 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_47 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_572 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_65 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_724 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_738 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_74 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_78 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_90 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_10 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1000 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1020 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1027 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1062 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1083 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1124 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1128 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1132 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1186 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1216 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1236 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1240 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1244 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1265 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1268 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1280 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1288 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1292 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_130 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1308 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1327 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1346 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1350 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1364 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1368 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1394 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_14 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1424 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1433 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1439 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1453 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1461 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1492 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1496 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1516 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1520 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1523 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1545 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1572 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1601 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1616 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1620 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1668 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1676 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1682 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1686 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1691 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1702 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1713 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1752 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1762 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1787 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1796 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_18 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_180 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1800 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1804 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1808 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1812 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1816 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_184 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1843 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1852 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1864 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_188 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1881 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1892 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1908 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1927 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1965 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1980 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1993 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2004 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2012 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2016 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2020 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2024 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2032 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2039 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2049 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2058 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_206 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2066 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2072 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2124 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2136 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2178 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_22 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2244 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2299 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2322 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2348 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_26 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_29 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_322 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_33 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_369 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_372 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_376 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_388 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_444 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_45 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_508 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_512 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_516 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_524 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_564 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_59 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_593 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_6 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_606 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_618 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_63 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_655 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_675 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_68 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_684 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_688 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_705 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_716 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_72 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_720 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_744 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_748 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_752 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_761 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_772 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_803 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_822 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_826 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_85 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_853 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_873 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_888 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_89 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_900 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_934 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_938 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_942 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_965 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_97 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_971 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_990 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_996 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1130 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1201 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_131 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1453 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1478 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1657 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1678 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1682 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1702 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1774 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1814 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_184 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1843 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2095 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2200 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2263 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2319 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_326 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_442 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_55 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_60 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_710 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_72 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_798 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_80 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_820 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_824 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_836 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_881 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_932 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_960 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_976 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1027 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1030 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1042 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1130 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1150 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1548 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1842 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2103 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2320 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_318 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_35 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_462 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_495 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_60 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_66 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_76 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_798 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_823 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_859 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_881 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_888 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_929 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_983 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_99 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1030 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1244 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1460 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1464 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_148 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1761 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_179 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1810 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1832 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1836 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1916 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2131 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_296 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_327 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_350 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_383 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_406 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_495 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_607 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_628 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_63 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_705 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_77 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_775 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_887 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_937 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_943 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1150 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1158 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1388 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1621 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1700 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1713 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1899 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_214 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2263 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2324 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_47 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_542 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_57 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_63 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_67 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_70 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_815 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_906 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_92 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_922 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_934 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_96 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_965 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1369 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1534 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1629 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1742 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1746 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1752 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1760 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1904 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2041 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2049 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2060 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2128 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2181 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_2193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2276 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2284 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2320 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_369 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_444 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_601 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_663 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_744 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_78 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_82 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_838 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_850 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_858 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_862 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_904 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_91 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_95 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_99 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1049 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1083 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1244 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1453 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1632 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1733 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1759 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1769 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1899 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1970 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1986 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_201 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2060 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_215 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_2273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_237 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_328 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_433 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_649 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_67 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_853 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_868 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_976 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1075 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1264 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1290 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1366 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1769 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1808 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1812 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1952 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1964 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2004 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_201 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2040 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2072 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2088 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2209 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_369 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_428 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_551 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_61 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_657 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_770 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_798 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_85 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_852 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_92 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_96 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_100 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1013 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1083 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1090 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1263 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1378 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1394 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1509 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1712 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1775 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1805 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1844 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1912 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1952 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1984 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1999 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2062 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_2108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_2193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_220 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2214 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_2225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_228 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2322 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2350 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_545 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_691 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_71 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_859 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_909 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_96 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_103 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1300 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1489 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1508 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1636 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1761 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1915 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1920 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1963 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2077 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2322 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_439 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_686 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_79 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_833 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_845 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_882 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_898 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_970 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1018 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1034 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1046 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1058 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1083 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1104 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1327 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1508 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1537 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1652 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1753 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1759 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1922 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1928 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2047 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2080 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2088 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_220 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2265 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_243 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_584 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_677 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_69 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_767 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_91 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_95 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_988 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1027 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1088 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_11 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1128 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1168 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1243 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1263 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1326 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1412 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1434 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1466 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1480 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1486 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1543 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_16 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1608 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1648 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1668 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1685 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1732 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1753 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1787 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1968 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2030 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2042 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2067 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2094 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2122 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2180 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2348 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_252 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_276 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_28 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_324 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_355 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_375 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_40 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_593 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_64 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_68 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_682 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_705 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_724 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_749 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_80 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_850 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_906 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_92 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_922 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_934 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_957 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_963 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1015 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1072 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1088 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_1128 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1201 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1291 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1901 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_2033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2040 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_2085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_2145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2150 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_2197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2322 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_288 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_292 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_91 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_938 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_95 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1318 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1328 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1397 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1749 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1908 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1912 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1942 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_2037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2040 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_299 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_658 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_77 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_776 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_815 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_823 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_909 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_934 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_98 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1166 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1293 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1466 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1515 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1536 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1564 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1574 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_2189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_2357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_495 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_777 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_798 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_833 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_840 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_844 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_85 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_873 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_886 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_89 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1433 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1438 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1442 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1454 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1657 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1662 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1678 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1752 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1828 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1844 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2021 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2095 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_833 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_836 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_873 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1008 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1080 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1893 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2123 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_663 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_805 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_840 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_844 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_878 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_904 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_908 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_943 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_964 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_1112 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1201 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1216 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1220 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_1345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1542 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1558 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1578 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_2004 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2008 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_2012 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_2105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_2133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_354 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_370 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_85 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_93 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1012 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1153 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1439 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1584 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1749 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1909 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2022 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2048 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2088 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_803 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_915 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_955 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1090 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_11 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_1345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1496 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1596 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1677 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1888 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_1898 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_2017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2148 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_23 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2316 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2320 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_35 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_47 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_621 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_646 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_7 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_797 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_822 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_826 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_853 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_858 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_862 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_882 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_886 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_901 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_926 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_957 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1075 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_1452 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1537 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_2041 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_2123 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_2146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_2235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_2325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_607 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_1185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1208 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_1689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1704 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1719 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1810 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1822 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1834 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_1990 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2002 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2160 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_2273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_2283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_635 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_892 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_49_989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1013 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1019 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1044 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1048 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1096 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1100 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1236 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1240 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1433 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1489 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1516 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1614 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1629 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1753 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1768 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1861 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1870 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1927 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_2009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2187 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2355 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_300 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_487 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_649 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_733 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_736 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_775 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_836 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_840 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_844 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_932 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_940 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_943 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_962 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_1069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_1137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_1586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_1693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_1729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_1829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1843 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1970 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2030 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2066 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2090 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_2121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2136 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_2264 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_850 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_862 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_899 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_920 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_50_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1237 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1405 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1601 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1604 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1861 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1870 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1957 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2022 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2062 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_2081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2089 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2092 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2151 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2318 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_2346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2360 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_454 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_478 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_57 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_61 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_73 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_886 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_51_989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1055 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1216 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1220 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_128 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1326 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1366 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1377 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1405 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1416 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1537 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1550 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1570 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1586 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1636 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1648 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1663 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1749 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1762 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_186 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1872 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_19 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1962 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_1975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2008 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2024 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2040 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_3 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_448 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_462 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_61 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_67 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_7 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_79 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_52_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_53_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1052 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_1071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1103 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1131 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1168 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1215 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1240 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1244 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1248 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1284 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1298 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1328 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1444 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_1463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1495 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_1502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1523 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1560 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_1575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1618 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1632 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1676 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1691 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1713 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1720 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1724 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1749 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1836 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_1855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1887 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1898 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1915 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1952 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2010 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2024 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2032 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2039 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2054 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2058 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2068 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2083 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2112 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2209 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2228 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2290 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_23 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2344 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2348 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_453 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_514 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_543 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_57 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_572 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_602 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_61 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_629 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_660 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_711 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_718 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_722 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_739 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_747 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_75 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_776 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_805 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_848 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_856 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_892 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_906 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_935 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_94 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_965 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_98 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_994 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1088 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1100 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1104 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1140 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1431 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1484 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1492 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1496 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_159 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1601 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1620 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_2059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2103 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_2115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2122 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_2193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2208 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_2212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_2220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_2363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_254 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_77 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_864 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_868 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_904 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_99 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1006 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_104 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1047 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1179 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1187 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1268 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1284 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1336 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1355 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1404 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1408 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1502 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1544 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1548 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1560 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1564 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1592 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1828 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1844 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2054 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2058 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2070 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2094 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_214 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_2359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_49 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_495 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_59 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_63 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_652 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_67 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_70 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_731 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_74 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_761 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_769 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_80 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_842 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_915 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_92 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_96 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_993 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_10 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1018 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1299 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1369 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1593 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1784 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2062 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_22 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2248 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_53 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_568 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_6 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_68 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_80 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1004 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1156 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1160 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1172 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1264 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1268 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1293 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1453 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1619 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1636 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1658 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1662 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1733 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1761 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1769 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1789 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1845 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1901 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1927 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_2007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_571 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_700 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_712 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_724 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_796 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_800 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_804 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_844 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_892 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_963 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1015 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1064 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1068 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1083 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1095 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1130 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1152 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1208 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1235 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1320 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1347 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1480 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1537 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1574 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1578 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1627 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1705 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1716 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1873 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1929 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_2007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_369 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_380 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_403 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_416 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_546 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_578 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_685 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_753 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_808 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_851 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_870 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_898 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_914 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_920 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_934 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_0 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_1 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_10 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_11 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_12 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_13 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_14 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_16 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_17 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_18 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_19 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_2 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_20 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_21 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_22 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_23 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_24 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_25 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_26 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_28 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_31 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_33 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_34 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_35 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_36 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_37 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_38 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_4 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_40 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_42 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_43 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_44 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_45 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_46 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_47 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_48 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_49 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_5 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_50 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_52 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_54 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_55 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_56 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_59 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_6 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_60 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_61 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_62 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_63 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_64 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_67 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_68 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_7 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_71 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_72 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_73 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_74 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_75 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_76 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_78 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_79 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_8 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_80 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_82 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_83 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_84 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_86 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_88 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_89 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_9 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_90 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_91 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_92 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_94 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_95 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_96 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_98 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_99 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1000 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1003 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1004 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1009 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1012 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1019 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1030 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1031 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1040 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1046 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1082 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1090 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1091 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1104 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1105 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1109 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1119 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1139 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1140 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1150 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1155 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1174 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1182 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1189 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1190 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1191 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1193 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_140 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_150 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_159 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_160 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1725 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1734 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1739 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1748 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1752 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1757 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1759 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1766 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1767 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1769 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1770 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1775 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1779 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1784 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1789 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1790 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1791 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1793 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1794 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1795 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1797 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1798 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1799 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_180 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1800 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1806 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1807 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1809 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1824 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1829 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1833 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1834 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1842 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1843 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1845 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1857 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1859 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1866 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1867 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1869 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1870 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1874 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1875 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1877 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1879 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1880 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1883 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1884 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1889 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1890 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1891 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1892 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1893 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1894 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1895 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1897 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1898 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1899 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_190 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1906 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1907 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1908 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1909 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1915 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1919 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1924 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1929 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1947 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1949 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1957 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1958 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1960 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1967 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1968 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1970 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1974 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1976 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1977 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1979 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1980 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1986 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1990 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1993 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1994 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1996 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1997 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1998 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2000 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2001 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2002 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2003 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2004 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2005 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2006 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2007 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2008 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2009 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2010 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2016 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2019 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2020 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2021 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2030 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2033 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2039 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2040 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2042 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2049 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2050 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2051 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2058 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2060 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2061 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2062 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2067 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2070 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2076 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2080 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2085 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2090 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2091 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2092 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2094 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2099 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2100 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2101 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2102 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2103 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2104 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2105 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2106 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2107 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2108 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2109 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2110 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2116 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2117 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2119 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2120 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2130 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2136 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2137 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2140 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2141 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2150 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2160 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2161 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2162 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2164 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2169 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2170 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2171 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2173 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2180 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2182 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2190 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2191 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_760 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_790 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_800 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_801 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_807 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_808 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_809 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_810 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_870 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_880 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_890 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_896 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_900 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_901 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_907 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_908 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_909 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_910 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_925 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_961 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_969 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_970 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_980 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_989 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_990 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_998 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_329_ net478 vssd vssd vccd vccd _291_ sky130_fd_sc_hd__inv_2
X_330_ net479 vssd vssd vccd vccd _292_ sky130_fd_sc_hd__clkinv_2
X_331_ net480 vssd vssd vccd vccd _293_ sky130_fd_sc_hd__inv_2
X_332_ net481 vssd vssd vccd vccd _294_ sky130_fd_sc_hd__inv_2
X_333_ net483 vssd vssd vccd vccd _296_ sky130_fd_sc_hd__clkinv_2
X_334_ net484 vssd vssd vccd vccd _297_ sky130_fd_sc_hd__clkinv_2
X_335_ net485 vssd vssd vccd vccd _298_ sky130_fd_sc_hd__clkinv_2
X_336_ net486 vssd vssd vccd vccd _299_ sky130_fd_sc_hd__clkinv_2
X_337_ net487 vssd vssd vccd vccd _300_ sky130_fd_sc_hd__clkinv_2
X_338_ net488 vssd vssd vccd vccd _301_ sky130_fd_sc_hd__clkinv_2
X_339_ net489 vssd vssd vccd vccd _302_ sky130_fd_sc_hd__inv_2
X_340_ net490 vssd vssd vccd vccd _303_ sky130_fd_sc_hd__clkinv_2
X_341_ net491 vssd vssd vccd vccd _304_ sky130_fd_sc_hd__clkinv_2
X_342_ net492 vssd vssd vccd vccd _305_ sky130_fd_sc_hd__clkinv_2
X_343_ net494 vssd vssd vccd vccd _307_ sky130_fd_sc_hd__clkinv_2
X_344_ net495 vssd vssd vccd vccd _308_ sky130_fd_sc_hd__inv_2
X_345_ net496 vssd vssd vccd vccd _309_ sky130_fd_sc_hd__clkinv_2
X_346_ net497 vssd vssd vccd vccd _310_ sky130_fd_sc_hd__clkinv_2
X_347_ net498 vssd vssd vccd vccd _311_ sky130_fd_sc_hd__inv_2
X_348_ net499 vssd vssd vccd vccd _312_ sky130_fd_sc_hd__inv_2
X_349_ net500 vssd vssd vccd vccd _313_ sky130_fd_sc_hd__inv_2
X_350_ net501 vssd vssd vccd vccd _314_ sky130_fd_sc_hd__inv_2
X_351_ net502 vssd vssd vccd vccd _315_ sky130_fd_sc_hd__inv_2
X_352_ net503 vssd vssd vccd vccd _316_ sky130_fd_sc_hd__clkinv_2
X_353_ net505 vssd vssd vccd vccd _318_ sky130_fd_sc_hd__clkinv_2
X_354_ net506 vssd vssd vccd vccd _319_ sky130_fd_sc_hd__clkinv_2
X_355_ net507 vssd vssd vccd vccd _320_ sky130_fd_sc_hd__clkinv_2
X_356_ net508 vssd vssd vccd vccd _321_ sky130_fd_sc_hd__inv_2
X_357_ net509 vssd vssd vccd vccd _322_ sky130_fd_sc_hd__inv_2
X_358_ net510 vssd vssd vccd vccd _323_ sky130_fd_sc_hd__inv_2
X_359_ net511 vssd vssd vccd vccd _324_ sky130_fd_sc_hd__inv_2
X_360_ net512 vssd vssd vccd vccd _325_ sky130_fd_sc_hd__inv_2
X_361_ net513 vssd vssd vccd vccd _326_ sky130_fd_sc_hd__inv_2
X_362_ net514 vssd vssd vccd vccd _327_ sky130_fd_sc_hd__inv_2
X_363_ net389 vssd vssd vccd vccd _202_ sky130_fd_sc_hd__inv_2
X_364_ net390 vssd vssd vccd vccd _203_ sky130_fd_sc_hd__clkinv_2
X_365_ net391 vssd vssd vccd vccd _204_ sky130_fd_sc_hd__inv_2
X_366_ net392 vssd vssd vccd vccd _205_ sky130_fd_sc_hd__clkinv_2
X_367_ net393 vssd vssd vccd vccd _206_ sky130_fd_sc_hd__clkinv_2
X_368_ net394 vssd vssd vccd vccd _207_ sky130_fd_sc_hd__inv_2
X_369_ net395 vssd vssd vccd vccd _208_ sky130_fd_sc_hd__clkinv_2
X_370_ net396 vssd vssd vccd vccd _209_ sky130_fd_sc_hd__inv_2
X_371_ net397 vssd vssd vccd vccd _210_ sky130_fd_sc_hd__inv_2
X_372_ net398 vssd vssd vccd vccd _211_ sky130_fd_sc_hd__inv_2
X_373_ net400 vssd vssd vccd vccd _213_ sky130_fd_sc_hd__inv_2
X_374_ net401 vssd vssd vccd vccd _214_ sky130_fd_sc_hd__inv_2
X_375_ net402 vssd vssd vccd vccd _215_ sky130_fd_sc_hd__inv_2
X_376_ net403 vssd vssd vccd vccd _216_ sky130_fd_sc_hd__inv_2
X_377_ net404 vssd vssd vccd vccd _217_ sky130_fd_sc_hd__inv_2
X_378_ net405 vssd vssd vccd vccd _218_ sky130_fd_sc_hd__clkinv_2
X_379_ net406 vssd vssd vccd vccd _219_ sky130_fd_sc_hd__clkinv_2
X_380_ net407 vssd vssd vccd vccd _220_ sky130_fd_sc_hd__inv_2
X_381_ net408 vssd vssd vccd vccd _221_ sky130_fd_sc_hd__inv_2
X_382_ net409 vssd vssd vccd vccd _222_ sky130_fd_sc_hd__clkinv_2
X_383_ net411 vssd vssd vccd vccd _224_ sky130_fd_sc_hd__inv_2
X_384_ net412 vssd vssd vccd vccd _225_ sky130_fd_sc_hd__clkinv_2
X_385_ net413 vssd vssd vccd vccd _226_ sky130_fd_sc_hd__clkinv_2
X_386_ net414 vssd vssd vccd vccd _227_ sky130_fd_sc_hd__clkinv_2
X_387_ net415 vssd vssd vccd vccd _228_ sky130_fd_sc_hd__inv_2
X_388_ net416 vssd vssd vccd vccd _229_ sky130_fd_sc_hd__clkinv_2
X_389_ net417 vssd vssd vccd vccd _230_ sky130_fd_sc_hd__inv_2
X_390_ net418 vssd vssd vccd vccd _231_ sky130_fd_sc_hd__inv_2
X_391_ net1 vssd vssd vccd vccd _000_ sky130_fd_sc_hd__clkinv_2
X_392_ net2 vssd vssd vccd vccd _001_ sky130_fd_sc_hd__inv_2
X_393_ net549 vssd vssd vccd vccd _002_ sky130_fd_sc_hd__inv_6
X_394_ net619 vssd vssd vccd vccd _003_ sky130_fd_sc_hd__inv_2
X_395_ net620 vssd vssd vccd vccd _004_ sky130_fd_sc_hd__clkinv_2
X_396_ net615 vssd vssd vccd vccd _005_ sky130_fd_sc_hd__clkinv_2
X_397_ net616 vssd vssd vccd vccd _006_ sky130_fd_sc_hd__inv_2
X_398_ net617 vssd vssd vccd vccd _007_ sky130_fd_sc_hd__clkinv_2
X_399_ net618 vssd vssd vccd vccd _008_ sky130_fd_sc_hd__clkinv_2
X_400_ net517 vssd vssd vccd vccd _009_ sky130_fd_sc_hd__clkinv_2
X_401_ net528 vssd vssd vccd vccd _020_ sky130_fd_sc_hd__inv_12
X_402_ net539 vssd vssd vccd vccd _031_ sky130_fd_sc_hd__inv_2
X_403_ net542 vssd vssd vccd vccd _034_ sky130_fd_sc_hd__inv_12
X_404_ net543 vssd vssd vccd vccd _035_ sky130_fd_sc_hd__inv_2
X_405_ net544 vssd vssd vccd vccd _036_ sky130_fd_sc_hd__inv_16
X_406_ net545 vssd vssd vccd vccd _037_ sky130_fd_sc_hd__clkinv_8
X_407_ net546 vssd vssd vccd vccd _038_ sky130_fd_sc_hd__inv_8
X_408_ net547 vssd vssd vccd vccd _039_ sky130_fd_sc_hd__clkinv_16
X_409_ net548 vssd vssd vccd vccd _040_ sky130_fd_sc_hd__inv_8
X_410_ net518 vssd vssd vccd vccd _010_ sky130_fd_sc_hd__inv_2
X_411_ net519 vssd vssd vccd vccd _011_ sky130_fd_sc_hd__inv_4
X_412_ net520 vssd vssd vccd vccd _012_ sky130_fd_sc_hd__inv_12
X_413_ net521 vssd vssd vccd vccd _013_ sky130_fd_sc_hd__inv_6
X_414_ net522 vssd vssd vccd vccd _014_ sky130_fd_sc_hd__clkinv_8
X_415_ net523 vssd vssd vccd vccd _015_ sky130_fd_sc_hd__inv_12
X_416_ net524 vssd vssd vccd vccd _016_ sky130_fd_sc_hd__inv_12
X_417_ net525 vssd vssd vccd vccd _017_ sky130_fd_sc_hd__inv_6
X_418_ net526 vssd vssd vccd vccd _018_ sky130_fd_sc_hd__inv_12
X_419_ net527 vssd vssd vccd vccd _019_ sky130_fd_sc_hd__inv_16
X_420_ net529 vssd vssd vccd vccd _021_ sky130_fd_sc_hd__clkinv_8
X_421_ net530 vssd vssd vccd vccd _022_ sky130_fd_sc_hd__inv_12
X_422_ net531 vssd vssd vccd vccd _023_ sky130_fd_sc_hd__inv_6
X_423_ net532 vssd vssd vccd vccd _024_ sky130_fd_sc_hd__inv_8
X_424_ net533 vssd vssd vccd vccd _025_ sky130_fd_sc_hd__clkinv_16
X_425_ net534 vssd vssd vccd vccd _026_ sky130_fd_sc_hd__inv_12
X_426_ net535 vssd vssd vccd vccd _027_ sky130_fd_sc_hd__inv_12
X_427_ net536 vssd vssd vccd vccd _028_ sky130_fd_sc_hd__clkinv_8
X_428_ net537 vssd vssd vccd vccd _029_ sky130_fd_sc_hd__inv_8
X_429_ net538 vssd vssd vccd vccd _030_ sky130_fd_sc_hd__inv_8
X_430_ net540 vssd vssd vccd vccd _032_ sky130_fd_sc_hd__clkinv_8
X_431_ net541 vssd vssd vccd vccd _033_ sky130_fd_sc_hd__inv_8
X_432_ net582 vssd vssd vccd vccd _041_ sky130_fd_sc_hd__clkinv_2
X_433_ net593 vssd vssd vccd vccd _052_ sky130_fd_sc_hd__inv_2
X_434_ net604 vssd vssd vccd vccd _063_ sky130_fd_sc_hd__inv_2
X_435_ net607 vssd vssd vccd vccd _066_ sky130_fd_sc_hd__inv_2
X_436_ net608 vssd vssd vccd vccd _067_ sky130_fd_sc_hd__clkinv_2
X_437_ net609 vssd vssd vccd vccd _068_ sky130_fd_sc_hd__inv_2
X_438_ net610 vssd vssd vccd vccd _069_ sky130_fd_sc_hd__inv_2
X_439_ net611 vssd vssd vccd vccd _070_ sky130_fd_sc_hd__clkinv_2
X_440_ net612 vssd vssd vccd vccd _071_ sky130_fd_sc_hd__inv_2
X_441_ net613 vssd vssd vccd vccd _072_ sky130_fd_sc_hd__clkinv_4
X_442_ net583 vssd vssd vccd vccd _042_ sky130_fd_sc_hd__clkinv_4
X_443_ net584 vssd vssd vccd vccd _043_ sky130_fd_sc_hd__clkinv_2
X_444_ net585 vssd vssd vccd vccd _044_ sky130_fd_sc_hd__clkinv_2
X_445_ net586 vssd vssd vccd vccd _045_ sky130_fd_sc_hd__clkinv_4
X_446_ net587 vssd vssd vccd vccd _046_ sky130_fd_sc_hd__clkinv_4
X_447_ net588 vssd vssd vccd vccd _047_ sky130_fd_sc_hd__clkinv_4
X_448_ net589 vssd vssd vccd vccd _048_ sky130_fd_sc_hd__clkinv_2
X_449_ net590 vssd vssd vccd vccd _049_ sky130_fd_sc_hd__inv_4
X_450_ net591 vssd vssd vccd vccd _050_ sky130_fd_sc_hd__inv_4
X_451_ net592 vssd vssd vccd vccd _051_ sky130_fd_sc_hd__inv_4
X_452_ net594 vssd vssd vccd vccd _053_ sky130_fd_sc_hd__inv_4
X_453_ net595 vssd vssd vccd vccd _054_ sky130_fd_sc_hd__inv_4
X_454_ net596 vssd vssd vccd vccd _055_ sky130_fd_sc_hd__inv_4
X_455_ net597 vssd vssd vccd vccd _056_ sky130_fd_sc_hd__inv_6
X_456_ net598 vssd vssd vccd vccd _057_ sky130_fd_sc_hd__inv_4
X_457_ net599 vssd vssd vccd vccd _058_ sky130_fd_sc_hd__inv_2
X_458_ net600 vssd vssd vccd vccd _059_ sky130_fd_sc_hd__inv_4
X_459_ net601 vssd vssd vccd vccd _060_ sky130_fd_sc_hd__inv_6
X_460_ net602 vssd vssd vccd vccd _061_ sky130_fd_sc_hd__clkinv_4
X_461_ net603 vssd vssd vccd vccd _062_ sky130_fd_sc_hd__clkinv_4
X_462_ net605 vssd vssd vccd vccd _064_ sky130_fd_sc_hd__inv_6
X_463_ net606 vssd vssd vccd vccd _065_ sky130_fd_sc_hd__clkinv_4
X_464_ net132 vssd vssd vccd vccd _073_ sky130_fd_sc_hd__inv_2
X_465_ net171 vssd vssd vccd vccd _112_ sky130_fd_sc_hd__clkinv_2
X_466_ net182 vssd vssd vccd vccd _123_ sky130_fd_sc_hd__clkinv_2
X_467_ net193 vssd vssd vccd vccd _134_ sky130_fd_sc_hd__clkinv_2
X_468_ net204 vssd vssd vccd vccd _145_ sky130_fd_sc_hd__clkinv_2
X_469_ net215 vssd vssd vccd vccd _156_ sky130_fd_sc_hd__inv_2
X_470_ net226 vssd vssd vccd vccd _167_ sky130_fd_sc_hd__inv_2
X_471_ net237 vssd vssd vccd vccd _178_ sky130_fd_sc_hd__clkinv_2
X_472_ net248 vssd vssd vccd vccd _189_ sky130_fd_sc_hd__inv_2
X_473_ net259 vssd vssd vccd vccd _200_ sky130_fd_sc_hd__clkinv_2
X_474_ net143 vssd vssd vccd vccd _084_ sky130_fd_sc_hd__clkinv_2
X_475_ net154 vssd vssd vccd vccd _095_ sky130_fd_sc_hd__clkinv_2
X_476_ net163 vssd vssd vccd vccd _104_ sky130_fd_sc_hd__clkinv_2
X_477_ net164 vssd vssd vccd vccd _105_ sky130_fd_sc_hd__clkinv_2
X_478_ net165 vssd vssd vccd vccd _106_ sky130_fd_sc_hd__inv_2
X_479_ net166 vssd vssd vccd vccd _107_ sky130_fd_sc_hd__inv_2
X_480_ net167 vssd vssd vccd vccd _108_ sky130_fd_sc_hd__clkinv_2
X_481_ net168 vssd vssd vccd vccd _109_ sky130_fd_sc_hd__clkinv_2
X_482_ net169 vssd vssd vccd vccd _110_ sky130_fd_sc_hd__clkinv_2
X_483_ net170 vssd vssd vccd vccd _111_ sky130_fd_sc_hd__inv_2
X_484_ net172 vssd vssd vccd vccd _113_ sky130_fd_sc_hd__inv_2
X_485_ net173 vssd vssd vccd vccd _114_ sky130_fd_sc_hd__clkinv_2
X_486_ net174 vssd vssd vccd vccd _115_ sky130_fd_sc_hd__clkinv_2
X_487_ net175 vssd vssd vccd vccd _116_ sky130_fd_sc_hd__clkinv_2
X_488_ net176 vssd vssd vccd vccd _117_ sky130_fd_sc_hd__inv_2
X_489_ net177 vssd vssd vccd vccd _118_ sky130_fd_sc_hd__clkinv_2
X_490_ net178 vssd vssd vccd vccd _119_ sky130_fd_sc_hd__inv_2
X_491_ net179 vssd vssd vccd vccd _120_ sky130_fd_sc_hd__clkinv_2
X_492_ net180 vssd vssd vccd vccd _121_ sky130_fd_sc_hd__inv_2
X_493_ net181 vssd vssd vccd vccd _122_ sky130_fd_sc_hd__clkinv_2
X_494_ net183 vssd vssd vccd vccd _124_ sky130_fd_sc_hd__clkinv_2
X_495_ net184 vssd vssd vccd vccd _125_ sky130_fd_sc_hd__clkinv_2
X_496_ net185 vssd vssd vccd vccd _126_ sky130_fd_sc_hd__clkinv_2
X_497_ net186 vssd vssd vccd vccd _127_ sky130_fd_sc_hd__clkinv_2
X_498_ net187 vssd vssd vccd vccd _128_ sky130_fd_sc_hd__clkinv_2
X_499_ net188 vssd vssd vccd vccd _129_ sky130_fd_sc_hd__clkinv_2
X_500_ net189 vssd vssd vccd vccd _130_ sky130_fd_sc_hd__clkinv_2
X_501_ net190 vssd vssd vccd vccd _131_ sky130_fd_sc_hd__clkinv_2
X_502_ net191 vssd vssd vccd vccd _132_ sky130_fd_sc_hd__inv_2
X_503_ net192 vssd vssd vccd vccd _133_ sky130_fd_sc_hd__clkinv_2
X_504_ net194 vssd vssd vccd vccd _135_ sky130_fd_sc_hd__inv_2
X_505_ net195 vssd vssd vccd vccd _136_ sky130_fd_sc_hd__clkinv_2
X_506_ net196 vssd vssd vccd vccd _137_ sky130_fd_sc_hd__clkinv_2
X_507_ net197 vssd vssd vccd vccd _138_ sky130_fd_sc_hd__clkinv_2
X_508_ net198 vssd vssd vccd vccd _139_ sky130_fd_sc_hd__clkinv_2
X_509_ net199 vssd vssd vccd vccd _140_ sky130_fd_sc_hd__inv_2
X_510_ net200 vssd vssd vccd vccd _141_ sky130_fd_sc_hd__clkinv_2
X_511_ net201 vssd vssd vccd vccd _142_ sky130_fd_sc_hd__clkinv_2
X_512_ net202 vssd vssd vccd vccd _143_ sky130_fd_sc_hd__clkinv_2
X_513_ net203 vssd vssd vccd vccd _144_ sky130_fd_sc_hd__clkinv_2
X_514_ net205 vssd vssd vccd vccd _146_ sky130_fd_sc_hd__clkinv_2
X_515_ net206 vssd vssd vccd vccd _147_ sky130_fd_sc_hd__clkinv_2
X_516_ net207 vssd vssd vccd vccd _148_ sky130_fd_sc_hd__inv_2
X_517_ net208 vssd vssd vccd vccd _149_ sky130_fd_sc_hd__clkinv_2
X_518_ net209 vssd vssd vccd vccd _150_ sky130_fd_sc_hd__inv_2
X_519_ net210 vssd vssd vccd vccd _151_ sky130_fd_sc_hd__clkinv_2
X_520_ net211 vssd vssd vccd vccd _152_ sky130_fd_sc_hd__clkinv_2
X_521_ net212 vssd vssd vccd vccd _153_ sky130_fd_sc_hd__inv_2
X_522_ net213 vssd vssd vccd vccd _154_ sky130_fd_sc_hd__inv_2
X_523_ net214 vssd vssd vccd vccd _155_ sky130_fd_sc_hd__clkinv_2
X_524_ net216 vssd vssd vccd vccd _157_ sky130_fd_sc_hd__inv_2
X_525_ net217 vssd vssd vccd vccd _158_ sky130_fd_sc_hd__inv_2
X_526_ net218 vssd vssd vccd vccd _159_ sky130_fd_sc_hd__clkinv_2
X_527_ net219 vssd vssd vccd vccd _160_ sky130_fd_sc_hd__clkinv_2
X_528_ net220 vssd vssd vccd vccd _161_ sky130_fd_sc_hd__clkinv_2
X_529_ net221 vssd vssd vccd vccd _162_ sky130_fd_sc_hd__clkinv_2
X_530_ net222 vssd vssd vccd vccd _163_ sky130_fd_sc_hd__clkinv_2
X_531_ net223 vssd vssd vccd vccd _164_ sky130_fd_sc_hd__inv_2
X_532_ net224 vssd vssd vccd vccd _165_ sky130_fd_sc_hd__clkinv_2
X_533_ net225 vssd vssd vccd vccd _166_ sky130_fd_sc_hd__clkinv_2
X_534_ net227 vssd vssd vccd vccd _168_ sky130_fd_sc_hd__clkinv_2
X_535_ net228 vssd vssd vccd vccd _169_ sky130_fd_sc_hd__inv_2
X_536_ net229 vssd vssd vccd vccd _170_ sky130_fd_sc_hd__clkinv_2
X_537_ net230 vssd vssd vccd vccd _171_ sky130_fd_sc_hd__inv_2
X_538_ net231 vssd vssd vccd vccd _172_ sky130_fd_sc_hd__clkinv_2
X_539_ net232 vssd vssd vccd vccd _173_ sky130_fd_sc_hd__inv_2
X_540_ net233 vssd vssd vccd vccd _174_ sky130_fd_sc_hd__clkinv_2
X_541_ net234 vssd vssd vccd vccd _175_ sky130_fd_sc_hd__inv_2
X_542_ net235 vssd vssd vccd vccd _176_ sky130_fd_sc_hd__clkinv_2
X_543_ net236 vssd vssd vccd vccd _177_ sky130_fd_sc_hd__clkinv_2
X_544_ net238 vssd vssd vccd vccd _179_ sky130_fd_sc_hd__clkinv_2
X_545_ net239 vssd vssd vccd vccd _180_ sky130_fd_sc_hd__clkinv_2
X_546_ net240 vssd vssd vccd vccd _181_ sky130_fd_sc_hd__clkinv_2
X_547_ net241 vssd vssd vccd vccd _182_ sky130_fd_sc_hd__clkinv_2
X_548_ net242 vssd vssd vccd vccd _183_ sky130_fd_sc_hd__clkinv_2
X_549_ net243 vssd vssd vccd vccd _184_ sky130_fd_sc_hd__clkinv_2
X_550_ net244 vssd vssd vccd vccd _185_ sky130_fd_sc_hd__inv_2
X_551_ net245 vssd vssd vccd vccd _186_ sky130_fd_sc_hd__inv_2
X_552_ net246 vssd vssd vccd vccd _187_ sky130_fd_sc_hd__clkinv_2
X_553_ net247 vssd vssd vccd vccd _188_ sky130_fd_sc_hd__inv_2
X_554_ net249 vssd vssd vccd vccd _190_ sky130_fd_sc_hd__inv_2
X_555_ net250 vssd vssd vccd vccd _191_ sky130_fd_sc_hd__inv_2
X_556_ net251 vssd vssd vccd vccd _192_ sky130_fd_sc_hd__inv_2
X_557_ net252 vssd vssd vccd vccd _193_ sky130_fd_sc_hd__clkinv_2
X_558_ net253 vssd vssd vccd vccd _194_ sky130_fd_sc_hd__inv_2
X_559_ net254 vssd vssd vccd vccd _195_ sky130_fd_sc_hd__inv_2
X_560_ net255 vssd vssd vccd vccd _196_ sky130_fd_sc_hd__clkinv_2
X_561_ net256 vssd vssd vccd vccd _197_ sky130_fd_sc_hd__clkinv_4
X_562_ net257 vssd vssd vccd vccd _198_ sky130_fd_sc_hd__clkinv_2
X_563_ net258 vssd vssd vccd vccd _199_ sky130_fd_sc_hd__clkinv_2
X_564_ net133 vssd vssd vccd vccd _074_ sky130_fd_sc_hd__inv_2
X_565_ net134 vssd vssd vccd vccd _075_ sky130_fd_sc_hd__clkinv_2
X_566_ net135 vssd vssd vccd vccd _076_ sky130_fd_sc_hd__inv_2
X_567_ net136 vssd vssd vccd vccd _077_ sky130_fd_sc_hd__clkinv_2
X_568_ net137 vssd vssd vccd vccd _078_ sky130_fd_sc_hd__clkinv_2
X_569_ net138 vssd vssd vccd vccd _079_ sky130_fd_sc_hd__clkinv_2
X_570_ net139 vssd vssd vccd vccd _080_ sky130_fd_sc_hd__clkinv_2
X_571_ net140 vssd vssd vccd vccd _081_ sky130_fd_sc_hd__inv_2
X_572_ net141 vssd vssd vccd vccd _082_ sky130_fd_sc_hd__inv_2
X_573_ net142 vssd vssd vccd vccd _083_ sky130_fd_sc_hd__inv_2
X_574_ net144 vssd vssd vccd vccd _085_ sky130_fd_sc_hd__inv_2
X_575_ net145 vssd vssd vccd vccd _086_ sky130_fd_sc_hd__clkinv_2
X_576_ net146 vssd vssd vccd vccd _087_ sky130_fd_sc_hd__inv_2
X_577_ net147 vssd vssd vccd vccd _088_ sky130_fd_sc_hd__inv_2
X_578_ net148 vssd vssd vccd vccd _089_ sky130_fd_sc_hd__inv_4
X_579_ net149 vssd vssd vccd vccd _090_ sky130_fd_sc_hd__clkinv_2
X_580_ net150 vssd vssd vccd vccd _091_ sky130_fd_sc_hd__inv_2
X_581_ net151 vssd vssd vccd vccd _092_ sky130_fd_sc_hd__clkinv_2
X_582_ net152 vssd vssd vccd vccd _093_ sky130_fd_sc_hd__inv_2
X_583_ net153 vssd vssd vccd vccd _094_ sky130_fd_sc_hd__inv_2
X_584_ net155 vssd vssd vccd vccd _096_ sky130_fd_sc_hd__clkinv_2
X_585_ net156 vssd vssd vccd vccd _097_ sky130_fd_sc_hd__inv_2
X_586_ net157 vssd vssd vccd vccd _098_ sky130_fd_sc_hd__inv_2
X_587_ net158 vssd vssd vccd vccd _099_ sky130_fd_sc_hd__clkinv_2
X_588_ net159 vssd vssd vccd vccd _100_ sky130_fd_sc_hd__clkinv_2
X_589_ net160 vssd vssd vccd vccd _101_ sky130_fd_sc_hd__inv_2
X_590_ net161 vssd vssd vccd vccd _102_ sky130_fd_sc_hd__inv_2
X_591_ net162 vssd vssd vccd vccd _103_ sky130_fd_sc_hd__clkinv_2
X_592_ net388 vssd vssd vccd vccd _201_ sky130_fd_sc_hd__clkinv_2
X_593_ net427 vssd vssd vccd vccd _240_ sky130_fd_sc_hd__clkinv_4
X_594_ net438 vssd vssd vccd vccd _251_ sky130_fd_sc_hd__clkinv_4
X_595_ net449 vssd vssd vccd vccd _262_ sky130_fd_sc_hd__inv_2
X_596_ net460 vssd vssd vccd vccd _273_ sky130_fd_sc_hd__clkinv_4
X_597_ net471 vssd vssd vccd vccd _284_ sky130_fd_sc_hd__clkinv_4
X_598_ net482 vssd vssd vccd vccd _295_ sky130_fd_sc_hd__clkinv_2
X_599_ net493 vssd vssd vccd vccd _306_ sky130_fd_sc_hd__clkinv_4
X_600_ net504 vssd vssd vccd vccd _317_ sky130_fd_sc_hd__clkinv_4
X_601_ net515 vssd vssd vccd vccd _328_ sky130_fd_sc_hd__inv_2
X_602_ net399 vssd vssd vccd vccd _212_ sky130_fd_sc_hd__clkinv_2
X_603_ net410 vssd vssd vccd vccd _223_ sky130_fd_sc_hd__inv_2
X_604_ net419 vssd vssd vccd vccd _232_ sky130_fd_sc_hd__clkinv_4
X_605_ net420 vssd vssd vccd vccd _233_ sky130_fd_sc_hd__clkinv_2
X_606_ net421 vssd vssd vccd vccd _234_ sky130_fd_sc_hd__clkinv_4
X_607_ net422 vssd vssd vccd vccd _235_ sky130_fd_sc_hd__clkinv_4
X_608_ net423 vssd vssd vccd vccd _236_ sky130_fd_sc_hd__inv_2
X_609_ net424 vssd vssd vccd vccd _237_ sky130_fd_sc_hd__inv_2
X_610_ net425 vssd vssd vccd vccd _238_ sky130_fd_sc_hd__clkinv_2
X_611_ net426 vssd vssd vccd vccd _239_ sky130_fd_sc_hd__clkinv_2
X_612_ net428 vssd vssd vccd vccd _241_ sky130_fd_sc_hd__clkinv_4
X_613_ net429 vssd vssd vccd vccd _242_ sky130_fd_sc_hd__clkinv_2
X_614_ net430 vssd vssd vccd vccd _243_ sky130_fd_sc_hd__inv_2
X_615_ net431 vssd vssd vccd vccd _244_ sky130_fd_sc_hd__inv_2
X_616_ net432 vssd vssd vccd vccd _245_ sky130_fd_sc_hd__clkinv_2
X_617_ net433 vssd vssd vccd vccd _246_ sky130_fd_sc_hd__clkinv_2
X_618_ net434 vssd vssd vccd vccd _247_ sky130_fd_sc_hd__inv_2
X_619_ net435 vssd vssd vccd vccd _248_ sky130_fd_sc_hd__clkinv_2
X_620_ net436 vssd vssd vccd vccd _249_ sky130_fd_sc_hd__clkinv_2
X_621_ net437 vssd vssd vccd vccd _250_ sky130_fd_sc_hd__inv_2
X_622_ net439 vssd vssd vccd vccd _252_ sky130_fd_sc_hd__clkinv_4
X_623_ net440 vssd vssd vccd vccd _253_ sky130_fd_sc_hd__clkinv_4
X_624_ net441 vssd vssd vccd vccd _254_ sky130_fd_sc_hd__clkinv_4
X_625_ net442 vssd vssd vccd vccd _255_ sky130_fd_sc_hd__clkinv_4
X_626_ net443 vssd vssd vccd vccd _256_ sky130_fd_sc_hd__inv_2
X_627_ net444 vssd vssd vccd vccd _257_ sky130_fd_sc_hd__clkinv_4
X_628_ net445 vssd vssd vccd vccd _258_ sky130_fd_sc_hd__inv_2
X_629_ net446 vssd vssd vccd vccd _259_ sky130_fd_sc_hd__clkinv_4
X_630_ net447 vssd vssd vccd vccd _260_ sky130_fd_sc_hd__clkinv_4
X_631_ net448 vssd vssd vccd vccd _261_ sky130_fd_sc_hd__inv_2
X_632_ net450 vssd vssd vccd vccd _263_ sky130_fd_sc_hd__clkinv_2
X_633_ net451 vssd vssd vccd vccd _264_ sky130_fd_sc_hd__inv_2
X_634_ net452 vssd vssd vccd vccd _265_ sky130_fd_sc_hd__inv_2
X_635_ net453 vssd vssd vccd vccd _266_ sky130_fd_sc_hd__clkinv_2
X_636_ net454 vssd vssd vccd vccd _267_ sky130_fd_sc_hd__clkinv_4
X_637_ net455 vssd vssd vccd vccd _268_ sky130_fd_sc_hd__inv_2
X_638_ net456 vssd vssd vccd vccd _269_ sky130_fd_sc_hd__clkinv_2
X_639_ net457 vssd vssd vccd vccd _270_ sky130_fd_sc_hd__clkinv_2
X_640_ net458 vssd vssd vccd vccd _271_ sky130_fd_sc_hd__clkinv_4
X_641_ net459 vssd vssd vccd vccd _272_ sky130_fd_sc_hd__clkinv_2
X_642_ net461 vssd vssd vccd vccd _274_ sky130_fd_sc_hd__inv_2
X_643_ net462 vssd vssd vccd vccd _275_ sky130_fd_sc_hd__clkinv_4
X_644_ net463 vssd vssd vccd vccd _276_ sky130_fd_sc_hd__inv_2
X_645_ net464 vssd vssd vccd vccd _277_ sky130_fd_sc_hd__clkinv_2
X_646_ net465 vssd vssd vccd vccd _278_ sky130_fd_sc_hd__inv_2
X_647_ net466 vssd vssd vccd vccd _279_ sky130_fd_sc_hd__clkinv_2
X_648_ net467 vssd vssd vccd vccd _280_ sky130_fd_sc_hd__clkinv_2
X_649_ net468 vssd vssd vccd vccd _281_ sky130_fd_sc_hd__inv_2
X_650_ net469 vssd vssd vccd vccd _282_ sky130_fd_sc_hd__clkinv_2
X_651_ net470 vssd vssd vccd vccd _283_ sky130_fd_sc_hd__inv_2
X_652_ net472 vssd vssd vccd vccd _285_ sky130_fd_sc_hd__inv_2
X_653_ net473 vssd vssd vccd vccd _286_ sky130_fd_sc_hd__inv_2
X_654_ net474 vssd vssd vccd vccd _287_ sky130_fd_sc_hd__clkinv_2
X_655_ net475 vssd vssd vccd vccd _288_ sky130_fd_sc_hd__inv_2
X_656_ net476 vssd vssd vccd vccd _289_ sky130_fd_sc_hd__inv_2
X_657_ net477 vssd vssd vccd vccd _290_ sky130_fd_sc_hd__inv_2
Xinput1 caravel_clk vssd vssd vccd vccd net1 sky130_fd_sc_hd__clkbuf_1
Xinput10 la_data_out_core[105] vssd vssd vccd vccd net10 sky130_fd_sc_hd__buf_4
Xinput100 la_data_out_core[71] vssd vssd vccd vccd net100 sky130_fd_sc_hd__buf_4
Xinput101 la_data_out_core[72] vssd vssd vccd vccd net101 sky130_fd_sc_hd__buf_4
Xinput102 la_data_out_core[73] vssd vssd vccd vccd net102 sky130_fd_sc_hd__buf_4
Xinput103 la_data_out_core[74] vssd vssd vccd vccd net103 sky130_fd_sc_hd__buf_4
Xinput104 la_data_out_core[75] vssd vssd vccd vccd net104 sky130_fd_sc_hd__buf_4
Xinput105 la_data_out_core[76] vssd vssd vccd vccd net105 sky130_fd_sc_hd__buf_4
Xinput106 la_data_out_core[77] vssd vssd vccd vccd net106 sky130_fd_sc_hd__buf_4
Xinput107 la_data_out_core[78] vssd vssd vccd vccd net107 sky130_fd_sc_hd__buf_4
Xinput108 la_data_out_core[79] vssd vssd vccd vccd net108 sky130_fd_sc_hd__buf_4
Xinput109 la_data_out_core[7] vssd vssd vccd vccd net109 sky130_fd_sc_hd__buf_2
Xinput11 la_data_out_core[106] vssd vssd vccd vccd net11 sky130_fd_sc_hd__buf_4
Xinput110 la_data_out_core[80] vssd vssd vccd vccd net110 sky130_fd_sc_hd__buf_4
Xinput111 la_data_out_core[81] vssd vssd vccd vccd net111 sky130_fd_sc_hd__buf_4
Xinput112 la_data_out_core[82] vssd vssd vccd vccd net112 sky130_fd_sc_hd__buf_4
Xinput113 la_data_out_core[83] vssd vssd vccd vccd net113 sky130_fd_sc_hd__buf_4
Xinput114 la_data_out_core[84] vssd vssd vccd vccd net114 sky130_fd_sc_hd__buf_4
Xinput115 la_data_out_core[85] vssd vssd vccd vccd net115 sky130_fd_sc_hd__buf_4
Xinput116 la_data_out_core[86] vssd vssd vccd vccd net116 sky130_fd_sc_hd__clkbuf_4
Xinput117 la_data_out_core[87] vssd vssd vccd vccd net117 sky130_fd_sc_hd__buf_4
Xinput118 la_data_out_core[88] vssd vssd vccd vccd net118 sky130_fd_sc_hd__buf_4
Xinput119 la_data_out_core[89] vssd vssd vccd vccd net119 sky130_fd_sc_hd__buf_4
Xinput12 la_data_out_core[107] vssd vssd vccd vccd net12 sky130_fd_sc_hd__clkbuf_4
Xinput120 la_data_out_core[8] vssd vssd vccd vccd net120 sky130_fd_sc_hd__buf_2
Xinput121 la_data_out_core[90] vssd vssd vccd vccd net121 sky130_fd_sc_hd__buf_4
Xinput122 la_data_out_core[91] vssd vssd vccd vccd net122 sky130_fd_sc_hd__buf_4
Xinput123 la_data_out_core[92] vssd vssd vccd vccd net123 sky130_fd_sc_hd__buf_4
Xinput124 la_data_out_core[93] vssd vssd vccd vccd net124 sky130_fd_sc_hd__buf_4
Xinput125 la_data_out_core[94] vssd vssd vccd vccd net125 sky130_fd_sc_hd__clkbuf_4
Xinput126 la_data_out_core[95] vssd vssd vccd vccd net126 sky130_fd_sc_hd__clkbuf_4
Xinput127 la_data_out_core[96] vssd vssd vccd vccd net127 sky130_fd_sc_hd__clkbuf_4
Xinput128 la_data_out_core[97] vssd vssd vccd vccd net128 sky130_fd_sc_hd__buf_4
Xinput129 la_data_out_core[98] vssd vssd vccd vccd net129 sky130_fd_sc_hd__clkbuf_4
Xinput13 la_data_out_core[108] vssd vssd vccd vccd net13 sky130_fd_sc_hd__buf_4
Xinput130 la_data_out_core[99] vssd vssd vccd vccd net130 sky130_fd_sc_hd__buf_4
Xinput131 la_data_out_core[9] vssd vssd vccd vccd net131 sky130_fd_sc_hd__buf_2
Xinput132 la_data_out_mprj[0] vssd vssd vccd vccd net132 sky130_fd_sc_hd__clkbuf_2
Xinput133 la_data_out_mprj[100] vssd vssd vccd vccd net133 sky130_fd_sc_hd__clkbuf_4
Xinput134 la_data_out_mprj[101] vssd vssd vccd vccd net134 sky130_fd_sc_hd__clkbuf_4
Xinput135 la_data_out_mprj[102] vssd vssd vccd vccd net135 sky130_fd_sc_hd__clkbuf_2
Xinput136 la_data_out_mprj[103] vssd vssd vccd vccd net136 sky130_fd_sc_hd__clkbuf_2
Xinput137 la_data_out_mprj[104] vssd vssd vccd vccd net137 sky130_fd_sc_hd__clkbuf_2
Xinput138 la_data_out_mprj[105] vssd vssd vccd vccd net138 sky130_fd_sc_hd__clkbuf_1
Xinput139 la_data_out_mprj[106] vssd vssd vccd vccd net139 sky130_fd_sc_hd__buf_2
Xinput14 la_data_out_core[109] vssd vssd vccd vccd net14 sky130_fd_sc_hd__clkbuf_4
Xinput140 la_data_out_mprj[107] vssd vssd vccd vccd net140 sky130_fd_sc_hd__clkbuf_4
Xinput141 la_data_out_mprj[108] vssd vssd vccd vccd net141 sky130_fd_sc_hd__clkbuf_4
Xinput142 la_data_out_mprj[109] vssd vssd vccd vccd net142 sky130_fd_sc_hd__clkbuf_4
Xinput143 la_data_out_mprj[10] vssd vssd vccd vccd net143 sky130_fd_sc_hd__clkbuf_2
Xinput144 la_data_out_mprj[110] vssd vssd vccd vccd net144 sky130_fd_sc_hd__clkbuf_4
Xinput145 la_data_out_mprj[111] vssd vssd vccd vccd net145 sky130_fd_sc_hd__buf_4
Xinput146 la_data_out_mprj[112] vssd vssd vccd vccd net146 sky130_fd_sc_hd__clkbuf_4
Xinput147 la_data_out_mprj[113] vssd vssd vccd vccd net147 sky130_fd_sc_hd__clkbuf_4
Xinput148 la_data_out_mprj[114] vssd vssd vccd vccd net148 sky130_fd_sc_hd__clkbuf_1
Xinput149 la_data_out_mprj[115] vssd vssd vccd vccd net149 sky130_fd_sc_hd__clkbuf_4
Xinput15 la_data_out_core[10] vssd vssd vccd vccd net15 sky130_fd_sc_hd__clkbuf_4
Xinput150 la_data_out_mprj[116] vssd vssd vccd vccd net150 sky130_fd_sc_hd__clkbuf_2
Xinput151 la_data_out_mprj[117] vssd vssd vccd vccd net151 sky130_fd_sc_hd__clkbuf_4
Xinput152 la_data_out_mprj[118] vssd vssd vccd vccd net152 sky130_fd_sc_hd__clkbuf_2
Xinput153 la_data_out_mprj[119] vssd vssd vccd vccd net153 sky130_fd_sc_hd__clkbuf_2
Xinput154 la_data_out_mprj[11] vssd vssd vccd vccd net154 sky130_fd_sc_hd__clkbuf_2
Xinput155 la_data_out_mprj[120] vssd vssd vccd vccd net155 sky130_fd_sc_hd__buf_2
Xinput156 la_data_out_mprj[121] vssd vssd vccd vccd net156 sky130_fd_sc_hd__clkbuf_2
Xinput157 la_data_out_mprj[122] vssd vssd vccd vccd net157 sky130_fd_sc_hd__clkbuf_4
Xinput158 la_data_out_mprj[123] vssd vssd vccd vccd net158 sky130_fd_sc_hd__buf_2
Xinput159 la_data_out_mprj[124] vssd vssd vccd vccd net159 sky130_fd_sc_hd__clkbuf_4
Xinput16 la_data_out_core[110] vssd vssd vccd vccd net16 sky130_fd_sc_hd__clkbuf_4
Xinput160 la_data_out_mprj[125] vssd vssd vccd vccd net160 sky130_fd_sc_hd__clkbuf_2
Xinput161 la_data_out_mprj[126] vssd vssd vccd vccd net161 sky130_fd_sc_hd__clkbuf_2
Xinput162 la_data_out_mprj[127] vssd vssd vccd vccd net162 sky130_fd_sc_hd__buf_2
Xinput163 la_data_out_mprj[12] vssd vssd vccd vccd net163 sky130_fd_sc_hd__clkbuf_2
Xinput164 la_data_out_mprj[13] vssd vssd vccd vccd net164 sky130_fd_sc_hd__clkbuf_2
Xinput165 la_data_out_mprj[14] vssd vssd vccd vccd net165 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput166 la_data_out_mprj[15] vssd vssd vccd vccd net166 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput167 la_data_out_mprj[16] vssd vssd vccd vccd net167 sky130_fd_sc_hd__clkbuf_2
Xinput168 la_data_out_mprj[17] vssd vssd vccd vccd net168 sky130_fd_sc_hd__clkbuf_2
Xinput169 la_data_out_mprj[18] vssd vssd vccd vccd net169 sky130_fd_sc_hd__clkbuf_2
Xinput17 la_data_out_core[111] vssd vssd vccd vccd net17 sky130_fd_sc_hd__clkbuf_4
Xinput170 la_data_out_mprj[19] vssd vssd vccd vccd net170 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput171 la_data_out_mprj[1] vssd vssd vccd vccd net171 sky130_fd_sc_hd__clkbuf_2
Xinput172 la_data_out_mprj[20] vssd vssd vccd vccd net172 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput173 la_data_out_mprj[21] vssd vssd vccd vccd net173 sky130_fd_sc_hd__clkbuf_2
Xinput174 la_data_out_mprj[22] vssd vssd vccd vccd net174 sky130_fd_sc_hd__clkbuf_2
Xinput175 la_data_out_mprj[23] vssd vssd vccd vccd net175 sky130_fd_sc_hd__clkbuf_2
Xinput176 la_data_out_mprj[24] vssd vssd vccd vccd net176 sky130_fd_sc_hd__clkbuf_2
Xinput177 la_data_out_mprj[25] vssd vssd vccd vccd net177 sky130_fd_sc_hd__clkbuf_2
Xinput178 la_data_out_mprj[26] vssd vssd vccd vccd net178 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput179 la_data_out_mprj[27] vssd vssd vccd vccd net179 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput18 la_data_out_core[112] vssd vssd vccd vccd net18 sky130_fd_sc_hd__clkbuf_4
Xinput180 la_data_out_mprj[28] vssd vssd vccd vccd net180 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput181 la_data_out_mprj[29] vssd vssd vccd vccd net181 sky130_fd_sc_hd__clkbuf_2
Xinput182 la_data_out_mprj[2] vssd vssd vccd vccd net182 sky130_fd_sc_hd__clkbuf_2
Xinput183 la_data_out_mprj[30] vssd vssd vccd vccd net183 sky130_fd_sc_hd__clkbuf_2
Xinput184 la_data_out_mprj[31] vssd vssd vccd vccd net184 sky130_fd_sc_hd__clkbuf_2
Xinput185 la_data_out_mprj[32] vssd vssd vccd vccd net185 sky130_fd_sc_hd__clkbuf_2
Xinput186 la_data_out_mprj[33] vssd vssd vccd vccd net186 sky130_fd_sc_hd__clkbuf_2
Xinput187 la_data_out_mprj[34] vssd vssd vccd vccd net187 sky130_fd_sc_hd__clkbuf_2
Xinput188 la_data_out_mprj[35] vssd vssd vccd vccd net188 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput189 la_data_out_mprj[36] vssd vssd vccd vccd net189 sky130_fd_sc_hd__clkbuf_1
Xinput19 la_data_out_core[113] vssd vssd vccd vccd net19 sky130_fd_sc_hd__clkbuf_4
Xinput190 la_data_out_mprj[37] vssd vssd vccd vccd net190 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput191 la_data_out_mprj[38] vssd vssd vccd vccd net191 sky130_fd_sc_hd__clkbuf_1
Xinput192 la_data_out_mprj[39] vssd vssd vccd vccd net192 sky130_fd_sc_hd__clkbuf_1
Xinput193 la_data_out_mprj[3] vssd vssd vccd vccd net193 sky130_fd_sc_hd__clkbuf_2
Xinput194 la_data_out_mprj[40] vssd vssd vccd vccd net194 sky130_fd_sc_hd__clkbuf_2
Xinput195 la_data_out_mprj[41] vssd vssd vccd vccd net195 sky130_fd_sc_hd__clkbuf_2
Xinput196 la_data_out_mprj[42] vssd vssd vccd vccd net196 sky130_fd_sc_hd__clkbuf_2
Xinput197 la_data_out_mprj[43] vssd vssd vccd vccd net197 sky130_fd_sc_hd__clkbuf_2
Xinput198 la_data_out_mprj[44] vssd vssd vccd vccd net198 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput199 la_data_out_mprj[45] vssd vssd vccd vccd net199 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput2 caravel_clk2 vssd vssd vccd vccd net2 sky130_fd_sc_hd__clkbuf_1
Xinput20 la_data_out_core[114] vssd vssd vccd vccd net20 sky130_fd_sc_hd__clkbuf_4
Xinput200 la_data_out_mprj[46] vssd vssd vccd vccd net200 sky130_fd_sc_hd__clkbuf_2
Xinput201 la_data_out_mprj[47] vssd vssd vccd vccd net201 sky130_fd_sc_hd__clkbuf_2
Xinput202 la_data_out_mprj[48] vssd vssd vccd vccd net202 sky130_fd_sc_hd__clkbuf_2
Xinput203 la_data_out_mprj[49] vssd vssd vccd vccd net203 sky130_fd_sc_hd__clkbuf_2
Xinput204 la_data_out_mprj[4] vssd vssd vccd vccd net204 sky130_fd_sc_hd__clkbuf_2
Xinput205 la_data_out_mprj[50] vssd vssd vccd vccd net205 sky130_fd_sc_hd__clkbuf_2
Xinput206 la_data_out_mprj[51] vssd vssd vccd vccd net206 sky130_fd_sc_hd__clkbuf_2
Xinput207 la_data_out_mprj[52] vssd vssd vccd vccd net207 sky130_fd_sc_hd__clkbuf_2
Xinput208 la_data_out_mprj[53] vssd vssd vccd vccd net208 sky130_fd_sc_hd__clkbuf_2
Xinput209 la_data_out_mprj[54] vssd vssd vccd vccd net209 sky130_fd_sc_hd__clkbuf_2
Xinput21 la_data_out_core[115] vssd vssd vccd vccd net21 sky130_fd_sc_hd__clkbuf_4
Xinput210 la_data_out_mprj[55] vssd vssd vccd vccd net210 sky130_fd_sc_hd__clkbuf_2
Xinput211 la_data_out_mprj[56] vssd vssd vccd vccd net211 sky130_fd_sc_hd__clkbuf_2
Xinput212 la_data_out_mprj[57] vssd vssd vccd vccd net212 sky130_fd_sc_hd__clkbuf_2
Xinput213 la_data_out_mprj[58] vssd vssd vccd vccd net213 sky130_fd_sc_hd__clkbuf_2
Xinput214 la_data_out_mprj[59] vssd vssd vccd vccd net214 sky130_fd_sc_hd__clkbuf_2
Xinput215 la_data_out_mprj[5] vssd vssd vccd vccd net215 sky130_fd_sc_hd__clkbuf_2
Xinput216 la_data_out_mprj[60] vssd vssd vccd vccd net216 sky130_fd_sc_hd__clkbuf_2
Xinput217 la_data_out_mprj[61] vssd vssd vccd vccd net217 sky130_fd_sc_hd__clkbuf_2
Xinput218 la_data_out_mprj[62] vssd vssd vccd vccd net218 sky130_fd_sc_hd__clkbuf_2
Xinput219 la_data_out_mprj[63] vssd vssd vccd vccd net219 sky130_fd_sc_hd__clkbuf_2
Xinput22 la_data_out_core[116] vssd vssd vccd vccd net22 sky130_fd_sc_hd__clkbuf_4
Xinput220 la_data_out_mprj[64] vssd vssd vccd vccd net220 sky130_fd_sc_hd__clkbuf_2
Xinput221 la_data_out_mprj[65] vssd vssd vccd vccd net221 sky130_fd_sc_hd__clkbuf_2
Xinput222 la_data_out_mprj[66] vssd vssd vccd vccd net222 sky130_fd_sc_hd__clkbuf_2
Xinput223 la_data_out_mprj[67] vssd vssd vccd vccd net223 sky130_fd_sc_hd__clkbuf_2
Xinput224 la_data_out_mprj[68] vssd vssd vccd vccd net224 sky130_fd_sc_hd__clkbuf_2
Xinput225 la_data_out_mprj[69] vssd vssd vccd vccd net225 sky130_fd_sc_hd__clkbuf_2
Xinput226 la_data_out_mprj[6] vssd vssd vccd vccd net226 sky130_fd_sc_hd__clkbuf_2
Xinput227 la_data_out_mprj[70] vssd vssd vccd vccd net227 sky130_fd_sc_hd__buf_2
Xinput228 la_data_out_mprj[71] vssd vssd vccd vccd net228 sky130_fd_sc_hd__clkbuf_2
Xinput229 la_data_out_mprj[72] vssd vssd vccd vccd net229 sky130_fd_sc_hd__clkbuf_2
Xinput23 la_data_out_core[117] vssd vssd vccd vccd net23 sky130_fd_sc_hd__clkbuf_4
Xinput230 la_data_out_mprj[73] vssd vssd vccd vccd net230 sky130_fd_sc_hd__buf_2
Xinput231 la_data_out_mprj[74] vssd vssd vccd vccd net231 sky130_fd_sc_hd__buf_2
Xinput232 la_data_out_mprj[75] vssd vssd vccd vccd net232 sky130_fd_sc_hd__buf_2
Xinput233 la_data_out_mprj[76] vssd vssd vccd vccd net233 sky130_fd_sc_hd__clkbuf_4
Xinput234 la_data_out_mprj[77] vssd vssd vccd vccd net234 sky130_fd_sc_hd__clkbuf_2
Xinput235 la_data_out_mprj[78] vssd vssd vccd vccd net235 sky130_fd_sc_hd__buf_2
Xinput236 la_data_out_mprj[79] vssd vssd vccd vccd net236 sky130_fd_sc_hd__clkbuf_4
Xinput237 la_data_out_mprj[7] vssd vssd vccd vccd net237 sky130_fd_sc_hd__clkbuf_2
Xinput238 la_data_out_mprj[80] vssd vssd vccd vccd net238 sky130_fd_sc_hd__clkbuf_4
Xinput239 la_data_out_mprj[81] vssd vssd vccd vccd net239 sky130_fd_sc_hd__clkbuf_4
Xinput24 la_data_out_core[118] vssd vssd vccd vccd net24 sky130_fd_sc_hd__clkbuf_4
Xinput240 la_data_out_mprj[82] vssd vssd vccd vccd net240 sky130_fd_sc_hd__buf_2
Xinput241 la_data_out_mprj[83] vssd vssd vccd vccd net241 sky130_fd_sc_hd__clkbuf_4
Xinput242 la_data_out_mprj[84] vssd vssd vccd vccd net242 sky130_fd_sc_hd__buf_4
Xinput243 la_data_out_mprj[85] vssd vssd vccd vccd net243 sky130_fd_sc_hd__clkbuf_4
Xinput244 la_data_out_mprj[86] vssd vssd vccd vccd net244 sky130_fd_sc_hd__clkbuf_4
Xinput245 la_data_out_mprj[87] vssd vssd vccd vccd net245 sky130_fd_sc_hd__clkbuf_2
Xinput246 la_data_out_mprj[88] vssd vssd vccd vccd net246 sky130_fd_sc_hd__buf_2
Xinput247 la_data_out_mprj[89] vssd vssd vccd vccd net247 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput248 la_data_out_mprj[8] vssd vssd vccd vccd net248 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput249 la_data_out_mprj[90] vssd vssd vccd vccd net249 sky130_fd_sc_hd__clkbuf_1
Xinput25 la_data_out_core[119] vssd vssd vccd vccd net25 sky130_fd_sc_hd__clkbuf_4
Xinput250 la_data_out_mprj[91] vssd vssd vccd vccd net250 sky130_fd_sc_hd__clkbuf_2
Xinput251 la_data_out_mprj[92] vssd vssd vccd vccd net251 sky130_fd_sc_hd__clkbuf_2
Xinput252 la_data_out_mprj[93] vssd vssd vccd vccd net252 sky130_fd_sc_hd__clkbuf_2
Xinput253 la_data_out_mprj[94] vssd vssd vccd vccd net253 sky130_fd_sc_hd__buf_2
Xinput254 la_data_out_mprj[95] vssd vssd vccd vccd net254 sky130_fd_sc_hd__buf_2
Xinput255 la_data_out_mprj[96] vssd vssd vccd vccd net255 sky130_fd_sc_hd__clkbuf_2
Xinput256 la_data_out_mprj[97] vssd vssd vccd vccd net256 sky130_fd_sc_hd__buf_2
Xinput257 la_data_out_mprj[98] vssd vssd vccd vccd net257 sky130_fd_sc_hd__buf_2
Xinput258 la_data_out_mprj[99] vssd vssd vccd vccd net258 sky130_fd_sc_hd__clkbuf_2
Xinput259 la_data_out_mprj[9] vssd vssd vccd vccd net259 sky130_fd_sc_hd__clkbuf_2
Xinput26 la_data_out_core[11] vssd vssd vccd vccd net26 sky130_fd_sc_hd__clkbuf_2
Xinput260 la_iena_mprj[0] vssd vssd vccd vccd net260 sky130_fd_sc_hd__clkbuf_1
Xinput261 la_iena_mprj[100] vssd vssd vccd vccd net261 sky130_fd_sc_hd__clkbuf_1
Xinput262 la_iena_mprj[101] vssd vssd vccd vccd net262 sky130_fd_sc_hd__clkbuf_1
Xinput263 la_iena_mprj[102] vssd vssd vccd vccd net263 sky130_fd_sc_hd__clkbuf_1
Xinput264 la_iena_mprj[103] vssd vssd vccd vccd net264 sky130_fd_sc_hd__clkbuf_1
Xinput265 la_iena_mprj[104] vssd vssd vccd vccd net265 sky130_fd_sc_hd__clkbuf_1
Xinput266 la_iena_mprj[105] vssd vssd vccd vccd net266 sky130_fd_sc_hd__clkbuf_1
Xinput267 la_iena_mprj[106] vssd vssd vccd vccd net267 sky130_fd_sc_hd__clkbuf_1
Xinput268 la_iena_mprj[107] vssd vssd vccd vccd net268 sky130_fd_sc_hd__clkbuf_1
Xinput269 la_iena_mprj[108] vssd vssd vccd vccd net269 sky130_fd_sc_hd__clkbuf_1
Xinput27 la_data_out_core[120] vssd vssd vccd vccd net27 sky130_fd_sc_hd__clkbuf_4
Xinput270 la_iena_mprj[109] vssd vssd vccd vccd net270 sky130_fd_sc_hd__clkbuf_1
Xinput271 la_iena_mprj[10] vssd vssd vccd vccd net271 sky130_fd_sc_hd__clkbuf_2
Xinput272 la_iena_mprj[110] vssd vssd vccd vccd net272 sky130_fd_sc_hd__clkbuf_1
Xinput273 la_iena_mprj[111] vssd vssd vccd vccd net273 sky130_fd_sc_hd__clkbuf_1
Xinput274 la_iena_mprj[112] vssd vssd vccd vccd net274 sky130_fd_sc_hd__clkbuf_1
Xinput275 la_iena_mprj[113] vssd vssd vccd vccd net275 sky130_fd_sc_hd__clkbuf_1
Xinput276 la_iena_mprj[114] vssd vssd vccd vccd net276 sky130_fd_sc_hd__clkbuf_1
Xinput277 la_iena_mprj[115] vssd vssd vccd vccd net277 sky130_fd_sc_hd__clkbuf_1
Xinput278 la_iena_mprj[116] vssd vssd vccd vccd net278 sky130_fd_sc_hd__clkbuf_1
Xinput279 la_iena_mprj[117] vssd vssd vccd vccd net279 sky130_fd_sc_hd__clkbuf_1
Xinput28 la_data_out_core[121] vssd vssd vccd vccd net28 sky130_fd_sc_hd__clkbuf_4
Xinput280 la_iena_mprj[118] vssd vssd vccd vccd net280 sky130_fd_sc_hd__clkbuf_1
Xinput281 la_iena_mprj[119] vssd vssd vccd vccd net281 sky130_fd_sc_hd__clkbuf_1
Xinput282 la_iena_mprj[11] vssd vssd vccd vccd net282 sky130_fd_sc_hd__clkbuf_4
Xinput283 la_iena_mprj[120] vssd vssd vccd vccd net283 sky130_fd_sc_hd__clkbuf_1
Xinput284 la_iena_mprj[121] vssd vssd vccd vccd net284 sky130_fd_sc_hd__clkbuf_1
Xinput285 la_iena_mprj[122] vssd vssd vccd vccd net285 sky130_fd_sc_hd__clkbuf_1
Xinput286 la_iena_mprj[123] vssd vssd vccd vccd net286 sky130_fd_sc_hd__clkbuf_1
Xinput287 la_iena_mprj[124] vssd vssd vccd vccd net287 sky130_fd_sc_hd__clkbuf_1
Xinput288 la_iena_mprj[125] vssd vssd vccd vccd net288 sky130_fd_sc_hd__clkbuf_1
Xinput289 la_iena_mprj[126] vssd vssd vccd vccd net289 sky130_fd_sc_hd__clkbuf_1
Xinput29 la_data_out_core[122] vssd vssd vccd vccd net29 sky130_fd_sc_hd__clkbuf_4
Xinput290 la_iena_mprj[127] vssd vssd vccd vccd net290 sky130_fd_sc_hd__clkbuf_1
Xinput291 la_iena_mprj[12] vssd vssd vccd vccd net291 sky130_fd_sc_hd__clkbuf_4
Xinput292 la_iena_mprj[13] vssd vssd vccd vccd net292 sky130_fd_sc_hd__clkbuf_1
Xinput293 la_iena_mprj[14] vssd vssd vccd vccd net293 sky130_fd_sc_hd__clkbuf_1
Xinput294 la_iena_mprj[15] vssd vssd vccd vccd net294 sky130_fd_sc_hd__clkbuf_1
Xinput295 la_iena_mprj[16] vssd vssd vccd vccd net295 sky130_fd_sc_hd__clkbuf_1
Xinput296 la_iena_mprj[17] vssd vssd vccd vccd net296 sky130_fd_sc_hd__clkbuf_1
Xinput297 la_iena_mprj[18] vssd vssd vccd vccd net297 sky130_fd_sc_hd__clkbuf_1
Xinput298 la_iena_mprj[19] vssd vssd vccd vccd net298 sky130_fd_sc_hd__clkbuf_1
Xinput299 la_iena_mprj[1] vssd vssd vccd vccd net299 sky130_fd_sc_hd__clkbuf_1
Xinput3 caravel_rstn vssd vssd vccd vccd net3 sky130_fd_sc_hd__clkbuf_2
Xinput30 la_data_out_core[123] vssd vssd vccd vccd net30 sky130_fd_sc_hd__clkbuf_4
Xinput300 la_iena_mprj[20] vssd vssd vccd vccd net300 sky130_fd_sc_hd__clkbuf_1
Xinput301 la_iena_mprj[21] vssd vssd vccd vccd net301 sky130_fd_sc_hd__clkbuf_1
Xinput302 la_iena_mprj[22] vssd vssd vccd vccd net302 sky130_fd_sc_hd__clkbuf_1
Xinput303 la_iena_mprj[23] vssd vssd vccd vccd net303 sky130_fd_sc_hd__clkbuf_1
Xinput304 la_iena_mprj[24] vssd vssd vccd vccd net304 sky130_fd_sc_hd__clkbuf_1
Xinput305 la_iena_mprj[25] vssd vssd vccd vccd net305 sky130_fd_sc_hd__clkbuf_1
Xinput306 la_iena_mprj[26] vssd vssd vccd vccd net306 sky130_fd_sc_hd__clkbuf_1
Xinput307 la_iena_mprj[27] vssd vssd vccd vccd net307 sky130_fd_sc_hd__clkbuf_1
Xinput308 la_iena_mprj[28] vssd vssd vccd vccd net308 sky130_fd_sc_hd__clkbuf_1
Xinput309 la_iena_mprj[29] vssd vssd vccd vccd net309 sky130_fd_sc_hd__clkbuf_1
Xinput31 la_data_out_core[124] vssd vssd vccd vccd net31 sky130_fd_sc_hd__clkbuf_4
Xinput310 la_iena_mprj[2] vssd vssd vccd vccd net310 sky130_fd_sc_hd__clkbuf_1
Xinput311 la_iena_mprj[30] vssd vssd vccd vccd net311 sky130_fd_sc_hd__clkbuf_1
Xinput312 la_iena_mprj[31] vssd vssd vccd vccd net312 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput313 la_iena_mprj[32] vssd vssd vccd vccd net313 sky130_fd_sc_hd__clkbuf_1
Xinput314 la_iena_mprj[33] vssd vssd vccd vccd net314 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput315 la_iena_mprj[34] vssd vssd vccd vccd net315 sky130_fd_sc_hd__clkbuf_1
Xinput316 la_iena_mprj[35] vssd vssd vccd vccd net316 sky130_fd_sc_hd__clkbuf_1
Xinput317 la_iena_mprj[36] vssd vssd vccd vccd net317 sky130_fd_sc_hd__clkbuf_1
Xinput318 la_iena_mprj[37] vssd vssd vccd vccd net318 sky130_fd_sc_hd__clkbuf_1
Xinput319 la_iena_mprj[38] vssd vssd vccd vccd net319 sky130_fd_sc_hd__clkbuf_1
Xinput32 la_data_out_core[125] vssd vssd vccd vccd net32 sky130_fd_sc_hd__clkbuf_4
Xinput320 la_iena_mprj[39] vssd vssd vccd vccd net320 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput321 la_iena_mprj[3] vssd vssd vccd vccd net321 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput322 la_iena_mprj[40] vssd vssd vccd vccd net322 sky130_fd_sc_hd__clkbuf_1
Xinput323 la_iena_mprj[41] vssd vssd vccd vccd net323 sky130_fd_sc_hd__clkbuf_1
Xinput324 la_iena_mprj[42] vssd vssd vccd vccd net324 sky130_fd_sc_hd__clkbuf_1
Xinput325 la_iena_mprj[43] vssd vssd vccd vccd net325 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput326 la_iena_mprj[44] vssd vssd vccd vccd net326 sky130_fd_sc_hd__clkbuf_1
Xinput327 la_iena_mprj[45] vssd vssd vccd vccd net327 sky130_fd_sc_hd__clkbuf_1
Xinput328 la_iena_mprj[46] vssd vssd vccd vccd net328 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput329 la_iena_mprj[47] vssd vssd vccd vccd net329 sky130_fd_sc_hd__clkbuf_1
Xinput33 la_data_out_core[126] vssd vssd vccd vccd net33 sky130_fd_sc_hd__clkbuf_4
Xinput330 la_iena_mprj[48] vssd vssd vccd vccd net330 sky130_fd_sc_hd__clkbuf_1
Xinput331 la_iena_mprj[49] vssd vssd vccd vccd net331 sky130_fd_sc_hd__clkbuf_1
Xinput332 la_iena_mprj[4] vssd vssd vccd vccd net332 sky130_fd_sc_hd__buf_2
Xinput333 la_iena_mprj[50] vssd vssd vccd vccd net333 sky130_fd_sc_hd__clkbuf_1
Xinput334 la_iena_mprj[51] vssd vssd vccd vccd net334 sky130_fd_sc_hd__clkbuf_1
Xinput335 la_iena_mprj[52] vssd vssd vccd vccd net335 sky130_fd_sc_hd__clkbuf_1
Xinput336 la_iena_mprj[53] vssd vssd vccd vccd net336 sky130_fd_sc_hd__clkbuf_1
Xinput337 la_iena_mprj[54] vssd vssd vccd vccd net337 sky130_fd_sc_hd__clkbuf_1
Xinput338 la_iena_mprj[55] vssd vssd vccd vccd net338 sky130_fd_sc_hd__clkbuf_1
Xinput339 la_iena_mprj[56] vssd vssd vccd vccd net339 sky130_fd_sc_hd__clkbuf_1
Xinput34 la_data_out_core[127] vssd vssd vccd vccd net34 sky130_fd_sc_hd__clkbuf_4
Xinput340 la_iena_mprj[57] vssd vssd vccd vccd net340 sky130_fd_sc_hd__clkbuf_1
Xinput341 la_iena_mprj[58] vssd vssd vccd vccd net341 sky130_fd_sc_hd__clkbuf_1
Xinput342 la_iena_mprj[59] vssd vssd vccd vccd net342 sky130_fd_sc_hd__clkbuf_1
Xinput343 la_iena_mprj[5] vssd vssd vccd vccd net343 sky130_fd_sc_hd__buf_2
Xinput344 la_iena_mprj[60] vssd vssd vccd vccd net344 sky130_fd_sc_hd__clkbuf_1
Xinput345 la_iena_mprj[61] vssd vssd vccd vccd net345 sky130_fd_sc_hd__clkbuf_1
Xinput346 la_iena_mprj[62] vssd vssd vccd vccd net346 sky130_fd_sc_hd__clkbuf_1
Xinput347 la_iena_mprj[63] vssd vssd vccd vccd net347 sky130_fd_sc_hd__clkbuf_1
Xinput348 la_iena_mprj[64] vssd vssd vccd vccd net348 sky130_fd_sc_hd__clkbuf_1
Xinput349 la_iena_mprj[65] vssd vssd vccd vccd net349 sky130_fd_sc_hd__clkbuf_1
Xinput35 la_data_out_core[12] vssd vssd vccd vccd net35 sky130_fd_sc_hd__clkbuf_2
Xinput350 la_iena_mprj[66] vssd vssd vccd vccd net350 sky130_fd_sc_hd__clkbuf_1
Xinput351 la_iena_mprj[67] vssd vssd vccd vccd net351 sky130_fd_sc_hd__clkbuf_1
Xinput352 la_iena_mprj[68] vssd vssd vccd vccd net352 sky130_fd_sc_hd__clkbuf_1
Xinput353 la_iena_mprj[69] vssd vssd vccd vccd net353 sky130_fd_sc_hd__clkbuf_1
Xinput354 la_iena_mprj[6] vssd vssd vccd vccd net354 sky130_fd_sc_hd__clkbuf_2
Xinput355 la_iena_mprj[70] vssd vssd vccd vccd net355 sky130_fd_sc_hd__clkbuf_1
Xinput356 la_iena_mprj[71] vssd vssd vccd vccd net356 sky130_fd_sc_hd__clkbuf_1
Xinput357 la_iena_mprj[72] vssd vssd vccd vccd net357 sky130_fd_sc_hd__clkbuf_1
Xinput358 la_iena_mprj[73] vssd vssd vccd vccd net358 sky130_fd_sc_hd__clkbuf_1
Xinput359 la_iena_mprj[74] vssd vssd vccd vccd net359 sky130_fd_sc_hd__clkbuf_1
Xinput36 la_data_out_core[13] vssd vssd vccd vccd net36 sky130_fd_sc_hd__buf_4
Xinput360 la_iena_mprj[75] vssd vssd vccd vccd net360 sky130_fd_sc_hd__clkbuf_1
Xinput361 la_iena_mprj[76] vssd vssd vccd vccd net361 sky130_fd_sc_hd__clkbuf_1
Xinput362 la_iena_mprj[77] vssd vssd vccd vccd net362 sky130_fd_sc_hd__clkbuf_1
Xinput363 la_iena_mprj[78] vssd vssd vccd vccd net363 sky130_fd_sc_hd__clkbuf_1
Xinput364 la_iena_mprj[79] vssd vssd vccd vccd net364 sky130_fd_sc_hd__clkbuf_1
Xinput365 la_iena_mprj[7] vssd vssd vccd vccd net365 sky130_fd_sc_hd__clkbuf_4
Xinput366 la_iena_mprj[80] vssd vssd vccd vccd net366 sky130_fd_sc_hd__clkbuf_1
Xinput367 la_iena_mprj[81] vssd vssd vccd vccd net367 sky130_fd_sc_hd__clkbuf_1
Xinput368 la_iena_mprj[82] vssd vssd vccd vccd net368 sky130_fd_sc_hd__clkbuf_1
Xinput369 la_iena_mprj[83] vssd vssd vccd vccd net369 sky130_fd_sc_hd__clkbuf_1
Xinput37 la_data_out_core[14] vssd vssd vccd vccd net37 sky130_fd_sc_hd__buf_4
Xinput370 la_iena_mprj[84] vssd vssd vccd vccd net370 sky130_fd_sc_hd__clkbuf_1
Xinput371 la_iena_mprj[85] vssd vssd vccd vccd net371 sky130_fd_sc_hd__clkbuf_1
Xinput372 la_iena_mprj[86] vssd vssd vccd vccd net372 sky130_fd_sc_hd__clkbuf_1
Xinput373 la_iena_mprj[87] vssd vssd vccd vccd net373 sky130_fd_sc_hd__clkbuf_1
Xinput374 la_iena_mprj[88] vssd vssd vccd vccd net374 sky130_fd_sc_hd__clkbuf_1
Xinput375 la_iena_mprj[89] vssd vssd vccd vccd net375 sky130_fd_sc_hd__clkbuf_1
Xinput376 la_iena_mprj[8] vssd vssd vccd vccd net376 sky130_fd_sc_hd__clkbuf_4
Xinput377 la_iena_mprj[90] vssd vssd vccd vccd net377 sky130_fd_sc_hd__clkbuf_1
Xinput378 la_iena_mprj[91] vssd vssd vccd vccd net378 sky130_fd_sc_hd__clkbuf_1
Xinput379 la_iena_mprj[92] vssd vssd vccd vccd net379 sky130_fd_sc_hd__clkbuf_1
Xinput38 la_data_out_core[15] vssd vssd vccd vccd net38 sky130_fd_sc_hd__buf_4
Xinput380 la_iena_mprj[93] vssd vssd vccd vccd net380 sky130_fd_sc_hd__clkbuf_1
Xinput381 la_iena_mprj[94] vssd vssd vccd vccd net381 sky130_fd_sc_hd__clkbuf_1
Xinput382 la_iena_mprj[95] vssd vssd vccd vccd net382 sky130_fd_sc_hd__clkbuf_1
Xinput383 la_iena_mprj[96] vssd vssd vccd vccd net383 sky130_fd_sc_hd__clkbuf_1
Xinput384 la_iena_mprj[97] vssd vssd vccd vccd net384 sky130_fd_sc_hd__clkbuf_1
Xinput385 la_iena_mprj[98] vssd vssd vccd vccd net385 sky130_fd_sc_hd__clkbuf_1
Xinput386 la_iena_mprj[99] vssd vssd vccd vccd net386 sky130_fd_sc_hd__clkbuf_1
Xinput387 la_iena_mprj[9] vssd vssd vccd vccd net387 sky130_fd_sc_hd__buf_2
Xinput388 la_oenb_mprj[0] vssd vssd vccd vccd net388 sky130_fd_sc_hd__clkbuf_2
Xinput389 la_oenb_mprj[100] vssd vssd vccd vccd net389 sky130_fd_sc_hd__clkbuf_4
Xinput39 la_data_out_core[16] vssd vssd vccd vccd net39 sky130_fd_sc_hd__clkbuf_4
Xinput390 la_oenb_mprj[101] vssd vssd vccd vccd net390 sky130_fd_sc_hd__clkbuf_4
Xinput391 la_oenb_mprj[102] vssd vssd vccd vccd net391 sky130_fd_sc_hd__clkbuf_4
Xinput392 la_oenb_mprj[103] vssd vssd vccd vccd net392 sky130_fd_sc_hd__clkbuf_4
Xinput393 la_oenb_mprj[104] vssd vssd vccd vccd net393 sky130_fd_sc_hd__buf_2
Xinput394 la_oenb_mprj[105] vssd vssd vccd vccd net394 sky130_fd_sc_hd__buf_4
Xinput395 la_oenb_mprj[106] vssd vssd vccd vccd net395 sky130_fd_sc_hd__buf_2
Xinput396 la_oenb_mprj[107] vssd vssd vccd vccd net396 sky130_fd_sc_hd__clkbuf_4
Xinput397 la_oenb_mprj[108] vssd vssd vccd vccd net397 sky130_fd_sc_hd__buf_4
Xinput398 la_oenb_mprj[109] vssd vssd vccd vccd net398 sky130_fd_sc_hd__clkbuf_4
Xinput399 la_oenb_mprj[10] vssd vssd vccd vccd net399 sky130_fd_sc_hd__clkbuf_2
Xinput4 la_data_out_core[0] vssd vssd vccd vccd net4 sky130_fd_sc_hd__buf_4
Xinput40 la_data_out_core[17] vssd vssd vccd vccd net40 sky130_fd_sc_hd__buf_4
Xinput400 la_oenb_mprj[110] vssd vssd vccd vccd net400 sky130_fd_sc_hd__clkbuf_4
Xinput401 la_oenb_mprj[111] vssd vssd vccd vccd net401 sky130_fd_sc_hd__buf_4
Xinput402 la_oenb_mprj[112] vssd vssd vccd vccd net402 sky130_fd_sc_hd__buf_2
Xinput403 la_oenb_mprj[113] vssd vssd vccd vccd net403 sky130_fd_sc_hd__clkbuf_4
Xinput404 la_oenb_mprj[114] vssd vssd vccd vccd net404 sky130_fd_sc_hd__clkbuf_4
Xinput405 la_oenb_mprj[115] vssd vssd vccd vccd net405 sky130_fd_sc_hd__clkbuf_4
Xinput406 la_oenb_mprj[116] vssd vssd vccd vccd net406 sky130_fd_sc_hd__clkbuf_4
Xinput407 la_oenb_mprj[117] vssd vssd vccd vccd net407 sky130_fd_sc_hd__clkbuf_4
Xinput408 la_oenb_mprj[118] vssd vssd vccd vccd net408 sky130_fd_sc_hd__clkbuf_4
Xinput409 la_oenb_mprj[119] vssd vssd vccd vccd net409 sky130_fd_sc_hd__clkbuf_4
Xinput41 la_data_out_core[18] vssd vssd vccd vccd net41 sky130_fd_sc_hd__buf_4
Xinput410 la_oenb_mprj[11] vssd vssd vccd vccd net410 sky130_fd_sc_hd__clkbuf_2
Xinput411 la_oenb_mprj[120] vssd vssd vccd vccd net411 sky130_fd_sc_hd__clkbuf_2
Xinput412 la_oenb_mprj[121] vssd vssd vccd vccd net412 sky130_fd_sc_hd__clkbuf_4
Xinput413 la_oenb_mprj[122] vssd vssd vccd vccd net413 sky130_fd_sc_hd__clkbuf_4
Xinput414 la_oenb_mprj[123] vssd vssd vccd vccd net414 sky130_fd_sc_hd__clkbuf_4
Xinput415 la_oenb_mprj[124] vssd vssd vccd vccd net415 sky130_fd_sc_hd__clkbuf_4
Xinput416 la_oenb_mprj[125] vssd vssd vccd vccd net416 sky130_fd_sc_hd__clkbuf_4
Xinput417 la_oenb_mprj[126] vssd vssd vccd vccd net417 sky130_fd_sc_hd__clkbuf_4
Xinput418 la_oenb_mprj[127] vssd vssd vccd vccd net418 sky130_fd_sc_hd__clkbuf_4
Xinput419 la_oenb_mprj[12] vssd vssd vccd vccd net419 sky130_fd_sc_hd__buf_2
Xinput42 la_data_out_core[19] vssd vssd vccd vccd net42 sky130_fd_sc_hd__buf_4
Xinput420 la_oenb_mprj[13] vssd vssd vccd vccd net420 sky130_fd_sc_hd__clkbuf_2
Xinput421 la_oenb_mprj[14] vssd vssd vccd vccd net421 sky130_fd_sc_hd__buf_2
Xinput422 la_oenb_mprj[15] vssd vssd vccd vccd net422 sky130_fd_sc_hd__clkbuf_2
Xinput423 la_oenb_mprj[16] vssd vssd vccd vccd net423 sky130_fd_sc_hd__clkbuf_2
Xinput424 la_oenb_mprj[17] vssd vssd vccd vccd net424 sky130_fd_sc_hd__buf_2
Xinput425 la_oenb_mprj[18] vssd vssd vccd vccd net425 sky130_fd_sc_hd__clkbuf_2
Xinput426 la_oenb_mprj[19] vssd vssd vccd vccd net426 sky130_fd_sc_hd__clkbuf_2
Xinput427 la_oenb_mprj[1] vssd vssd vccd vccd net427 sky130_fd_sc_hd__buf_2
Xinput428 la_oenb_mprj[20] vssd vssd vccd vccd net428 sky130_fd_sc_hd__clkbuf_2
Xinput429 la_oenb_mprj[21] vssd vssd vccd vccd net429 sky130_fd_sc_hd__buf_2
Xinput43 la_data_out_core[1] vssd vssd vccd vccd net43 sky130_fd_sc_hd__buf_4
Xinput430 la_oenb_mprj[22] vssd vssd vccd vccd net430 sky130_fd_sc_hd__clkbuf_2
Xinput431 la_oenb_mprj[23] vssd vssd vccd vccd net431 sky130_fd_sc_hd__buf_2
Xinput432 la_oenb_mprj[24] vssd vssd vccd vccd net432 sky130_fd_sc_hd__clkbuf_4
Xinput433 la_oenb_mprj[25] vssd vssd vccd vccd net433 sky130_fd_sc_hd__buf_2
Xinput434 la_oenb_mprj[26] vssd vssd vccd vccd net434 sky130_fd_sc_hd__clkbuf_2
Xinput435 la_oenb_mprj[27] vssd vssd vccd vccd net435 sky130_fd_sc_hd__buf_2
Xinput436 la_oenb_mprj[28] vssd vssd vccd vccd net436 sky130_fd_sc_hd__clkbuf_4
Xinput437 la_oenb_mprj[29] vssd vssd vccd vccd net437 sky130_fd_sc_hd__buf_2
Xinput438 la_oenb_mprj[2] vssd vssd vccd vccd net438 sky130_fd_sc_hd__buf_2
Xinput439 la_oenb_mprj[30] vssd vssd vccd vccd net439 sky130_fd_sc_hd__buf_2
Xinput44 la_data_out_core[20] vssd vssd vccd vccd net44 sky130_fd_sc_hd__clkbuf_4
Xinput440 la_oenb_mprj[31] vssd vssd vccd vccd net440 sky130_fd_sc_hd__buf_2
Xinput441 la_oenb_mprj[32] vssd vssd vccd vccd net441 sky130_fd_sc_hd__buf_2
Xinput442 la_oenb_mprj[33] vssd vssd vccd vccd net442 sky130_fd_sc_hd__buf_2
Xinput443 la_oenb_mprj[34] vssd vssd vccd vccd net443 sky130_fd_sc_hd__clkbuf_2
Xinput444 la_oenb_mprj[35] vssd vssd vccd vccd net444 sky130_fd_sc_hd__clkbuf_2
Xinput445 la_oenb_mprj[36] vssd vssd vccd vccd net445 sky130_fd_sc_hd__clkbuf_2
Xinput446 la_oenb_mprj[37] vssd vssd vccd vccd net446 sky130_fd_sc_hd__clkbuf_2
Xinput447 la_oenb_mprj[38] vssd vssd vccd vccd net447 sky130_fd_sc_hd__clkbuf_2
Xinput448 la_oenb_mprj[39] vssd vssd vccd vccd net448 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput449 la_oenb_mprj[3] vssd vssd vccd vccd net449 sky130_fd_sc_hd__clkbuf_2
Xinput45 la_data_out_core[21] vssd vssd vccd vccd net45 sky130_fd_sc_hd__clkbuf_4
Xinput450 la_oenb_mprj[40] vssd vssd vccd vccd net450 sky130_fd_sc_hd__buf_4
Xinput451 la_oenb_mprj[41] vssd vssd vccd vccd net451 sky130_fd_sc_hd__clkbuf_2
Xinput452 la_oenb_mprj[42] vssd vssd vccd vccd net452 sky130_fd_sc_hd__clkbuf_4
Xinput453 la_oenb_mprj[43] vssd vssd vccd vccd net453 sky130_fd_sc_hd__buf_4
Xinput454 la_oenb_mprj[44] vssd vssd vccd vccd net454 sky130_fd_sc_hd__buf_2
Xinput455 la_oenb_mprj[45] vssd vssd vccd vccd net455 sky130_fd_sc_hd__clkbuf_2
Xinput456 la_oenb_mprj[46] vssd vssd vccd vccd net456 sky130_fd_sc_hd__buf_4
Xinput457 la_oenb_mprj[47] vssd vssd vccd vccd net457 sky130_fd_sc_hd__buf_4
Xinput458 la_oenb_mprj[48] vssd vssd vccd vccd net458 sky130_fd_sc_hd__buf_2
Xinput459 la_oenb_mprj[49] vssd vssd vccd vccd net459 sky130_fd_sc_hd__clkbuf_4
Xinput46 la_data_out_core[22] vssd vssd vccd vccd net46 sky130_fd_sc_hd__buf_4
Xinput460 la_oenb_mprj[4] vssd vssd vccd vccd net460 sky130_fd_sc_hd__buf_2
Xinput461 la_oenb_mprj[50] vssd vssd vccd vccd net461 sky130_fd_sc_hd__clkbuf_2
Xinput462 la_oenb_mprj[51] vssd vssd vccd vccd net462 sky130_fd_sc_hd__buf_2
Xinput463 la_oenb_mprj[52] vssd vssd vccd vccd net463 sky130_fd_sc_hd__clkbuf_2
Xinput464 la_oenb_mprj[53] vssd vssd vccd vccd net464 sky130_fd_sc_hd__buf_2
Xinput465 la_oenb_mprj[54] vssd vssd vccd vccd net465 sky130_fd_sc_hd__clkbuf_2
Xinput466 la_oenb_mprj[55] vssd vssd vccd vccd net466 sky130_fd_sc_hd__buf_2
Xinput467 la_oenb_mprj[56] vssd vssd vccd vccd net467 sky130_fd_sc_hd__clkbuf_2
Xinput468 la_oenb_mprj[57] vssd vssd vccd vccd net468 sky130_fd_sc_hd__clkbuf_2
Xinput469 la_oenb_mprj[58] vssd vssd vccd vccd net469 sky130_fd_sc_hd__buf_2
Xinput47 la_data_out_core[23] vssd vssd vccd vccd net47 sky130_fd_sc_hd__buf_4
Xinput470 la_oenb_mprj[59] vssd vssd vccd vccd net470 sky130_fd_sc_hd__clkbuf_2
Xinput471 la_oenb_mprj[5] vssd vssd vccd vccd net471 sky130_fd_sc_hd__buf_2
Xinput472 la_oenb_mprj[60] vssd vssd vccd vccd net472 sky130_fd_sc_hd__buf_2
Xinput473 la_oenb_mprj[61] vssd vssd vccd vccd net473 sky130_fd_sc_hd__buf_2
Xinput474 la_oenb_mprj[62] vssd vssd vccd vccd net474 sky130_fd_sc_hd__buf_2
Xinput475 la_oenb_mprj[63] vssd vssd vccd vccd net475 sky130_fd_sc_hd__clkbuf_2
Xinput476 la_oenb_mprj[64] vssd vssd vccd vccd net476 sky130_fd_sc_hd__buf_2
Xinput477 la_oenb_mprj[65] vssd vssd vccd vccd net477 sky130_fd_sc_hd__clkbuf_2
Xinput478 la_oenb_mprj[66] vssd vssd vccd vccd net478 sky130_fd_sc_hd__buf_4
Xinput479 la_oenb_mprj[67] vssd vssd vccd vccd net479 sky130_fd_sc_hd__buf_4
Xinput48 la_data_out_core[24] vssd vssd vccd vccd net48 sky130_fd_sc_hd__buf_4
Xinput480 la_oenb_mprj[68] vssd vssd vccd vccd net480 sky130_fd_sc_hd__clkbuf_2
Xinput481 la_oenb_mprj[69] vssd vssd vccd vccd net481 sky130_fd_sc_hd__clkbuf_2
Xinput482 la_oenb_mprj[6] vssd vssd vccd vccd net482 sky130_fd_sc_hd__clkbuf_2
Xinput483 la_oenb_mprj[70] vssd vssd vccd vccd net483 sky130_fd_sc_hd__buf_2
Xinput484 la_oenb_mprj[71] vssd vssd vccd vccd net484 sky130_fd_sc_hd__clkbuf_2
Xinput485 la_oenb_mprj[72] vssd vssd vccd vccd net485 sky130_fd_sc_hd__buf_2
Xinput486 la_oenb_mprj[73] vssd vssd vccd vccd net486 sky130_fd_sc_hd__clkbuf_4
Xinput487 la_oenb_mprj[74] vssd vssd vccd vccd net487 sky130_fd_sc_hd__buf_2
Xinput488 la_oenb_mprj[75] vssd vssd vccd vccd net488 sky130_fd_sc_hd__buf_2
Xinput489 la_oenb_mprj[76] vssd vssd vccd vccd net489 sky130_fd_sc_hd__clkbuf_4
Xinput49 la_data_out_core[25] vssd vssd vccd vccd net49 sky130_fd_sc_hd__buf_4
Xinput490 la_oenb_mprj[77] vssd vssd vccd vccd net490 sky130_fd_sc_hd__clkbuf_4
Xinput491 la_oenb_mprj[78] vssd vssd vccd vccd net491 sky130_fd_sc_hd__clkbuf_4
Xinput492 la_oenb_mprj[79] vssd vssd vccd vccd net492 sky130_fd_sc_hd__clkbuf_4
Xinput493 la_oenb_mprj[7] vssd vssd vccd vccd net493 sky130_fd_sc_hd__buf_2
Xinput494 la_oenb_mprj[80] vssd vssd vccd vccd net494 sky130_fd_sc_hd__clkbuf_4
Xinput495 la_oenb_mprj[81] vssd vssd vccd vccd net495 sky130_fd_sc_hd__buf_4
Xinput496 la_oenb_mprj[82] vssd vssd vccd vccd net496 sky130_fd_sc_hd__clkbuf_4
Xinput497 la_oenb_mprj[83] vssd vssd vccd vccd net497 sky130_fd_sc_hd__buf_4
Xinput498 la_oenb_mprj[84] vssd vssd vccd vccd net498 sky130_fd_sc_hd__buf_4
Xinput499 la_oenb_mprj[85] vssd vssd vccd vccd net499 sky130_fd_sc_hd__buf_4
Xinput5 la_data_out_core[100] vssd vssd vccd vccd net5 sky130_fd_sc_hd__clkbuf_4
Xinput50 la_data_out_core[26] vssd vssd vccd vccd net50 sky130_fd_sc_hd__buf_4
Xinput500 la_oenb_mprj[86] vssd vssd vccd vccd net500 sky130_fd_sc_hd__buf_4
Xinput501 la_oenb_mprj[87] vssd vssd vccd vccd net501 sky130_fd_sc_hd__clkbuf_4
Xinput502 la_oenb_mprj[88] vssd vssd vccd vccd net502 sky130_fd_sc_hd__buf_4
Xinput503 la_oenb_mprj[89] vssd vssd vccd vccd net503 sky130_fd_sc_hd__buf_4
Xinput504 la_oenb_mprj[8] vssd vssd vccd vccd net504 sky130_fd_sc_hd__buf_2
Xinput505 la_oenb_mprj[90] vssd vssd vccd vccd net505 sky130_fd_sc_hd__clkbuf_4
Xinput506 la_oenb_mprj[91] vssd vssd vccd vccd net506 sky130_fd_sc_hd__clkbuf_4
Xinput507 la_oenb_mprj[92] vssd vssd vccd vccd net507 sky130_fd_sc_hd__clkbuf_4
Xinput508 la_oenb_mprj[93] vssd vssd vccd vccd net508 sky130_fd_sc_hd__buf_2
Xinput509 la_oenb_mprj[94] vssd vssd vccd vccd net509 sky130_fd_sc_hd__buf_4
Xinput51 la_data_out_core[27] vssd vssd vccd vccd net51 sky130_fd_sc_hd__clkbuf_4
Xinput510 la_oenb_mprj[95] vssd vssd vccd vccd net510 sky130_fd_sc_hd__clkbuf_4
Xinput511 la_oenb_mprj[96] vssd vssd vccd vccd net511 sky130_fd_sc_hd__clkbuf_2
Xinput512 la_oenb_mprj[97] vssd vssd vccd vccd net512 sky130_fd_sc_hd__clkbuf_4
Xinput513 la_oenb_mprj[98] vssd vssd vccd vccd net513 sky130_fd_sc_hd__clkbuf_4
Xinput514 la_oenb_mprj[99] vssd vssd vccd vccd net514 sky130_fd_sc_hd__clkbuf_4
Xinput515 la_oenb_mprj[9] vssd vssd vccd vccd net515 sky130_fd_sc_hd__clkbuf_2
Xinput516 mprj_ack_i_user vssd vssd vccd vccd net516 sky130_fd_sc_hd__buf_8
Xinput517 mprj_adr_o_core[0] vssd vssd vccd vccd net517 sky130_fd_sc_hd__buf_12
Xinput518 mprj_adr_o_core[10] vssd vssd vccd vccd net518 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput519 mprj_adr_o_core[11] vssd vssd vccd vccd net519 sky130_fd_sc_hd__clkbuf_1
Xinput52 la_data_out_core[28] vssd vssd vccd vccd net52 sky130_fd_sc_hd__clkbuf_4
Xinput520 mprj_adr_o_core[12] vssd vssd vccd vccd net520 sky130_fd_sc_hd__buf_2
Xinput521 mprj_adr_o_core[13] vssd vssd vccd vccd net521 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput522 mprj_adr_o_core[14] vssd vssd vccd vccd net522 sky130_fd_sc_hd__clkbuf_2
Xinput523 mprj_adr_o_core[15] vssd vssd vccd vccd net523 sky130_fd_sc_hd__buf_2
Xinput524 mprj_adr_o_core[16] vssd vssd vccd vccd net524 sky130_fd_sc_hd__buf_2
Xinput525 mprj_adr_o_core[17] vssd vssd vccd vccd net525 sky130_fd_sc_hd__clkbuf_2
Xinput526 mprj_adr_o_core[18] vssd vssd vccd vccd net526 sky130_fd_sc_hd__buf_2
Xinput527 mprj_adr_o_core[19] vssd vssd vccd vccd net527 sky130_fd_sc_hd__clkbuf_4
Xinput528 mprj_adr_o_core[1] vssd vssd vccd vccd net528 sky130_fd_sc_hd__buf_2
Xinput529 mprj_adr_o_core[20] vssd vssd vccd vccd net529 sky130_fd_sc_hd__clkbuf_2
Xinput53 la_data_out_core[29] vssd vssd vccd vccd net53 sky130_fd_sc_hd__clkbuf_4
Xinput530 mprj_adr_o_core[21] vssd vssd vccd vccd net530 sky130_fd_sc_hd__buf_2
Xinput531 mprj_adr_o_core[22] vssd vssd vccd vccd net531 sky130_fd_sc_hd__clkbuf_2
Xinput532 mprj_adr_o_core[23] vssd vssd vccd vccd net532 sky130_fd_sc_hd__clkbuf_2
Xinput533 mprj_adr_o_core[24] vssd vssd vccd vccd net533 sky130_fd_sc_hd__buf_4
Xinput534 mprj_adr_o_core[25] vssd vssd vccd vccd net534 sky130_fd_sc_hd__clkbuf_4
Xinput535 mprj_adr_o_core[26] vssd vssd vccd vccd net535 sky130_fd_sc_hd__clkbuf_4
Xinput536 mprj_adr_o_core[27] vssd vssd vccd vccd net536 sky130_fd_sc_hd__buf_2
Xinput537 mprj_adr_o_core[28] vssd vssd vccd vccd net537 sky130_fd_sc_hd__buf_2
Xinput538 mprj_adr_o_core[29] vssd vssd vccd vccd net538 sky130_fd_sc_hd__buf_2
Xinput539 mprj_adr_o_core[2] vssd vssd vccd vccd net539 sky130_fd_sc_hd__buf_12
Xinput54 la_data_out_core[2] vssd vssd vccd vccd net54 sky130_fd_sc_hd__buf_4
Xinput540 mprj_adr_o_core[30] vssd vssd vccd vccd net540 sky130_fd_sc_hd__buf_2
Xinput541 mprj_adr_o_core[31] vssd vssd vccd vccd net541 sky130_fd_sc_hd__clkbuf_2
Xinput542 mprj_adr_o_core[3] vssd vssd vccd vccd net542 sky130_fd_sc_hd__buf_2
Xinput543 mprj_adr_o_core[4] vssd vssd vccd vccd net543 sky130_fd_sc_hd__buf_12
Xinput544 mprj_adr_o_core[5] vssd vssd vccd vccd net544 sky130_fd_sc_hd__clkbuf_4
Xinput545 mprj_adr_o_core[6] vssd vssd vccd vccd net545 sky130_fd_sc_hd__clkbuf_2
Xinput546 mprj_adr_o_core[7] vssd vssd vccd vccd net546 sky130_fd_sc_hd__clkbuf_2
Xinput547 mprj_adr_o_core[8] vssd vssd vccd vccd net547 sky130_fd_sc_hd__clkbuf_4
Xinput548 mprj_adr_o_core[9] vssd vssd vccd vccd net548 sky130_fd_sc_hd__clkbuf_2
Xinput549 mprj_cyc_o_core vssd vssd vccd vccd net549 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput55 la_data_out_core[30] vssd vssd vccd vccd net55 sky130_fd_sc_hd__buf_4
Xinput550 mprj_dat_i_user[0] vssd vssd vccd vccd net550 sky130_fd_sc_hd__buf_8
Xinput551 mprj_dat_i_user[10] vssd vssd vccd vccd net551 sky130_fd_sc_hd__buf_8
Xinput552 mprj_dat_i_user[11] vssd vssd vccd vccd net552 sky130_fd_sc_hd__buf_12
Xinput553 mprj_dat_i_user[12] vssd vssd vccd vccd net553 sky130_fd_sc_hd__buf_8
Xinput554 mprj_dat_i_user[13] vssd vssd vccd vccd net554 sky130_fd_sc_hd__buf_8
Xinput555 mprj_dat_i_user[14] vssd vssd vccd vccd net555 sky130_fd_sc_hd__buf_12
Xinput556 mprj_dat_i_user[15] vssd vssd vccd vccd net556 sky130_fd_sc_hd__buf_12
Xinput557 mprj_dat_i_user[16] vssd vssd vccd vccd net557 sky130_fd_sc_hd__clkbuf_16
Xinput558 mprj_dat_i_user[17] vssd vssd vccd vccd net558 sky130_fd_sc_hd__buf_12
Xinput559 mprj_dat_i_user[18] vssd vssd vccd vccd net559 sky130_fd_sc_hd__buf_12
Xinput56 la_data_out_core[31] vssd vssd vccd vccd net56 sky130_fd_sc_hd__clkbuf_4
Xinput560 mprj_dat_i_user[19] vssd vssd vccd vccd net560 sky130_fd_sc_hd__buf_8
Xinput561 mprj_dat_i_user[1] vssd vssd vccd vccd net561 sky130_fd_sc_hd__buf_8
Xinput562 mprj_dat_i_user[20] vssd vssd vccd vccd net562 sky130_fd_sc_hd__clkbuf_16
Xinput563 mprj_dat_i_user[21] vssd vssd vccd vccd net563 sky130_fd_sc_hd__buf_12
Xinput564 mprj_dat_i_user[22] vssd vssd vccd vccd net564 sky130_fd_sc_hd__buf_12
Xinput565 mprj_dat_i_user[23] vssd vssd vccd vccd net565 sky130_fd_sc_hd__buf_12
Xinput566 mprj_dat_i_user[24] vssd vssd vccd vccd net566 sky130_fd_sc_hd__buf_12
Xinput567 mprj_dat_i_user[25] vssd vssd vccd vccd net567 sky130_fd_sc_hd__buf_12
Xinput568 mprj_dat_i_user[26] vssd vssd vccd vccd net568 sky130_fd_sc_hd__buf_8
Xinput569 mprj_dat_i_user[27] vssd vssd vccd vccd net569 sky130_fd_sc_hd__buf_8
Xinput57 la_data_out_core[32] vssd vssd vccd vccd net57 sky130_fd_sc_hd__buf_4
Xinput570 mprj_dat_i_user[28] vssd vssd vccd vccd net570 sky130_fd_sc_hd__buf_8
Xinput571 mprj_dat_i_user[29] vssd vssd vccd vccd net571 sky130_fd_sc_hd__clkbuf_16
Xinput572 mprj_dat_i_user[2] vssd vssd vccd vccd net572 sky130_fd_sc_hd__buf_8
Xinput573 mprj_dat_i_user[30] vssd vssd vccd vccd net573 sky130_fd_sc_hd__buf_12
Xinput574 mprj_dat_i_user[31] vssd vssd vccd vccd net574 sky130_fd_sc_hd__buf_12
Xinput575 mprj_dat_i_user[3] vssd vssd vccd vccd net575 sky130_fd_sc_hd__buf_6
Xinput576 mprj_dat_i_user[4] vssd vssd vccd vccd net576 sky130_fd_sc_hd__buf_6
Xinput577 mprj_dat_i_user[5] vssd vssd vccd vccd net577 sky130_fd_sc_hd__buf_8
Xinput578 mprj_dat_i_user[6] vssd vssd vccd vccd net578 sky130_fd_sc_hd__buf_8
Xinput579 mprj_dat_i_user[7] vssd vssd vccd vccd net579 sky130_fd_sc_hd__buf_8
Xinput58 la_data_out_core[33] vssd vssd vccd vccd net58 sky130_fd_sc_hd__clkbuf_4
Xinput580 mprj_dat_i_user[8] vssd vssd vccd vccd net580 sky130_fd_sc_hd__buf_8
Xinput581 mprj_dat_i_user[9] vssd vssd vccd vccd net581 sky130_fd_sc_hd__buf_8
Xinput582 mprj_dat_o_core[0] vssd vssd vccd vccd net582 sky130_fd_sc_hd__clkbuf_8
Xinput583 mprj_dat_o_core[10] vssd vssd vccd vccd net583 sky130_fd_sc_hd__clkbuf_4
Xinput584 mprj_dat_o_core[11] vssd vssd vccd vccd net584 sky130_fd_sc_hd__clkbuf_4
Xinput585 mprj_dat_o_core[12] vssd vssd vccd vccd net585 sky130_fd_sc_hd__clkbuf_4
Xinput586 mprj_dat_o_core[13] vssd vssd vccd vccd net586 sky130_fd_sc_hd__clkbuf_4
Xinput587 mprj_dat_o_core[14] vssd vssd vccd vccd net587 sky130_fd_sc_hd__buf_4
Xinput588 mprj_dat_o_core[15] vssd vssd vccd vccd net588 sky130_fd_sc_hd__buf_4
Xinput589 mprj_dat_o_core[16] vssd vssd vccd vccd net589 sky130_fd_sc_hd__clkbuf_4
Xinput59 la_data_out_core[34] vssd vssd vccd vccd net59 sky130_fd_sc_hd__clkbuf_4
Xinput590 mprj_dat_o_core[17] vssd vssd vccd vccd net590 sky130_fd_sc_hd__clkbuf_2
Xinput591 mprj_dat_o_core[18] vssd vssd vccd vccd net591 sky130_fd_sc_hd__clkbuf_2
Xinput592 mprj_dat_o_core[19] vssd vssd vccd vccd net592 sky130_fd_sc_hd__clkbuf_2
Xinput593 mprj_dat_o_core[1] vssd vssd vccd vccd net593 sky130_fd_sc_hd__clkbuf_4
Xinput594 mprj_dat_o_core[20] vssd vssd vccd vccd net594 sky130_fd_sc_hd__clkbuf_2
Xinput595 mprj_dat_o_core[21] vssd vssd vccd vccd net595 sky130_fd_sc_hd__clkbuf_2
Xinput596 mprj_dat_o_core[22] vssd vssd vccd vccd net596 sky130_fd_sc_hd__clkbuf_2
Xinput597 mprj_dat_o_core[23] vssd vssd vccd vccd net597 sky130_fd_sc_hd__buf_2
Xinput598 mprj_dat_o_core[24] vssd vssd vccd vccd net598 sky130_fd_sc_hd__clkbuf_2
Xinput599 mprj_dat_o_core[25] vssd vssd vccd vccd net599 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput6 la_data_out_core[101] vssd vssd vccd vccd net6 sky130_fd_sc_hd__clkbuf_4
Xinput60 la_data_out_core[35] vssd vssd vccd vccd net60 sky130_fd_sc_hd__buf_4
Xinput600 mprj_dat_o_core[26] vssd vssd vccd vccd net600 sky130_fd_sc_hd__clkbuf_2
Xinput601 mprj_dat_o_core[27] vssd vssd vccd vccd net601 sky130_fd_sc_hd__buf_2
Xinput602 mprj_dat_o_core[28] vssd vssd vccd vccd net602 sky130_fd_sc_hd__clkbuf_2
Xinput603 mprj_dat_o_core[29] vssd vssd vccd vccd net603 sky130_fd_sc_hd__clkbuf_2
Xinput604 mprj_dat_o_core[2] vssd vssd vccd vccd net604 sky130_fd_sc_hd__buf_4
Xinput605 mprj_dat_o_core[30] vssd vssd vccd vccd net605 sky130_fd_sc_hd__buf_2
Xinput606 mprj_dat_o_core[31] vssd vssd vccd vccd net606 sky130_fd_sc_hd__clkbuf_2
Xinput607 mprj_dat_o_core[3] vssd vssd vccd vccd net607 sky130_fd_sc_hd__buf_2
Xinput608 mprj_dat_o_core[4] vssd vssd vccd vccd net608 sky130_fd_sc_hd__buf_4
Xinput609 mprj_dat_o_core[5] vssd vssd vccd vccd net609 sky130_fd_sc_hd__clkbuf_4
Xinput61 la_data_out_core[36] vssd vssd vccd vccd net61 sky130_fd_sc_hd__clkbuf_4
Xinput610 mprj_dat_o_core[6] vssd vssd vccd vccd net610 sky130_fd_sc_hd__clkbuf_4
Xinput611 mprj_dat_o_core[7] vssd vssd vccd vccd net611 sky130_fd_sc_hd__buf_4
Xinput612 mprj_dat_o_core[8] vssd vssd vccd vccd net612 sky130_fd_sc_hd__buf_2
Xinput613 mprj_dat_o_core[9] vssd vssd vccd vccd net613 sky130_fd_sc_hd__clkbuf_4
Xinput614 mprj_iena_wb vssd vssd vccd vccd net614 sky130_fd_sc_hd__buf_2
Xinput615 mprj_sel_o_core[0] vssd vssd vccd vccd net615 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput616 mprj_sel_o_core[1] vssd vssd vccd vccd net616 sky130_fd_sc_hd__clkbuf_2
Xinput617 mprj_sel_o_core[2] vssd vssd vccd vccd net617 sky130_fd_sc_hd__clkbuf_2
Xinput618 mprj_sel_o_core[3] vssd vssd vccd vccd net618 sky130_fd_sc_hd__clkbuf_2
Xinput619 mprj_stb_o_core vssd vssd vccd vccd net619 sky130_fd_sc_hd__buf_4
Xinput62 la_data_out_core[37] vssd vssd vccd vccd net62 sky130_fd_sc_hd__clkbuf_4
Xinput620 mprj_we_o_core vssd vssd vccd vccd net620 sky130_fd_sc_hd__clkbuf_2
Xinput621 user_irq_core[0] vssd vssd vccd vccd net621 sky130_fd_sc_hd__clkbuf_1
Xinput622 user_irq_core[1] vssd vssd vccd vccd net622 sky130_fd_sc_hd__clkbuf_1
Xinput623 user_irq_core[2] vssd vssd vccd vccd net623 sky130_fd_sc_hd__clkbuf_1
Xinput624 user_irq_ena[0] vssd vssd vccd vccd net624 sky130_fd_sc_hd__clkbuf_1
Xinput625 user_irq_ena[1] vssd vssd vccd vccd net625 sky130_fd_sc_hd__clkbuf_1
Xinput626 user_irq_ena[2] vssd vssd vccd vccd net626 sky130_fd_sc_hd__clkbuf_1
Xinput63 la_data_out_core[38] vssd vssd vccd vccd net63 sky130_fd_sc_hd__clkbuf_4
Xinput64 la_data_out_core[39] vssd vssd vccd vccd net64 sky130_fd_sc_hd__clkbuf_4
Xinput65 la_data_out_core[3] vssd vssd vccd vccd net65 sky130_fd_sc_hd__clkbuf_4
Xinput66 la_data_out_core[40] vssd vssd vccd vccd net66 sky130_fd_sc_hd__clkbuf_4
Xinput67 la_data_out_core[41] vssd vssd vccd vccd net67 sky130_fd_sc_hd__buf_4
Xinput68 la_data_out_core[42] vssd vssd vccd vccd net68 sky130_fd_sc_hd__clkbuf_4
Xinput69 la_data_out_core[43] vssd vssd vccd vccd net69 sky130_fd_sc_hd__clkbuf_4
Xinput7 la_data_out_core[102] vssd vssd vccd vccd net7 sky130_fd_sc_hd__buf_4
Xinput70 la_data_out_core[44] vssd vssd vccd vccd net70 sky130_fd_sc_hd__clkbuf_4
Xinput71 la_data_out_core[45] vssd vssd vccd vccd net71 sky130_fd_sc_hd__buf_4
Xinput72 la_data_out_core[46] vssd vssd vccd vccd net72 sky130_fd_sc_hd__clkbuf_4
Xinput73 la_data_out_core[47] vssd vssd vccd vccd net73 sky130_fd_sc_hd__buf_4
Xinput74 la_data_out_core[48] vssd vssd vccd vccd net74 sky130_fd_sc_hd__buf_4
Xinput75 la_data_out_core[49] vssd vssd vccd vccd net75 sky130_fd_sc_hd__buf_4
Xinput76 la_data_out_core[4] vssd vssd vccd vccd net76 sky130_fd_sc_hd__clkbuf_4
Xinput77 la_data_out_core[50] vssd vssd vccd vccd net77 sky130_fd_sc_hd__buf_4
Xinput78 la_data_out_core[51] vssd vssd vccd vccd net78 sky130_fd_sc_hd__buf_4
Xinput79 la_data_out_core[52] vssd vssd vccd vccd net79 sky130_fd_sc_hd__buf_4
Xinput8 la_data_out_core[103] vssd vssd vccd vccd net8 sky130_fd_sc_hd__buf_4
Xinput80 la_data_out_core[53] vssd vssd vccd vccd net80 sky130_fd_sc_hd__buf_4
Xinput81 la_data_out_core[54] vssd vssd vccd vccd net81 sky130_fd_sc_hd__buf_4
Xinput82 la_data_out_core[55] vssd vssd vccd vccd net82 sky130_fd_sc_hd__buf_4
Xinput83 la_data_out_core[56] vssd vssd vccd vccd net83 sky130_fd_sc_hd__clkbuf_4
Xinput84 la_data_out_core[57] vssd vssd vccd vccd net84 sky130_fd_sc_hd__clkbuf_4
Xinput85 la_data_out_core[58] vssd vssd vccd vccd net85 sky130_fd_sc_hd__buf_4
Xinput86 la_data_out_core[59] vssd vssd vccd vccd net86 sky130_fd_sc_hd__buf_4
Xinput87 la_data_out_core[5] vssd vssd vccd vccd net87 sky130_fd_sc_hd__buf_2
Xinput88 la_data_out_core[60] vssd vssd vccd vccd net88 sky130_fd_sc_hd__clkbuf_4
Xinput89 la_data_out_core[61] vssd vssd vccd vccd net89 sky130_fd_sc_hd__buf_4
Xinput9 la_data_out_core[104] vssd vssd vccd vccd net9 sky130_fd_sc_hd__buf_4
Xinput90 la_data_out_core[62] vssd vssd vccd vccd net90 sky130_fd_sc_hd__buf_4
Xinput91 la_data_out_core[63] vssd vssd vccd vccd net91 sky130_fd_sc_hd__buf_4
Xinput92 la_data_out_core[64] vssd vssd vccd vccd net92 sky130_fd_sc_hd__buf_4
Xinput93 la_data_out_core[65] vssd vssd vccd vccd net93 sky130_fd_sc_hd__buf_4
Xinput94 la_data_out_core[66] vssd vssd vccd vccd net94 sky130_fd_sc_hd__clkbuf_4
Xinput95 la_data_out_core[67] vssd vssd vccd vccd net95 sky130_fd_sc_hd__clkbuf_4
Xinput96 la_data_out_core[68] vssd vssd vccd vccd net96 sky130_fd_sc_hd__clkbuf_4
Xinput97 la_data_out_core[69] vssd vssd vccd vccd net97 sky130_fd_sc_hd__buf_4
Xinput98 la_data_out_core[6] vssd vssd vccd vccd net98 sky130_fd_sc_hd__clkbuf_4
Xinput99 la_data_out_core[70] vssd vssd vccd vccd net99 sky130_fd_sc_hd__buf_4
X\la_buf[0]  _073_ \la_data_out_enable[0]\ vssd vssd vccd vccd la_data_in_core[0] sky130_fd_sc_hd__einvp_8
X\la_buf[100]  _074_ \la_data_out_enable[100]\ vssd vssd vccd vccd la_data_in_core[100] sky130_fd_sc_hd__einvp_8
X\la_buf[101]  _075_ \la_data_out_enable[101]\ vssd vssd vccd vccd la_data_in_core[101] sky130_fd_sc_hd__einvp_8
X\la_buf[102]  _076_ \la_data_out_enable[102]\ vssd vssd vccd vccd la_data_in_core[102] sky130_fd_sc_hd__einvp_8
X\la_buf[103]  _077_ \la_data_out_enable[103]\ vssd vssd vccd vccd la_data_in_core[103] sky130_fd_sc_hd__einvp_8
X\la_buf[104]  _078_ \la_data_out_enable[104]\ vssd vssd vccd vccd la_data_in_core[104] sky130_fd_sc_hd__einvp_8
X\la_buf[105]  _079_ \la_data_out_enable[105]\ vssd vssd vccd vccd la_data_in_core[105] sky130_fd_sc_hd__einvp_8
X\la_buf[106]  _080_ \la_data_out_enable[106]\ vssd vssd vccd vccd la_data_in_core[106] sky130_fd_sc_hd__einvp_8
X\la_buf[107]  _081_ \la_data_out_enable[107]\ vssd vssd vccd vccd la_data_in_core[107] sky130_fd_sc_hd__einvp_8
X\la_buf[108]  _082_ \la_data_out_enable[108]\ vssd vssd vccd vccd la_data_in_core[108] sky130_fd_sc_hd__einvp_8
X\la_buf[109]  _083_ \la_data_out_enable[109]\ vssd vssd vccd vccd la_data_in_core[109] sky130_fd_sc_hd__einvp_8
X\la_buf[10]  _084_ \la_data_out_enable[10]\ vssd vssd vccd vccd la_data_in_core[10] sky130_fd_sc_hd__einvp_8
X\la_buf[110]  _085_ \la_data_out_enable[110]\ vssd vssd vccd vccd la_data_in_core[110] sky130_fd_sc_hd__einvp_8
X\la_buf[111]  _086_ \la_data_out_enable[111]\ vssd vssd vccd vccd la_data_in_core[111] sky130_fd_sc_hd__einvp_8
X\la_buf[112]  _087_ \la_data_out_enable[112]\ vssd vssd vccd vccd la_data_in_core[112] sky130_fd_sc_hd__einvp_8
X\la_buf[113]  _088_ \la_data_out_enable[113]\ vssd vssd vccd vccd la_data_in_core[113] sky130_fd_sc_hd__einvp_8
X\la_buf[114]  _089_ \la_data_out_enable[114]\ vssd vssd vccd vccd la_data_in_core[114] sky130_fd_sc_hd__einvp_8
X\la_buf[115]  _090_ \la_data_out_enable[115]\ vssd vssd vccd vccd la_data_in_core[115] sky130_fd_sc_hd__einvp_8
X\la_buf[116]  _091_ \la_data_out_enable[116]\ vssd vssd vccd vccd la_data_in_core[116] sky130_fd_sc_hd__einvp_8
X\la_buf[117]  _092_ \la_data_out_enable[117]\ vssd vssd vccd vccd la_data_in_core[117] sky130_fd_sc_hd__einvp_8
X\la_buf[118]  _093_ \la_data_out_enable[118]\ vssd vssd vccd vccd la_data_in_core[118] sky130_fd_sc_hd__einvp_8
X\la_buf[119]  _094_ \la_data_out_enable[119]\ vssd vssd vccd vccd la_data_in_core[119] sky130_fd_sc_hd__einvp_8
X\la_buf[11]  _095_ \la_data_out_enable[11]\ vssd vssd vccd vccd la_data_in_core[11] sky130_fd_sc_hd__einvp_8
X\la_buf[120]  _096_ \la_data_out_enable[120]\ vssd vssd vccd vccd la_data_in_core[120] sky130_fd_sc_hd__einvp_8
X\la_buf[121]  _097_ \la_data_out_enable[121]\ vssd vssd vccd vccd la_data_in_core[121] sky130_fd_sc_hd__einvp_8
X\la_buf[122]  _098_ \la_data_out_enable[122]\ vssd vssd vccd vccd la_data_in_core[122] sky130_fd_sc_hd__einvp_8
X\la_buf[123]  _099_ \la_data_out_enable[123]\ vssd vssd vccd vccd la_data_in_core[123] sky130_fd_sc_hd__einvp_8
X\la_buf[124]  _100_ \la_data_out_enable[124]\ vssd vssd vccd vccd la_data_in_core[124] sky130_fd_sc_hd__einvp_8
X\la_buf[125]  _101_ \la_data_out_enable[125]\ vssd vssd vccd vccd la_data_in_core[125] sky130_fd_sc_hd__einvp_8
X\la_buf[126]  _102_ \la_data_out_enable[126]\ vssd vssd vccd vccd la_data_in_core[126] sky130_fd_sc_hd__einvp_8
X\la_buf[127]  _103_ \la_data_out_enable[127]\ vssd vssd vccd vccd la_data_in_core[127] sky130_fd_sc_hd__einvp_8
X\la_buf[12]  _104_ \la_data_out_enable[12]\ vssd vssd vccd vccd la_data_in_core[12] sky130_fd_sc_hd__einvp_8
X\la_buf[13]  _105_ \la_data_out_enable[13]\ vssd vssd vccd vccd la_data_in_core[13] sky130_fd_sc_hd__einvp_8
X\la_buf[14]  _106_ \la_data_out_enable[14]\ vssd vssd vccd vccd la_data_in_core[14] sky130_fd_sc_hd__einvp_8
X\la_buf[15]  _107_ \la_data_out_enable[15]\ vssd vssd vccd vccd la_data_in_core[15] sky130_fd_sc_hd__einvp_8
X\la_buf[16]  _108_ \la_data_out_enable[16]\ vssd vssd vccd vccd la_data_in_core[16] sky130_fd_sc_hd__einvp_8
X\la_buf[17]  _109_ \la_data_out_enable[17]\ vssd vssd vccd vccd la_data_in_core[17] sky130_fd_sc_hd__einvp_8
X\la_buf[18]  _110_ \la_data_out_enable[18]\ vssd vssd vccd vccd la_data_in_core[18] sky130_fd_sc_hd__einvp_8
X\la_buf[19]  _111_ \la_data_out_enable[19]\ vssd vssd vccd vccd la_data_in_core[19] sky130_fd_sc_hd__einvp_8
X\la_buf[1]  _112_ \la_data_out_enable[1]\ vssd vssd vccd vccd la_data_in_core[1] sky130_fd_sc_hd__einvp_8
X\la_buf[20]  _113_ \la_data_out_enable[20]\ vssd vssd vccd vccd la_data_in_core[20] sky130_fd_sc_hd__einvp_8
X\la_buf[21]  _114_ \la_data_out_enable[21]\ vssd vssd vccd vccd la_data_in_core[21] sky130_fd_sc_hd__einvp_8
X\la_buf[22]  _115_ \la_data_out_enable[22]\ vssd vssd vccd vccd la_data_in_core[22] sky130_fd_sc_hd__einvp_8
X\la_buf[23]  _116_ \la_data_out_enable[23]\ vssd vssd vccd vccd la_data_in_core[23] sky130_fd_sc_hd__einvp_8
X\la_buf[24]  _117_ \la_data_out_enable[24]\ vssd vssd vccd vccd la_data_in_core[24] sky130_fd_sc_hd__einvp_8
X\la_buf[25]  _118_ \la_data_out_enable[25]\ vssd vssd vccd vccd la_data_in_core[25] sky130_fd_sc_hd__einvp_8
X\la_buf[26]  _119_ \la_data_out_enable[26]\ vssd vssd vccd vccd la_data_in_core[26] sky130_fd_sc_hd__einvp_8
X\la_buf[27]  _120_ \la_data_out_enable[27]\ vssd vssd vccd vccd la_data_in_core[27] sky130_fd_sc_hd__einvp_8
X\la_buf[28]  _121_ \la_data_out_enable[28]\ vssd vssd vccd vccd la_data_in_core[28] sky130_fd_sc_hd__einvp_8
X\la_buf[29]  _122_ \la_data_out_enable[29]\ vssd vssd vccd vccd la_data_in_core[29] sky130_fd_sc_hd__einvp_8
X\la_buf[2]  _123_ \la_data_out_enable[2]\ vssd vssd vccd vccd la_data_in_core[2] sky130_fd_sc_hd__einvp_8
X\la_buf[30]  _124_ \la_data_out_enable[30]\ vssd vssd vccd vccd la_data_in_core[30] sky130_fd_sc_hd__einvp_8
X\la_buf[31]  _125_ \la_data_out_enable[31]\ vssd vssd vccd vccd la_data_in_core[31] sky130_fd_sc_hd__einvp_8
X\la_buf[32]  _126_ \la_data_out_enable[32]\ vssd vssd vccd vccd la_data_in_core[32] sky130_fd_sc_hd__einvp_8
X\la_buf[33]  _127_ \la_data_out_enable[33]\ vssd vssd vccd vccd la_data_in_core[33] sky130_fd_sc_hd__einvp_8
X\la_buf[34]  _128_ \la_data_out_enable[34]\ vssd vssd vccd vccd la_data_in_core[34] sky130_fd_sc_hd__einvp_8
X\la_buf[35]  _129_ \la_data_out_enable[35]\ vssd vssd vccd vccd la_data_in_core[35] sky130_fd_sc_hd__einvp_8
X\la_buf[36]  _130_ \la_data_out_enable[36]\ vssd vssd vccd vccd la_data_in_core[36] sky130_fd_sc_hd__einvp_8
X\la_buf[37]  _131_ \la_data_out_enable[37]\ vssd vssd vccd vccd la_data_in_core[37] sky130_fd_sc_hd__einvp_8
X\la_buf[38]  _132_ \la_data_out_enable[38]\ vssd vssd vccd vccd la_data_in_core[38] sky130_fd_sc_hd__einvp_8
X\la_buf[39]  _133_ \la_data_out_enable[39]\ vssd vssd vccd vccd la_data_in_core[39] sky130_fd_sc_hd__einvp_8
X\la_buf[3]  _134_ \la_data_out_enable[3]\ vssd vssd vccd vccd la_data_in_core[3] sky130_fd_sc_hd__einvp_8
X\la_buf[40]  _135_ \la_data_out_enable[40]\ vssd vssd vccd vccd la_data_in_core[40] sky130_fd_sc_hd__einvp_8
X\la_buf[41]  _136_ \la_data_out_enable[41]\ vssd vssd vccd vccd la_data_in_core[41] sky130_fd_sc_hd__einvp_8
X\la_buf[42]  _137_ \la_data_out_enable[42]\ vssd vssd vccd vccd la_data_in_core[42] sky130_fd_sc_hd__einvp_8
X\la_buf[43]  _138_ \la_data_out_enable[43]\ vssd vssd vccd vccd la_data_in_core[43] sky130_fd_sc_hd__einvp_8
X\la_buf[44]  _139_ \la_data_out_enable[44]\ vssd vssd vccd vccd la_data_in_core[44] sky130_fd_sc_hd__einvp_8
X\la_buf[45]  _140_ \la_data_out_enable[45]\ vssd vssd vccd vccd la_data_in_core[45] sky130_fd_sc_hd__einvp_8
X\la_buf[46]  _141_ \la_data_out_enable[46]\ vssd vssd vccd vccd la_data_in_core[46] sky130_fd_sc_hd__einvp_8
X\la_buf[47]  _142_ \la_data_out_enable[47]\ vssd vssd vccd vccd la_data_in_core[47] sky130_fd_sc_hd__einvp_8
X\la_buf[48]  _143_ \la_data_out_enable[48]\ vssd vssd vccd vccd la_data_in_core[48] sky130_fd_sc_hd__einvp_8
X\la_buf[49]  _144_ \la_data_out_enable[49]\ vssd vssd vccd vccd la_data_in_core[49] sky130_fd_sc_hd__einvp_8
X\la_buf[4]  _145_ \la_data_out_enable[4]\ vssd vssd vccd vccd la_data_in_core[4] sky130_fd_sc_hd__einvp_8
X\la_buf[50]  _146_ \la_data_out_enable[50]\ vssd vssd vccd vccd la_data_in_core[50] sky130_fd_sc_hd__einvp_8
X\la_buf[51]  _147_ \la_data_out_enable[51]\ vssd vssd vccd vccd la_data_in_core[51] sky130_fd_sc_hd__einvp_8
X\la_buf[52]  _148_ \la_data_out_enable[52]\ vssd vssd vccd vccd la_data_in_core[52] sky130_fd_sc_hd__einvp_8
X\la_buf[53]  _149_ \la_data_out_enable[53]\ vssd vssd vccd vccd la_data_in_core[53] sky130_fd_sc_hd__einvp_8
X\la_buf[54]  _150_ \la_data_out_enable[54]\ vssd vssd vccd vccd la_data_in_core[54] sky130_fd_sc_hd__einvp_8
X\la_buf[55]  _151_ \la_data_out_enable[55]\ vssd vssd vccd vccd la_data_in_core[55] sky130_fd_sc_hd__einvp_8
X\la_buf[56]  _152_ \la_data_out_enable[56]\ vssd vssd vccd vccd la_data_in_core[56] sky130_fd_sc_hd__einvp_8
X\la_buf[57]  _153_ \la_data_out_enable[57]\ vssd vssd vccd vccd la_data_in_core[57] sky130_fd_sc_hd__einvp_8
X\la_buf[58]  _154_ \la_data_out_enable[58]\ vssd vssd vccd vccd la_data_in_core[58] sky130_fd_sc_hd__einvp_8
X\la_buf[59]  _155_ \la_data_out_enable[59]\ vssd vssd vccd vccd la_data_in_core[59] sky130_fd_sc_hd__einvp_8
X\la_buf[5]  _156_ \la_data_out_enable[5]\ vssd vssd vccd vccd la_data_in_core[5] sky130_fd_sc_hd__einvp_8
X\la_buf[60]  _157_ \la_data_out_enable[60]\ vssd vssd vccd vccd la_data_in_core[60] sky130_fd_sc_hd__einvp_8
X\la_buf[61]  _158_ \la_data_out_enable[61]\ vssd vssd vccd vccd la_data_in_core[61] sky130_fd_sc_hd__einvp_8
X\la_buf[62]  _159_ \la_data_out_enable[62]\ vssd vssd vccd vccd la_data_in_core[62] sky130_fd_sc_hd__einvp_8
X\la_buf[63]  _160_ \la_data_out_enable[63]\ vssd vssd vccd vccd la_data_in_core[63] sky130_fd_sc_hd__einvp_8
X\la_buf[64]  _161_ \la_data_out_enable[64]\ vssd vssd vccd vccd la_data_in_core[64] sky130_fd_sc_hd__einvp_8
X\la_buf[65]  _162_ \la_data_out_enable[65]\ vssd vssd vccd vccd la_data_in_core[65] sky130_fd_sc_hd__einvp_8
X\la_buf[66]  _163_ \la_data_out_enable[66]\ vssd vssd vccd vccd la_data_in_core[66] sky130_fd_sc_hd__einvp_8
X\la_buf[67]  _164_ \la_data_out_enable[67]\ vssd vssd vccd vccd la_data_in_core[67] sky130_fd_sc_hd__einvp_8
X\la_buf[68]  _165_ \la_data_out_enable[68]\ vssd vssd vccd vccd la_data_in_core[68] sky130_fd_sc_hd__einvp_8
X\la_buf[69]  _166_ \la_data_out_enable[69]\ vssd vssd vccd vccd la_data_in_core[69] sky130_fd_sc_hd__einvp_8
X\la_buf[6]  _167_ \la_data_out_enable[6]\ vssd vssd vccd vccd la_data_in_core[6] sky130_fd_sc_hd__einvp_8
X\la_buf[70]  _168_ \la_data_out_enable[70]\ vssd vssd vccd vccd la_data_in_core[70] sky130_fd_sc_hd__einvp_8
X\la_buf[71]  _169_ \la_data_out_enable[71]\ vssd vssd vccd vccd la_data_in_core[71] sky130_fd_sc_hd__einvp_8
X\la_buf[72]  _170_ \la_data_out_enable[72]\ vssd vssd vccd vccd la_data_in_core[72] sky130_fd_sc_hd__einvp_8
X\la_buf[73]  _171_ \la_data_out_enable[73]\ vssd vssd vccd vccd la_data_in_core[73] sky130_fd_sc_hd__einvp_8
X\la_buf[74]  _172_ \la_data_out_enable[74]\ vssd vssd vccd vccd la_data_in_core[74] sky130_fd_sc_hd__einvp_8
X\la_buf[75]  _173_ \la_data_out_enable[75]\ vssd vssd vccd vccd la_data_in_core[75] sky130_fd_sc_hd__einvp_8
X\la_buf[76]  _174_ \la_data_out_enable[76]\ vssd vssd vccd vccd la_data_in_core[76] sky130_fd_sc_hd__einvp_8
X\la_buf[77]  _175_ \la_data_out_enable[77]\ vssd vssd vccd vccd la_data_in_core[77] sky130_fd_sc_hd__einvp_8
X\la_buf[78]  _176_ \la_data_out_enable[78]\ vssd vssd vccd vccd la_data_in_core[78] sky130_fd_sc_hd__einvp_8
X\la_buf[79]  _177_ \la_data_out_enable[79]\ vssd vssd vccd vccd la_data_in_core[79] sky130_fd_sc_hd__einvp_8
X\la_buf[7]  _178_ \la_data_out_enable[7]\ vssd vssd vccd vccd la_data_in_core[7] sky130_fd_sc_hd__einvp_8
X\la_buf[80]  _179_ \la_data_out_enable[80]\ vssd vssd vccd vccd la_data_in_core[80] sky130_fd_sc_hd__einvp_8
X\la_buf[81]  _180_ \la_data_out_enable[81]\ vssd vssd vccd vccd la_data_in_core[81] sky130_fd_sc_hd__einvp_8
X\la_buf[82]  _181_ \la_data_out_enable[82]\ vssd vssd vccd vccd la_data_in_core[82] sky130_fd_sc_hd__einvp_8
X\la_buf[83]  _182_ \la_data_out_enable[83]\ vssd vssd vccd vccd la_data_in_core[83] sky130_fd_sc_hd__einvp_8
X\la_buf[84]  _183_ \la_data_out_enable[84]\ vssd vssd vccd vccd la_data_in_core[84] sky130_fd_sc_hd__einvp_8
X\la_buf[85]  _184_ \la_data_out_enable[85]\ vssd vssd vccd vccd la_data_in_core[85] sky130_fd_sc_hd__einvp_8
X\la_buf[86]  _185_ \la_data_out_enable[86]\ vssd vssd vccd vccd la_data_in_core[86] sky130_fd_sc_hd__einvp_8
X\la_buf[87]  _186_ \la_data_out_enable[87]\ vssd vssd vccd vccd la_data_in_core[87] sky130_fd_sc_hd__einvp_8
X\la_buf[88]  _187_ \la_data_out_enable[88]\ vssd vssd vccd vccd la_data_in_core[88] sky130_fd_sc_hd__einvp_8
X\la_buf[89]  _188_ \la_data_out_enable[89]\ vssd vssd vccd vccd la_data_in_core[89] sky130_fd_sc_hd__einvp_8
X\la_buf[8]  _189_ \la_data_out_enable[8]\ vssd vssd vccd vccd la_data_in_core[8] sky130_fd_sc_hd__einvp_8
X\la_buf[90]  _190_ \la_data_out_enable[90]\ vssd vssd vccd vccd la_data_in_core[90] sky130_fd_sc_hd__einvp_8
X\la_buf[91]  _191_ \la_data_out_enable[91]\ vssd vssd vccd vccd la_data_in_core[91] sky130_fd_sc_hd__einvp_8
X\la_buf[92]  _192_ \la_data_out_enable[92]\ vssd vssd vccd vccd la_data_in_core[92] sky130_fd_sc_hd__einvp_8
X\la_buf[93]  _193_ \la_data_out_enable[93]\ vssd vssd vccd vccd la_data_in_core[93] sky130_fd_sc_hd__einvp_8
X\la_buf[94]  _194_ \la_data_out_enable[94]\ vssd vssd vccd vccd la_data_in_core[94] sky130_fd_sc_hd__einvp_8
X\la_buf[95]  _195_ \la_data_out_enable[95]\ vssd vssd vccd vccd la_data_in_core[95] sky130_fd_sc_hd__einvp_8
X\la_buf[96]  _196_ \la_data_out_enable[96]\ vssd vssd vccd vccd la_data_in_core[96] sky130_fd_sc_hd__einvp_8
X\la_buf[97]  _197_ \la_data_out_enable[97]\ vssd vssd vccd vccd la_data_in_core[97] sky130_fd_sc_hd__einvp_8
X\la_buf[98]  _198_ \la_data_out_enable[98]\ vssd vssd vccd vccd la_data_in_core[98] sky130_fd_sc_hd__einvp_8
X\la_buf[99]  _199_ \la_data_out_enable[99]\ vssd vssd vccd vccd la_data_in_core[99] sky130_fd_sc_hd__einvp_8
X\la_buf[9]  _200_ \la_data_out_enable[9]\ vssd vssd vccd vccd la_data_in_core[9] sky130_fd_sc_hd__einvp_8
X\la_buf_enable[0]  net388 \mprj_logic1[74]\ vssd vssd vccd vccd \la_data_out_enable[0]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[100]  net389 \mprj_logic1[174]\ vssd vssd vccd vccd \la_data_out_enable[100]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[101]  net390 \mprj_logic1[175]\ vssd vssd vccd vccd \la_data_out_enable[101]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[102]  net391 \mprj_logic1[176]\ vssd vssd vccd vccd \la_data_out_enable[102]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[103]  net392 \mprj_logic1[177]\ vssd vssd vccd vccd \la_data_out_enable[103]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[104]  net393 \mprj_logic1[178]\ vssd vssd vccd vccd \la_data_out_enable[104]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[105]  net394 \mprj_logic1[179]\ vssd vssd vccd vccd \la_data_out_enable[105]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[106]  net395 \mprj_logic1[180]\ vssd vssd vccd vccd \la_data_out_enable[106]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[107]  net396 \mprj_logic1[181]\ vssd vssd vccd vccd \la_data_out_enable[107]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[108]  net397 \mprj_logic1[182]\ vssd vssd vccd vccd \la_data_out_enable[108]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[109]  net398 \mprj_logic1[183]\ vssd vssd vccd vccd \la_data_out_enable[109]\ sky130_fd_sc_hd__and2b_2
X\la_buf_enable[10]  net399 \mprj_logic1[84]\ vssd vssd vccd vccd \la_data_out_enable[10]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[110]  net400 \mprj_logic1[184]\ vssd vssd vccd vccd \la_data_out_enable[110]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[111]  net401 \mprj_logic1[185]\ vssd vssd vccd vccd \la_data_out_enable[111]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[112]  net402 \mprj_logic1[186]\ vssd vssd vccd vccd \la_data_out_enable[112]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[113]  net403 \mprj_logic1[187]\ vssd vssd vccd vccd \la_data_out_enable[113]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[114]  net404 \mprj_logic1[188]\ vssd vssd vccd vccd \la_data_out_enable[114]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[115]  net405 \mprj_logic1[189]\ vssd vssd vccd vccd \la_data_out_enable[115]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[116]  net406 \mprj_logic1[190]\ vssd vssd vccd vccd \la_data_out_enable[116]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[117]  net407 \mprj_logic1[191]\ vssd vssd vccd vccd \la_data_out_enable[117]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[118]  net408 \mprj_logic1[192]\ vssd vssd vccd vccd \la_data_out_enable[118]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[119]  net409 \mprj_logic1[193]\ vssd vssd vccd vccd \la_data_out_enable[119]\ sky130_fd_sc_hd__and2b_2
X\la_buf_enable[11]  net410 \mprj_logic1[85]\ vssd vssd vccd vccd \la_data_out_enable[11]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[120]  net411 \mprj_logic1[194]\ vssd vssd vccd vccd \la_data_out_enable[120]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[121]  net412 \mprj_logic1[195]\ vssd vssd vccd vccd \la_data_out_enable[121]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[122]  net413 \mprj_logic1[196]\ vssd vssd vccd vccd \la_data_out_enable[122]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[123]  net414 \mprj_logic1[197]\ vssd vssd vccd vccd \la_data_out_enable[123]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[124]  net415 \mprj_logic1[198]\ vssd vssd vccd vccd \la_data_out_enable[124]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[125]  net416 \mprj_logic1[199]\ vssd vssd vccd vccd \la_data_out_enable[125]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[126]  net417 \mprj_logic1[200]\ vssd vssd vccd vccd \la_data_out_enable[126]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[127]  net418 \mprj_logic1[201]\ vssd vssd vccd vccd \la_data_out_enable[127]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[12]  net419 \mprj_logic1[86]\ vssd vssd vccd vccd \la_data_out_enable[12]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[13]  net420 \mprj_logic1[87]\ vssd vssd vccd vccd \la_data_out_enable[13]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[14]  net421 \mprj_logic1[88]\ vssd vssd vccd vccd \la_data_out_enable[14]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[15]  net422 \mprj_logic1[89]\ vssd vssd vccd vccd \la_data_out_enable[15]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[16]  net423 \mprj_logic1[90]\ vssd vssd vccd vccd \la_data_out_enable[16]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[17]  net424 \mprj_logic1[91]\ vssd vssd vccd vccd \la_data_out_enable[17]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[18]  net425 \mprj_logic1[92]\ vssd vssd vccd vccd \la_data_out_enable[18]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[19]  net426 \mprj_logic1[93]\ vssd vssd vccd vccd \la_data_out_enable[19]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[1]  net427 \mprj_logic1[75]\ vssd vssd vccd vccd \la_data_out_enable[1]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[20]  net428 \mprj_logic1[94]\ vssd vssd vccd vccd \la_data_out_enable[20]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[21]  net429 \mprj_logic1[95]\ vssd vssd vccd vccd \la_data_out_enable[21]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[22]  net430 \mprj_logic1[96]\ vssd vssd vccd vccd \la_data_out_enable[22]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[23]  net431 \mprj_logic1[97]\ vssd vssd vccd vccd \la_data_out_enable[23]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[24]  net432 \mprj_logic1[98]\ vssd vssd vccd vccd \la_data_out_enable[24]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[25]  net433 \mprj_logic1[99]\ vssd vssd vccd vccd \la_data_out_enable[25]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[26]  net434 \mprj_logic1[100]\ vssd vssd vccd vccd \la_data_out_enable[26]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[27]  net435 \mprj_logic1[101]\ vssd vssd vccd vccd \la_data_out_enable[27]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[28]  net436 \mprj_logic1[102]\ vssd vssd vccd vccd \la_data_out_enable[28]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[29]  net437 \mprj_logic1[103]\ vssd vssd vccd vccd \la_data_out_enable[29]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[2]  net438 \mprj_logic1[76]\ vssd vssd vccd vccd \la_data_out_enable[2]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[30]  net439 \mprj_logic1[104]\ vssd vssd vccd vccd \la_data_out_enable[30]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[31]  net440 \mprj_logic1[105]\ vssd vssd vccd vccd \la_data_out_enable[31]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[32]  net441 \mprj_logic1[106]\ vssd vssd vccd vccd \la_data_out_enable[32]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[33]  net442 \mprj_logic1[107]\ vssd vssd vccd vccd \la_data_out_enable[33]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[34]  net443 \mprj_logic1[108]\ vssd vssd vccd vccd \la_data_out_enable[34]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[35]  net444 \mprj_logic1[109]\ vssd vssd vccd vccd \la_data_out_enable[35]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[36]  net445 \mprj_logic1[110]\ vssd vssd vccd vccd \la_data_out_enable[36]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[37]  net446 \mprj_logic1[111]\ vssd vssd vccd vccd \la_data_out_enable[37]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[38]  net447 \mprj_logic1[112]\ vssd vssd vccd vccd \la_data_out_enable[38]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[39]  net448 \mprj_logic1[113]\ vssd vssd vccd vccd \la_data_out_enable[39]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[3]  net449 \mprj_logic1[77]\ vssd vssd vccd vccd \la_data_out_enable[3]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[40]  net450 \mprj_logic1[114]\ vssd vssd vccd vccd \la_data_out_enable[40]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[41]  net451 \mprj_logic1[115]\ vssd vssd vccd vccd \la_data_out_enable[41]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[42]  net452 \mprj_logic1[116]\ vssd vssd vccd vccd \la_data_out_enable[42]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[43]  net453 \mprj_logic1[117]\ vssd vssd vccd vccd \la_data_out_enable[43]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[44]  net454 \mprj_logic1[118]\ vssd vssd vccd vccd \la_data_out_enable[44]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[45]  net455 \mprj_logic1[119]\ vssd vssd vccd vccd \la_data_out_enable[45]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[46]  net456 \mprj_logic1[120]\ vssd vssd vccd vccd \la_data_out_enable[46]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[47]  net457 \mprj_logic1[121]\ vssd vssd vccd vccd \la_data_out_enable[47]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[48]  net458 \mprj_logic1[122]\ vssd vssd vccd vccd \la_data_out_enable[48]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[49]  net459 \mprj_logic1[123]\ vssd vssd vccd vccd \la_data_out_enable[49]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[4]  net460 \mprj_logic1[78]\ vssd vssd vccd vccd \la_data_out_enable[4]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[50]  net461 \mprj_logic1[124]\ vssd vssd vccd vccd \la_data_out_enable[50]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[51]  net462 \mprj_logic1[125]\ vssd vssd vccd vccd \la_data_out_enable[51]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[52]  net463 \mprj_logic1[126]\ vssd vssd vccd vccd \la_data_out_enable[52]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[53]  net464 \mprj_logic1[127]\ vssd vssd vccd vccd \la_data_out_enable[53]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[54]  net465 \mprj_logic1[128]\ vssd vssd vccd vccd \la_data_out_enable[54]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[55]  net466 \mprj_logic1[129]\ vssd vssd vccd vccd \la_data_out_enable[55]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[56]  net467 \mprj_logic1[130]\ vssd vssd vccd vccd \la_data_out_enable[56]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[57]  net468 \mprj_logic1[131]\ vssd vssd vccd vccd \la_data_out_enable[57]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[58]  net469 \mprj_logic1[132]\ vssd vssd vccd vccd \la_data_out_enable[58]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[59]  net470 \mprj_logic1[133]\ vssd vssd vccd vccd \la_data_out_enable[59]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[5]  net471 \mprj_logic1[79]\ vssd vssd vccd vccd \la_data_out_enable[5]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[60]  net472 \mprj_logic1[134]\ vssd vssd vccd vccd \la_data_out_enable[60]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[61]  net473 \mprj_logic1[135]\ vssd vssd vccd vccd \la_data_out_enable[61]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[62]  net474 \mprj_logic1[136]\ vssd vssd vccd vccd \la_data_out_enable[62]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[63]  net475 \mprj_logic1[137]\ vssd vssd vccd vccd \la_data_out_enable[63]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[64]  net476 \mprj_logic1[138]\ vssd vssd vccd vccd \la_data_out_enable[64]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[65]  net477 \mprj_logic1[139]\ vssd vssd vccd vccd \la_data_out_enable[65]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[66]  net478 \mprj_logic1[140]\ vssd vssd vccd vccd \la_data_out_enable[66]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[67]  net479 \mprj_logic1[141]\ vssd vssd vccd vccd \la_data_out_enable[67]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[68]  net480 \mprj_logic1[142]\ vssd vssd vccd vccd \la_data_out_enable[68]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[69]  net481 \mprj_logic1[143]\ vssd vssd vccd vccd \la_data_out_enable[69]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[6]  net482 \mprj_logic1[80]\ vssd vssd vccd vccd \la_data_out_enable[6]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[70]  net483 \mprj_logic1[144]\ vssd vssd vccd vccd \la_data_out_enable[70]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[71]  net484 \mprj_logic1[145]\ vssd vssd vccd vccd \la_data_out_enable[71]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[72]  net485 \mprj_logic1[146]\ vssd vssd vccd vccd \la_data_out_enable[72]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[73]  net486 \mprj_logic1[147]\ vssd vssd vccd vccd \la_data_out_enable[73]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[74]  net487 \mprj_logic1[148]\ vssd vssd vccd vccd \la_data_out_enable[74]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[75]  net488 \mprj_logic1[149]\ vssd vssd vccd vccd \la_data_out_enable[75]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[76]  net489 \mprj_logic1[150]\ vssd vssd vccd vccd \la_data_out_enable[76]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[77]  net490 \mprj_logic1[151]\ vssd vssd vccd vccd \la_data_out_enable[77]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[78]  net491 \mprj_logic1[152]\ vssd vssd vccd vccd \la_data_out_enable[78]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[79]  net492 \mprj_logic1[153]\ vssd vssd vccd vccd \la_data_out_enable[79]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[7]  net493 \mprj_logic1[81]\ vssd vssd vccd vccd \la_data_out_enable[7]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[80]  net494 \mprj_logic1[154]\ vssd vssd vccd vccd \la_data_out_enable[80]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[81]  net495 \mprj_logic1[155]\ vssd vssd vccd vccd \la_data_out_enable[81]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[82]  net496 \mprj_logic1[156]\ vssd vssd vccd vccd \la_data_out_enable[82]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[83]  net497 \mprj_logic1[157]\ vssd vssd vccd vccd \la_data_out_enable[83]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[84]  net498 \mprj_logic1[158]\ vssd vssd vccd vccd \la_data_out_enable[84]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[85]  net499 \mprj_logic1[159]\ vssd vssd vccd vccd \la_data_out_enable[85]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[86]  net500 \mprj_logic1[160]\ vssd vssd vccd vccd \la_data_out_enable[86]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[87]  net501 \mprj_logic1[161]\ vssd vssd vccd vccd \la_data_out_enable[87]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[88]  net502 \mprj_logic1[162]\ vssd vssd vccd vccd \la_data_out_enable[88]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[89]  net503 \mprj_logic1[163]\ vssd vssd vccd vccd \la_data_out_enable[89]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[8]  net504 \mprj_logic1[82]\ vssd vssd vccd vccd \la_data_out_enable[8]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[90]  net505 \mprj_logic1[164]\ vssd vssd vccd vccd \la_data_out_enable[90]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[91]  net506 \mprj_logic1[165]\ vssd vssd vccd vccd \la_data_out_enable[91]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[92]  net507 \mprj_logic1[166]\ vssd vssd vccd vccd \la_data_out_enable[92]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[93]  net508 \mprj_logic1[167]\ vssd vssd vccd vccd \la_data_out_enable[93]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[94]  net509 \mprj_logic1[168]\ vssd vssd vccd vccd \la_data_out_enable[94]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[95]  net510 \mprj_logic1[169]\ vssd vssd vccd vccd \la_data_out_enable[95]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[96]  net511 \mprj_logic1[170]\ vssd vssd vccd vccd \la_data_out_enable[96]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[97]  net512 \mprj_logic1[171]\ vssd vssd vccd vccd \la_data_out_enable[97]\ sky130_fd_sc_hd__and2b_2
X\la_buf_enable[98]  net513 \mprj_logic1[172]\ vssd vssd vccd vccd \la_data_out_enable[98]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[99]  net514 \mprj_logic1[173]\ vssd vssd vccd vccd \la_data_out_enable[99]\ sky130_fd_sc_hd__and2b_1
X\la_buf_enable[9]  net515 \mprj_logic1[83]\ vssd vssd vccd vccd \la_data_out_enable[9]\ sky130_fd_sc_hd__and2b_1
Xmprj2_logic_high_inst mprj2_logic1 vccd2 vssd2 mprj2_logic_high
Xmprj2_pwrgood mprj2_logic1 vssd vssd vccd vccd net790 sky130_fd_sc_hd__buf_12
Xmprj2_vdd_pwrgood mprj2_vdd_logic1 vssd vssd vccd vccd net791 sky130_fd_sc_hd__buf_6
X\mprj_adr_buf[0]  _009_ \mprj_logic1[10]\ vssd vssd vccd vccd mprj_adr_o_user[0] sky130_fd_sc_hd__einvp_8
X\mprj_adr_buf[10]  _010_ \mprj_logic1[20]\ vssd vssd vccd vccd mprj_adr_o_user[10] sky130_fd_sc_hd__einvp_8
X\mprj_adr_buf[11]  _011_ \mprj_logic1[21]\ vssd vssd vccd vccd mprj_adr_o_user[11] sky130_fd_sc_hd__einvp_8
X\mprj_adr_buf[12]  _012_ \mprj_logic1[22]\ vssd vssd vccd vccd mprj_adr_o_user[12] sky130_fd_sc_hd__einvp_8
X\mprj_adr_buf[13]  _013_ \mprj_logic1[23]\ vssd vssd vccd vccd mprj_adr_o_user[13] sky130_fd_sc_hd__einvp_8
X\mprj_adr_buf[14]  _014_ \mprj_logic1[24]\ vssd vssd vccd vccd mprj_adr_o_user[14] sky130_fd_sc_hd__einvp_8
X\mprj_adr_buf[15]  _015_ \mprj_logic1[25]\ vssd vssd vccd vccd mprj_adr_o_user[15] sky130_fd_sc_hd__einvp_8
X\mprj_adr_buf[16]  _016_ \mprj_logic1[26]\ vssd vssd vccd vccd mprj_adr_o_user[16] sky130_fd_sc_hd__einvp_8
X\mprj_adr_buf[17]  _017_ \mprj_logic1[27]\ vssd vssd vccd vccd mprj_adr_o_user[17] sky130_fd_sc_hd__einvp_8
X\mprj_adr_buf[18]  _018_ \mprj_logic1[28]\ vssd vssd vccd vccd mprj_adr_o_user[18] sky130_fd_sc_hd__einvp_8
X\mprj_adr_buf[19]  _019_ \mprj_logic1[29]\ vssd vssd vccd vccd mprj_adr_o_user[19] sky130_fd_sc_hd__einvp_8
X\mprj_adr_buf[1]  _020_ \mprj_logic1[11]\ vssd vssd vccd vccd mprj_adr_o_user[1] sky130_fd_sc_hd__einvp_8
X\mprj_adr_buf[20]  _021_ \mprj_logic1[30]\ vssd vssd vccd vccd mprj_adr_o_user[20] sky130_fd_sc_hd__einvp_8
X\mprj_adr_buf[21]  _022_ \mprj_logic1[31]\ vssd vssd vccd vccd mprj_adr_o_user[21] sky130_fd_sc_hd__einvp_8
X\mprj_adr_buf[22]  _023_ \mprj_logic1[32]\ vssd vssd vccd vccd mprj_adr_o_user[22] sky130_fd_sc_hd__einvp_8
X\mprj_adr_buf[23]  _024_ \mprj_logic1[33]\ vssd vssd vccd vccd mprj_adr_o_user[23] sky130_fd_sc_hd__einvp_8
X\mprj_adr_buf[24]  _025_ \mprj_logic1[34]\ vssd vssd vccd vccd mprj_adr_o_user[24] sky130_fd_sc_hd__einvp_8
X\mprj_adr_buf[25]  _026_ \mprj_logic1[35]\ vssd vssd vccd vccd mprj_adr_o_user[25] sky130_fd_sc_hd__einvp_8
X\mprj_adr_buf[26]  _027_ \mprj_logic1[36]\ vssd vssd vccd vccd mprj_adr_o_user[26] sky130_fd_sc_hd__einvp_8
X\mprj_adr_buf[27]  _028_ \mprj_logic1[37]\ vssd vssd vccd vccd mprj_adr_o_user[27] sky130_fd_sc_hd__einvp_8
X\mprj_adr_buf[28]  _029_ \mprj_logic1[38]\ vssd vssd vccd vccd mprj_adr_o_user[28] sky130_fd_sc_hd__einvp_8
X\mprj_adr_buf[29]  _030_ \mprj_logic1[39]\ vssd vssd vccd vccd mprj_adr_o_user[29] sky130_fd_sc_hd__einvp_8
X\mprj_adr_buf[2]  _031_ \mprj_logic1[12]\ vssd vssd vccd vccd mprj_adr_o_user[2] sky130_fd_sc_hd__einvp_8
X\mprj_adr_buf[30]  _032_ \mprj_logic1[40]\ vssd vssd vccd vccd mprj_adr_o_user[30] sky130_fd_sc_hd__einvp_8
X\mprj_adr_buf[31]  _033_ \mprj_logic1[41]\ vssd vssd vccd vccd mprj_adr_o_user[31] sky130_fd_sc_hd__einvp_8
X\mprj_adr_buf[3]  _034_ \mprj_logic1[13]\ vssd vssd vccd vccd mprj_adr_o_user[3] sky130_fd_sc_hd__einvp_8
X\mprj_adr_buf[4]  _035_ \mprj_logic1[14]\ vssd vssd vccd vccd mprj_adr_o_user[4] sky130_fd_sc_hd__einvp_8
X\mprj_adr_buf[5]  _036_ \mprj_logic1[15]\ vssd vssd vccd vccd mprj_adr_o_user[5] sky130_fd_sc_hd__einvp_8
X\mprj_adr_buf[6]  _037_ \mprj_logic1[16]\ vssd vssd vccd vccd mprj_adr_o_user[6] sky130_fd_sc_hd__einvp_8
X\mprj_adr_buf[7]  _038_ \mprj_logic1[17]\ vssd vssd vccd vccd mprj_adr_o_user[7] sky130_fd_sc_hd__einvp_8
X\mprj_adr_buf[8]  _039_ \mprj_logic1[18]\ vssd vssd vccd vccd mprj_adr_o_user[8] sky130_fd_sc_hd__einvp_8
X\mprj_adr_buf[9]  _040_ \mprj_logic1[19]\ vssd vssd vccd vccd mprj_adr_o_user[9] sky130_fd_sc_hd__einvp_8
Xmprj_clk2_buf _001_ \mprj_logic1[2]\ vssd vssd vccd vccd user_clock2 sky130_fd_sc_hd__einvp_8
Xmprj_clk_buf _000_ \mprj_logic1[1]\ vssd vssd vccd vccd user_clock sky130_fd_sc_hd__einvp_8
Xmprj_cyc_buf _002_ \mprj_logic1[3]\ vssd vssd vccd vccd mprj_cyc_o_user sky130_fd_sc_hd__einvp_8
X\mprj_dat_buf[0]  _041_ \mprj_logic1[42]\ vssd vssd vccd vccd mprj_dat_o_user[0] sky130_fd_sc_hd__einvp_8
X\mprj_dat_buf[10]  _042_ \mprj_logic1[52]\ vssd vssd vccd vccd mprj_dat_o_user[10] sky130_fd_sc_hd__einvp_8
X\mprj_dat_buf[11]  _043_ \mprj_logic1[53]\ vssd vssd vccd vccd mprj_dat_o_user[11] sky130_fd_sc_hd__einvp_8
X\mprj_dat_buf[12]  _044_ \mprj_logic1[54]\ vssd vssd vccd vccd mprj_dat_o_user[12] sky130_fd_sc_hd__einvp_8
X\mprj_dat_buf[13]  _045_ \mprj_logic1[55]\ vssd vssd vccd vccd mprj_dat_o_user[13] sky130_fd_sc_hd__einvp_8
X\mprj_dat_buf[14]  _046_ \mprj_logic1[56]\ vssd vssd vccd vccd mprj_dat_o_user[14] sky130_fd_sc_hd__einvp_8
X\mprj_dat_buf[15]  _047_ \mprj_logic1[57]\ vssd vssd vccd vccd mprj_dat_o_user[15] sky130_fd_sc_hd__einvp_8
X\mprj_dat_buf[16]  _048_ \mprj_logic1[58]\ vssd vssd vccd vccd mprj_dat_o_user[16] sky130_fd_sc_hd__einvp_8
X\mprj_dat_buf[17]  _049_ \mprj_logic1[59]\ vssd vssd vccd vccd mprj_dat_o_user[17] sky130_fd_sc_hd__einvp_8
X\mprj_dat_buf[18]  _050_ \mprj_logic1[60]\ vssd vssd vccd vccd mprj_dat_o_user[18] sky130_fd_sc_hd__einvp_8
X\mprj_dat_buf[19]  _051_ \mprj_logic1[61]\ vssd vssd vccd vccd mprj_dat_o_user[19] sky130_fd_sc_hd__einvp_8
X\mprj_dat_buf[1]  _052_ \mprj_logic1[43]\ vssd vssd vccd vccd mprj_dat_o_user[1] sky130_fd_sc_hd__einvp_8
X\mprj_dat_buf[20]  _053_ \mprj_logic1[62]\ vssd vssd vccd vccd mprj_dat_o_user[20] sky130_fd_sc_hd__einvp_8
X\mprj_dat_buf[21]  _054_ \mprj_logic1[63]\ vssd vssd vccd vccd mprj_dat_o_user[21] sky130_fd_sc_hd__einvp_8
X\mprj_dat_buf[22]  _055_ \mprj_logic1[64]\ vssd vssd vccd vccd mprj_dat_o_user[22] sky130_fd_sc_hd__einvp_8
X\mprj_dat_buf[23]  _056_ \mprj_logic1[65]\ vssd vssd vccd vccd mprj_dat_o_user[23] sky130_fd_sc_hd__einvp_8
X\mprj_dat_buf[24]  _057_ \mprj_logic1[66]\ vssd vssd vccd vccd mprj_dat_o_user[24] sky130_fd_sc_hd__einvp_8
X\mprj_dat_buf[25]  _058_ \mprj_logic1[67]\ vssd vssd vccd vccd mprj_dat_o_user[25] sky130_fd_sc_hd__einvp_8
X\mprj_dat_buf[26]  _059_ \mprj_logic1[68]\ vssd vssd vccd vccd mprj_dat_o_user[26] sky130_fd_sc_hd__einvp_8
X\mprj_dat_buf[27]  _060_ \mprj_logic1[69]\ vssd vssd vccd vccd mprj_dat_o_user[27] sky130_fd_sc_hd__einvp_8
X\mprj_dat_buf[28]  _061_ \mprj_logic1[70]\ vssd vssd vccd vccd mprj_dat_o_user[28] sky130_fd_sc_hd__einvp_8
X\mprj_dat_buf[29]  _062_ \mprj_logic1[71]\ vssd vssd vccd vccd mprj_dat_o_user[29] sky130_fd_sc_hd__einvp_8
X\mprj_dat_buf[2]  _063_ \mprj_logic1[44]\ vssd vssd vccd vccd mprj_dat_o_user[2] sky130_fd_sc_hd__einvp_8
X\mprj_dat_buf[30]  _064_ \mprj_logic1[72]\ vssd vssd vccd vccd mprj_dat_o_user[30] sky130_fd_sc_hd__einvp_8
X\mprj_dat_buf[31]  _065_ \mprj_logic1[73]\ vssd vssd vccd vccd mprj_dat_o_user[31] sky130_fd_sc_hd__einvp_8
X\mprj_dat_buf[3]  _066_ \mprj_logic1[45]\ vssd vssd vccd vccd mprj_dat_o_user[3] sky130_fd_sc_hd__einvp_8
X\mprj_dat_buf[4]  _067_ \mprj_logic1[46]\ vssd vssd vccd vccd mprj_dat_o_user[4] sky130_fd_sc_hd__einvp_8
X\mprj_dat_buf[5]  _068_ \mprj_logic1[47]\ vssd vssd vccd vccd mprj_dat_o_user[5] sky130_fd_sc_hd__einvp_8
X\mprj_dat_buf[6]  _069_ \mprj_logic1[48]\ vssd vssd vccd vccd mprj_dat_o_user[6] sky130_fd_sc_hd__einvp_8
X\mprj_dat_buf[7]  _070_ \mprj_logic1[49]\ vssd vssd vccd vccd mprj_dat_o_user[7] sky130_fd_sc_hd__einvp_8
X\mprj_dat_buf[8]  _071_ \mprj_logic1[50]\ vssd vssd vccd vccd mprj_dat_o_user[8] sky130_fd_sc_hd__einvp_8
X\mprj_dat_buf[9]  _072_ \mprj_logic1[51]\ vssd vssd vccd vccd mprj_dat_o_user[9] sky130_fd_sc_hd__einvp_8
Xmprj_logic_high_inst vccd1 vssd1 {\mprj_logic1[462] ,\mprj_logic1[461] ,\mprj_logic1[460] ,\mprj_logic1[459] ,\mprj_logic1[458] ,\mprj_logic1[457] ,\mprj_logic1[456] ,\mprj_logic1[455] ,\mprj_logic1[454] ,\mprj_logic1[453] ,\mprj_logic1[452] ,\mprj_logic1[451] ,\mprj_logic1[450] ,\mprj_logic1[449] ,\mprj_logic1[448] ,\mprj_logic1[447] ,\mprj_logic1[446] ,\mprj_logic1[445] ,\mprj_logic1[444] ,\mprj_logic1[443] ,\mprj_logic1[442] ,\mprj_logic1[441] ,\mprj_logic1[440] ,\mprj_logic1[439] ,\mprj_logic1[438] ,\mprj_logic1[437] ,\mprj_logic1[436] ,\mprj_logic1[435] ,\mprj_logic1[434] ,\mprj_logic1[433] ,\mprj_logic1[432] ,\mprj_logic1[431] ,\mprj_logic1[430] ,\mprj_logic1[429] ,\mprj_logic1[428] ,\mprj_logic1[427] ,\mprj_logic1[426] ,\mprj_logic1[425] ,\mprj_logic1[424] ,\mprj_logic1[423] ,\mprj_logic1[422] ,\mprj_logic1[421] ,\mprj_logic1[420] ,\mprj_logic1[419] ,\mprj_logic1[418] ,\mprj_logic1[417] ,\mprj_logic1[416] ,\mprj_logic1[415] ,\mprj_logic1[414] ,\mprj_logic1[413] ,\mprj_logic1[412] ,\mprj_logic1[411] ,\mprj_logic1[410] ,\mprj_logic1[409] ,\mprj_logic1[408] ,\mprj_logic1[407] ,\mprj_logic1[406] ,\mprj_logic1[405] ,\mprj_logic1[404] ,\mprj_logic1[403] ,\mprj_logic1[402] ,\mprj_logic1[401] ,\mprj_logic1[400] ,\mprj_logic1[399] ,\mprj_logic1[398] ,\mprj_logic1[397] ,\mprj_logic1[396] ,\mprj_logic1[395] ,\mprj_logic1[394] ,\mprj_logic1[393] ,\mprj_logic1[392] ,\mprj_logic1[391] ,\mprj_logic1[390] ,\mprj_logic1[389] ,\mprj_logic1[388] ,\mprj_logic1[387] ,\mprj_logic1[386] ,\mprj_logic1[385] ,\mprj_logic1[384] ,\mprj_logic1[383] ,\mprj_logic1[382] ,\mprj_logic1[381] ,\mprj_logic1[380] ,\mprj_logic1[379] ,\mprj_logic1[378] ,\mprj_logic1[377] ,\mprj_logic1[376] ,\mprj_logic1[375] ,\mprj_logic1[374] ,\mprj_logic1[373] ,\mprj_logic1[372] ,\mprj_logic1[371] ,\mprj_logic1[370] ,\mprj_logic1[369] ,\mprj_logic1[368] ,\mprj_logic1[367] ,\mprj_logic1[366] ,\mprj_logic1[365] ,\mprj_logic1[364] ,\mprj_logic1[363] ,\mprj_logic1[362] ,\mprj_logic1[361] ,\mprj_logic1[360] ,\mprj_logic1[359] ,\mprj_logic1[358] ,\mprj_logic1[357] ,\mprj_logic1[356] ,\mprj_logic1[355] ,\mprj_logic1[354] ,\mprj_logic1[353] ,\mprj_logic1[352] ,\mprj_logic1[351] ,\mprj_logic1[350] ,\mprj_logic1[349] ,\mprj_logic1[348] ,\mprj_logic1[347] ,\mprj_logic1[346] ,\mprj_logic1[345] ,\mprj_logic1[344] ,\mprj_logic1[343] ,\mprj_logic1[342] ,\mprj_logic1[341] ,\mprj_logic1[340] ,\mprj_logic1[339] ,\mprj_logic1[338] ,\mprj_logic1[337] ,\mprj_logic1[336] ,\mprj_logic1[335] ,\mprj_logic1[334] ,\mprj_logic1[333] ,\mprj_logic1[332] ,\mprj_logic1[331] ,\mprj_logic1[330] ,\mprj_logic1[329] ,\mprj_logic1[328] ,\mprj_logic1[327] ,\mprj_logic1[326] ,\mprj_logic1[325] ,\mprj_logic1[324] ,\mprj_logic1[323] ,\mprj_logic1[322] ,\mprj_logic1[321] ,\mprj_logic1[320] ,\mprj_logic1[319] ,\mprj_logic1[318] ,\mprj_logic1[317] ,\mprj_logic1[316] ,\mprj_logic1[315] ,\mprj_logic1[314] ,\mprj_logic1[313] ,\mprj_logic1[312] ,\mprj_logic1[311] ,\mprj_logic1[310] ,\mprj_logic1[309] ,\mprj_logic1[308] ,\mprj_logic1[307] ,\mprj_logic1[306] ,\mprj_logic1[305] ,\mprj_logic1[304] ,\mprj_logic1[303] ,\mprj_logic1[302] ,\mprj_logic1[301] ,\mprj_logic1[300] ,\mprj_logic1[299] ,\mprj_logic1[298] ,\mprj_logic1[297] ,\mprj_logic1[296] ,\mprj_logic1[295] ,\mprj_logic1[294] ,\mprj_logic1[293] ,\mprj_logic1[292] ,\mprj_logic1[291] ,\mprj_logic1[290] ,\mprj_logic1[289] ,\mprj_logic1[288] ,\mprj_logic1[287] ,\mprj_logic1[286] ,\mprj_logic1[285] ,\mprj_logic1[284] ,\mprj_logic1[283] ,\mprj_logic1[282] ,\mprj_logic1[281] ,\mprj_logic1[280] ,\mprj_logic1[279] ,\mprj_logic1[278] ,\mprj_logic1[277] ,\mprj_logic1[276] ,\mprj_logic1[275] ,\mprj_logic1[274] ,\mprj_logic1[273] ,\mprj_logic1[272] ,\mprj_logic1[271] ,\mprj_logic1[270] ,\mprj_logic1[269] ,\mprj_logic1[268] ,\mprj_logic1[267] ,\mprj_logic1[266] ,\mprj_logic1[265] ,\mprj_logic1[264] ,\mprj_logic1[263] ,\mprj_logic1[262] ,\mprj_logic1[261] ,\mprj_logic1[260] ,\mprj_logic1[259] ,\mprj_logic1[258] ,\mprj_logic1[257] ,\mprj_logic1[256] ,\mprj_logic1[255] ,\mprj_logic1[254] ,\mprj_logic1[253] ,\mprj_logic1[252] ,\mprj_logic1[251] ,\mprj_logic1[250] ,\mprj_logic1[249] ,\mprj_logic1[248] ,\mprj_logic1[247] ,\mprj_logic1[246] ,\mprj_logic1[245] ,\mprj_logic1[244] ,\mprj_logic1[243] ,\mprj_logic1[242] ,\mprj_logic1[241] ,\mprj_logic1[240] ,\mprj_logic1[239] ,\mprj_logic1[238] ,\mprj_logic1[237] ,\mprj_logic1[236] ,\mprj_logic1[235] ,\mprj_logic1[234] ,\mprj_logic1[233] ,\mprj_logic1[232] ,\mprj_logic1[231] ,\mprj_logic1[230] ,\mprj_logic1[229] ,\mprj_logic1[228] ,\mprj_logic1[227] ,\mprj_logic1[226] ,\mprj_logic1[225] ,\mprj_logic1[224] ,\mprj_logic1[223] ,\mprj_logic1[222] ,\mprj_logic1[221] ,\mprj_logic1[220] ,\mprj_logic1[219] ,\mprj_logic1[218] ,\mprj_logic1[217] ,\mprj_logic1[216] ,\mprj_logic1[215] ,\mprj_logic1[214] ,\mprj_logic1[213] ,\mprj_logic1[212] ,\mprj_logic1[211] ,\mprj_logic1[210] ,\mprj_logic1[209] ,\mprj_logic1[208] ,\mprj_logic1[207] ,\mprj_logic1[206] ,\mprj_logic1[205] ,\mprj_logic1[204] ,\mprj_logic1[203] ,\mprj_logic1[202] ,\mprj_logic1[201] ,\mprj_logic1[200] ,\mprj_logic1[199] ,\mprj_logic1[198] ,\mprj_logic1[197] ,\mprj_logic1[196] ,\mprj_logic1[195] ,\mprj_logic1[194] ,\mprj_logic1[193] ,\mprj_logic1[192] ,\mprj_logic1[191] ,\mprj_logic1[190] ,\mprj_logic1[189] ,\mprj_logic1[188] ,\mprj_logic1[187] ,\mprj_logic1[186] ,\mprj_logic1[185] ,\mprj_logic1[184] ,\mprj_logic1[183] ,\mprj_logic1[182] ,\mprj_logic1[181] ,\mprj_logic1[180] ,\mprj_logic1[179] ,\mprj_logic1[178] ,\mprj_logic1[177] ,\mprj_logic1[176] ,\mprj_logic1[175] ,\mprj_logic1[174] ,\mprj_logic1[173] ,\mprj_logic1[172] ,\mprj_logic1[171] ,\mprj_logic1[170] ,\mprj_logic1[169] ,\mprj_logic1[168] ,\mprj_logic1[167] ,\mprj_logic1[166] ,\mprj_logic1[165] ,\mprj_logic1[164] ,\mprj_logic1[163] ,\mprj_logic1[162] ,\mprj_logic1[161] ,\mprj_logic1[160] ,\mprj_logic1[159] ,\mprj_logic1[158] ,\mprj_logic1[157] ,\mprj_logic1[156] ,\mprj_logic1[155] ,\mprj_logic1[154] ,\mprj_logic1[153] ,\mprj_logic1[152] ,\mprj_logic1[151] ,\mprj_logic1[150] ,\mprj_logic1[149] ,\mprj_logic1[148] ,\mprj_logic1[147] ,\mprj_logic1[146] ,\mprj_logic1[145] ,\mprj_logic1[144] ,\mprj_logic1[143] ,\mprj_logic1[142] ,\mprj_logic1[141] ,\mprj_logic1[140] ,\mprj_logic1[139] ,\mprj_logic1[138] ,\mprj_logic1[137] ,\mprj_logic1[136] ,\mprj_logic1[135] ,\mprj_logic1[134] ,\mprj_logic1[133] ,\mprj_logic1[132] ,\mprj_logic1[131] ,\mprj_logic1[130] ,\mprj_logic1[129] ,\mprj_logic1[128] ,\mprj_logic1[127] ,\mprj_logic1[126] ,\mprj_logic1[125] ,\mprj_logic1[124] ,\mprj_logic1[123] ,\mprj_logic1[122] ,\mprj_logic1[121] ,\mprj_logic1[120] ,\mprj_logic1[119] ,\mprj_logic1[118] ,\mprj_logic1[117] ,\mprj_logic1[116] ,\mprj_logic1[115] ,\mprj_logic1[114] ,\mprj_logic1[113] ,\mprj_logic1[112] ,\mprj_logic1[111] ,\mprj_logic1[110] ,\mprj_logic1[109] ,\mprj_logic1[108] ,\mprj_logic1[107] ,\mprj_logic1[106] ,\mprj_logic1[105] ,\mprj_logic1[104] ,\mprj_logic1[103] ,\mprj_logic1[102] ,\mprj_logic1[101] ,\mprj_logic1[100] ,\mprj_logic1[99] ,\mprj_logic1[98] ,\mprj_logic1[97] ,\mprj_logic1[96] ,\mprj_logic1[95] ,\mprj_logic1[94] ,\mprj_logic1[93] ,\mprj_logic1[92] ,\mprj_logic1[91] ,\mprj_logic1[90] ,\mprj_logic1[89] ,\mprj_logic1[88] ,\mprj_logic1[87] ,\mprj_logic1[86] ,\mprj_logic1[85] ,\mprj_logic1[84] ,\mprj_logic1[83] ,\mprj_logic1[82] ,\mprj_logic1[81] ,\mprj_logic1[80] ,\mprj_logic1[79] ,\mprj_logic1[78] ,\mprj_logic1[77] ,\mprj_logic1[76] ,\mprj_logic1[75] ,\mprj_logic1[74] ,\mprj_logic1[73] ,\mprj_logic1[72] ,\mprj_logic1[71] ,\mprj_logic1[70] ,\mprj_logic1[69] ,\mprj_logic1[68] ,\mprj_logic1[67] ,\mprj_logic1[66] ,\mprj_logic1[65] ,\mprj_logic1[64] ,\mprj_logic1[63] ,\mprj_logic1[62] ,\mprj_logic1[61] ,\mprj_logic1[60] ,\mprj_logic1[59] ,\mprj_logic1[58] ,\mprj_logic1[57] ,\mprj_logic1[56] ,\mprj_logic1[55] ,\mprj_logic1[54] ,\mprj_logic1[53] ,\mprj_logic1[52] ,\mprj_logic1[51] ,\mprj_logic1[50] ,\mprj_logic1[49] ,\mprj_logic1[48] ,\mprj_logic1[47] ,\mprj_logic1[46] ,\mprj_logic1[45] ,\mprj_logic1[44] ,\mprj_logic1[43] ,\mprj_logic1[42] ,\mprj_logic1[41] ,\mprj_logic1[40] ,\mprj_logic1[39] ,\mprj_logic1[38] ,\mprj_logic1[37] ,\mprj_logic1[36] ,\mprj_logic1[35] ,\mprj_logic1[34] ,\mprj_logic1[33] ,\mprj_logic1[32] ,\mprj_logic1[31] ,\mprj_logic1[30] ,\mprj_logic1[29] ,\mprj_logic1[28] ,\mprj_logic1[27] ,\mprj_logic1[26] ,\mprj_logic1[25] ,\mprj_logic1[24] ,\mprj_logic1[23] ,\mprj_logic1[22] ,\mprj_logic1[21] ,\mprj_logic1[20] ,\mprj_logic1[19] ,\mprj_logic1[18] ,\mprj_logic1[17] ,\mprj_logic1[16] ,\mprj_logic1[15] ,\mprj_logic1[14] ,\mprj_logic1[13] ,\mprj_logic1[12] ,\mprj_logic1[11] ,\mprj_logic1[10] ,\mprj_logic1[9] ,\mprj_logic1[8] ,\mprj_logic1[7] ,\mprj_logic1[6] ,\mprj_logic1[5] ,\mprj_logic1[4] ,\mprj_logic1[3] ,\mprj_logic1[2] ,\mprj_logic1[1] ,\mprj_logic1[0] } mprj_logic_high
Xmprj_pwrgood \mprj_logic1[461]\ vssd vssd vccd vccd net788 sky130_fd_sc_hd__buf_6
Xmprj_rstn_buf net3 \mprj_logic1[0]\ vssd vssd vccd vccd user_reset sky130_fd_sc_hd__einvp_8
X\mprj_sel_buf[0]  _005_ \mprj_logic1[6]\ vssd vssd vccd vccd mprj_sel_o_user[0] sky130_fd_sc_hd__einvp_8
X\mprj_sel_buf[1]  _006_ \mprj_logic1[7]\ vssd vssd vccd vccd mprj_sel_o_user[1] sky130_fd_sc_hd__einvp_8
X\mprj_sel_buf[2]  _007_ \mprj_logic1[8]\ vssd vssd vccd vccd mprj_sel_o_user[2] sky130_fd_sc_hd__einvp_8
X\mprj_sel_buf[3]  _008_ \mprj_logic1[9]\ vssd vssd vccd vccd mprj_sel_o_user[3] sky130_fd_sc_hd__einvp_8
Xmprj_stb_buf _003_ \mprj_logic1[4]\ vssd vssd vccd vccd mprj_stb_o_user sky130_fd_sc_hd__einvp_8
Xmprj_vdd_pwrgood mprj_vdd_logic1 vssd vssd vccd vccd net789 sky130_fd_sc_hd__buf_6
Xmprj_we_buf _004_ \mprj_logic1[5]\ vssd vssd vccd vccd mprj_we_o_user sky130_fd_sc_hd__einvp_8
Xoutput627 net627 vssd vssd vccd vccd la_data_in_mprj[0] sky130_fd_sc_hd__buf_2
Xoutput628 net628 vssd vssd vccd vccd la_data_in_mprj[100] sky130_fd_sc_hd__buf_2
Xoutput629 net629 vssd vssd vccd vccd la_data_in_mprj[101] sky130_fd_sc_hd__buf_2
Xoutput630 net630 vssd vssd vccd vccd la_data_in_mprj[102] sky130_fd_sc_hd__buf_2
Xoutput631 net631 vssd vssd vccd vccd la_data_in_mprj[103] sky130_fd_sc_hd__buf_2
Xoutput632 net632 vssd vssd vccd vccd la_data_in_mprj[104] sky130_fd_sc_hd__buf_2
Xoutput633 net633 vssd vssd vccd vccd la_data_in_mprj[105] sky130_fd_sc_hd__buf_2
Xoutput634 net634 vssd vssd vccd vccd la_data_in_mprj[106] sky130_fd_sc_hd__buf_2
Xoutput635 net635 vssd vssd vccd vccd la_data_in_mprj[107] sky130_fd_sc_hd__buf_2
Xoutput636 net636 vssd vssd vccd vccd la_data_in_mprj[108] sky130_fd_sc_hd__buf_2
Xoutput637 net637 vssd vssd vccd vccd la_data_in_mprj[109] sky130_fd_sc_hd__buf_2
Xoutput638 net638 vssd vssd vccd vccd la_data_in_mprj[10] sky130_fd_sc_hd__buf_2
Xoutput639 net639 vssd vssd vccd vccd la_data_in_mprj[110] sky130_fd_sc_hd__buf_2
Xoutput640 net640 vssd vssd vccd vccd la_data_in_mprj[111] sky130_fd_sc_hd__buf_2
Xoutput641 net641 vssd vssd vccd vccd la_data_in_mprj[112] sky130_fd_sc_hd__buf_2
Xoutput642 net642 vssd vssd vccd vccd la_data_in_mprj[113] sky130_fd_sc_hd__buf_2
Xoutput643 net643 vssd vssd vccd vccd la_data_in_mprj[114] sky130_fd_sc_hd__buf_2
Xoutput644 net644 vssd vssd vccd vccd la_data_in_mprj[115] sky130_fd_sc_hd__buf_2
Xoutput645 net645 vssd vssd vccd vccd la_data_in_mprj[116] sky130_fd_sc_hd__buf_2
Xoutput646 net646 vssd vssd vccd vccd la_data_in_mprj[117] sky130_fd_sc_hd__buf_2
Xoutput647 net647 vssd vssd vccd vccd la_data_in_mprj[118] sky130_fd_sc_hd__buf_2
Xoutput648 net648 vssd vssd vccd vccd la_data_in_mprj[119] sky130_fd_sc_hd__buf_2
Xoutput649 net649 vssd vssd vccd vccd la_data_in_mprj[11] sky130_fd_sc_hd__buf_2
Xoutput650 net650 vssd vssd vccd vccd la_data_in_mprj[120] sky130_fd_sc_hd__buf_2
Xoutput651 net651 vssd vssd vccd vccd la_data_in_mprj[121] sky130_fd_sc_hd__buf_2
Xoutput652 net652 vssd vssd vccd vccd la_data_in_mprj[122] sky130_fd_sc_hd__buf_2
Xoutput653 net653 vssd vssd vccd vccd la_data_in_mprj[123] sky130_fd_sc_hd__buf_2
Xoutput654 net654 vssd vssd vccd vccd la_data_in_mprj[124] sky130_fd_sc_hd__buf_2
Xoutput655 net655 vssd vssd vccd vccd la_data_in_mprj[125] sky130_fd_sc_hd__buf_2
Xoutput656 net656 vssd vssd vccd vccd la_data_in_mprj[126] sky130_fd_sc_hd__buf_2
Xoutput657 net657 vssd vssd vccd vccd la_data_in_mprj[127] sky130_fd_sc_hd__buf_2
Xoutput658 net658 vssd vssd vccd vccd la_data_in_mprj[12] sky130_fd_sc_hd__buf_2
Xoutput659 net659 vssd vssd vccd vccd la_data_in_mprj[13] sky130_fd_sc_hd__buf_2
Xoutput660 net660 vssd vssd vccd vccd la_data_in_mprj[14] sky130_fd_sc_hd__buf_2
Xoutput661 net661 vssd vssd vccd vccd la_data_in_mprj[15] sky130_fd_sc_hd__buf_2
Xoutput662 net662 vssd vssd vccd vccd la_data_in_mprj[16] sky130_fd_sc_hd__buf_2
Xoutput663 net663 vssd vssd vccd vccd la_data_in_mprj[17] sky130_fd_sc_hd__buf_2
Xoutput664 net664 vssd vssd vccd vccd la_data_in_mprj[18] sky130_fd_sc_hd__buf_2
Xoutput665 net665 vssd vssd vccd vccd la_data_in_mprj[19] sky130_fd_sc_hd__buf_2
Xoutput666 net666 vssd vssd vccd vccd la_data_in_mprj[1] sky130_fd_sc_hd__buf_2
Xoutput667 net667 vssd vssd vccd vccd la_data_in_mprj[20] sky130_fd_sc_hd__buf_2
Xoutput668 net668 vssd vssd vccd vccd la_data_in_mprj[21] sky130_fd_sc_hd__buf_2
Xoutput669 net669 vssd vssd vccd vccd la_data_in_mprj[22] sky130_fd_sc_hd__buf_2
Xoutput670 net670 vssd vssd vccd vccd la_data_in_mprj[23] sky130_fd_sc_hd__buf_2
Xoutput671 net671 vssd vssd vccd vccd la_data_in_mprj[24] sky130_fd_sc_hd__buf_2
Xoutput672 net672 vssd vssd vccd vccd la_data_in_mprj[25] sky130_fd_sc_hd__buf_2
Xoutput673 net673 vssd vssd vccd vccd la_data_in_mprj[26] sky130_fd_sc_hd__buf_2
Xoutput674 net674 vssd vssd vccd vccd la_data_in_mprj[27] sky130_fd_sc_hd__buf_2
Xoutput675 net675 vssd vssd vccd vccd la_data_in_mprj[28] sky130_fd_sc_hd__buf_2
Xoutput676 net676 vssd vssd vccd vccd la_data_in_mprj[29] sky130_fd_sc_hd__buf_2
Xoutput677 net677 vssd vssd vccd vccd la_data_in_mprj[2] sky130_fd_sc_hd__buf_2
Xoutput678 net678 vssd vssd vccd vccd la_data_in_mprj[30] sky130_fd_sc_hd__buf_2
Xoutput679 net679 vssd vssd vccd vccd la_data_in_mprj[31] sky130_fd_sc_hd__buf_2
Xoutput680 net680 vssd vssd vccd vccd la_data_in_mprj[32] sky130_fd_sc_hd__buf_2
Xoutput681 net681 vssd vssd vccd vccd la_data_in_mprj[33] sky130_fd_sc_hd__buf_2
Xoutput682 net682 vssd vssd vccd vccd la_data_in_mprj[34] sky130_fd_sc_hd__buf_2
Xoutput683 net683 vssd vssd vccd vccd la_data_in_mprj[35] sky130_fd_sc_hd__buf_2
Xoutput684 net684 vssd vssd vccd vccd la_data_in_mprj[36] sky130_fd_sc_hd__buf_2
Xoutput685 net685 vssd vssd vccd vccd la_data_in_mprj[37] sky130_fd_sc_hd__buf_2
Xoutput686 net686 vssd vssd vccd vccd la_data_in_mprj[38] sky130_fd_sc_hd__buf_2
Xoutput687 net687 vssd vssd vccd vccd la_data_in_mprj[39] sky130_fd_sc_hd__buf_2
Xoutput688 net688 vssd vssd vccd vccd la_data_in_mprj[3] sky130_fd_sc_hd__buf_2
Xoutput689 net689 vssd vssd vccd vccd la_data_in_mprj[40] sky130_fd_sc_hd__buf_2
Xoutput690 net690 vssd vssd vccd vccd la_data_in_mprj[41] sky130_fd_sc_hd__buf_2
Xoutput691 net691 vssd vssd vccd vccd la_data_in_mprj[42] sky130_fd_sc_hd__buf_2
Xoutput692 net692 vssd vssd vccd vccd la_data_in_mprj[43] sky130_fd_sc_hd__buf_2
Xoutput693 net693 vssd vssd vccd vccd la_data_in_mprj[44] sky130_fd_sc_hd__buf_2
Xoutput694 net694 vssd vssd vccd vccd la_data_in_mprj[45] sky130_fd_sc_hd__buf_2
Xoutput695 net695 vssd vssd vccd vccd la_data_in_mprj[46] sky130_fd_sc_hd__buf_2
Xoutput696 net696 vssd vssd vccd vccd la_data_in_mprj[47] sky130_fd_sc_hd__buf_2
Xoutput697 net697 vssd vssd vccd vccd la_data_in_mprj[48] sky130_fd_sc_hd__buf_2
Xoutput698 net698 vssd vssd vccd vccd la_data_in_mprj[49] sky130_fd_sc_hd__buf_2
Xoutput699 net699 vssd vssd vccd vccd la_data_in_mprj[4] sky130_fd_sc_hd__buf_2
Xoutput700 net700 vssd vssd vccd vccd la_data_in_mprj[50] sky130_fd_sc_hd__buf_2
Xoutput701 net701 vssd vssd vccd vccd la_data_in_mprj[51] sky130_fd_sc_hd__buf_2
Xoutput702 net702 vssd vssd vccd vccd la_data_in_mprj[52] sky130_fd_sc_hd__buf_2
Xoutput703 net703 vssd vssd vccd vccd la_data_in_mprj[53] sky130_fd_sc_hd__buf_2
Xoutput704 net704 vssd vssd vccd vccd la_data_in_mprj[54] sky130_fd_sc_hd__buf_2
Xoutput705 net705 vssd vssd vccd vccd la_data_in_mprj[55] sky130_fd_sc_hd__buf_2
Xoutput706 net706 vssd vssd vccd vccd la_data_in_mprj[56] sky130_fd_sc_hd__buf_2
Xoutput707 net707 vssd vssd vccd vccd la_data_in_mprj[57] sky130_fd_sc_hd__buf_2
Xoutput708 net708 vssd vssd vccd vccd la_data_in_mprj[58] sky130_fd_sc_hd__buf_2
Xoutput709 net709 vssd vssd vccd vccd la_data_in_mprj[59] sky130_fd_sc_hd__buf_2
Xoutput710 net710 vssd vssd vccd vccd la_data_in_mprj[5] sky130_fd_sc_hd__buf_2
Xoutput711 net711 vssd vssd vccd vccd la_data_in_mprj[60] sky130_fd_sc_hd__buf_2
Xoutput712 net712 vssd vssd vccd vccd la_data_in_mprj[61] sky130_fd_sc_hd__buf_2
Xoutput713 net713 vssd vssd vccd vccd la_data_in_mprj[62] sky130_fd_sc_hd__buf_2
Xoutput714 net714 vssd vssd vccd vccd la_data_in_mprj[63] sky130_fd_sc_hd__buf_2
Xoutput715 net715 vssd vssd vccd vccd la_data_in_mprj[64] sky130_fd_sc_hd__buf_2
Xoutput716 net716 vssd vssd vccd vccd la_data_in_mprj[65] sky130_fd_sc_hd__buf_2
Xoutput717 net717 vssd vssd vccd vccd la_data_in_mprj[66] sky130_fd_sc_hd__buf_2
Xoutput718 net718 vssd vssd vccd vccd la_data_in_mprj[67] sky130_fd_sc_hd__buf_2
Xoutput719 net719 vssd vssd vccd vccd la_data_in_mprj[68] sky130_fd_sc_hd__buf_2
Xoutput720 net720 vssd vssd vccd vccd la_data_in_mprj[69] sky130_fd_sc_hd__buf_2
Xoutput721 net721 vssd vssd vccd vccd la_data_in_mprj[6] sky130_fd_sc_hd__buf_2
Xoutput722 net722 vssd vssd vccd vccd la_data_in_mprj[70] sky130_fd_sc_hd__buf_2
Xoutput723 net723 vssd vssd vccd vccd la_data_in_mprj[71] sky130_fd_sc_hd__buf_2
Xoutput724 net724 vssd vssd vccd vccd la_data_in_mprj[72] sky130_fd_sc_hd__buf_2
Xoutput725 net725 vssd vssd vccd vccd la_data_in_mprj[73] sky130_fd_sc_hd__buf_2
Xoutput726 net726 vssd vssd vccd vccd la_data_in_mprj[74] sky130_fd_sc_hd__buf_2
Xoutput727 net727 vssd vssd vccd vccd la_data_in_mprj[75] sky130_fd_sc_hd__buf_2
Xoutput728 net728 vssd vssd vccd vccd la_data_in_mprj[76] sky130_fd_sc_hd__buf_2
Xoutput729 net729 vssd vssd vccd vccd la_data_in_mprj[77] sky130_fd_sc_hd__buf_2
Xoutput730 net730 vssd vssd vccd vccd la_data_in_mprj[78] sky130_fd_sc_hd__buf_2
Xoutput731 net731 vssd vssd vccd vccd la_data_in_mprj[79] sky130_fd_sc_hd__buf_2
Xoutput732 net732 vssd vssd vccd vccd la_data_in_mprj[7] sky130_fd_sc_hd__buf_2
Xoutput733 net733 vssd vssd vccd vccd la_data_in_mprj[80] sky130_fd_sc_hd__buf_2
Xoutput734 net734 vssd vssd vccd vccd la_data_in_mprj[81] sky130_fd_sc_hd__buf_2
Xoutput735 net735 vssd vssd vccd vccd la_data_in_mprj[82] sky130_fd_sc_hd__buf_2
Xoutput736 net736 vssd vssd vccd vccd la_data_in_mprj[83] sky130_fd_sc_hd__buf_2
Xoutput737 net737 vssd vssd vccd vccd la_data_in_mprj[84] sky130_fd_sc_hd__buf_2
Xoutput738 net738 vssd vssd vccd vccd la_data_in_mprj[85] sky130_fd_sc_hd__buf_2
Xoutput739 net739 vssd vssd vccd vccd la_data_in_mprj[86] sky130_fd_sc_hd__buf_2
Xoutput740 net740 vssd vssd vccd vccd la_data_in_mprj[87] sky130_fd_sc_hd__buf_2
Xoutput741 net741 vssd vssd vccd vccd la_data_in_mprj[88] sky130_fd_sc_hd__buf_2
Xoutput742 net742 vssd vssd vccd vccd la_data_in_mprj[89] sky130_fd_sc_hd__buf_2
Xoutput743 net743 vssd vssd vccd vccd la_data_in_mprj[8] sky130_fd_sc_hd__buf_2
Xoutput744 net744 vssd vssd vccd vccd la_data_in_mprj[90] sky130_fd_sc_hd__buf_2
Xoutput745 net745 vssd vssd vccd vccd la_data_in_mprj[91] sky130_fd_sc_hd__buf_2
Xoutput746 net746 vssd vssd vccd vccd la_data_in_mprj[92] sky130_fd_sc_hd__buf_2
Xoutput747 net747 vssd vssd vccd vccd la_data_in_mprj[93] sky130_fd_sc_hd__buf_2
Xoutput748 net748 vssd vssd vccd vccd la_data_in_mprj[94] sky130_fd_sc_hd__buf_2
Xoutput749 net749 vssd vssd vccd vccd la_data_in_mprj[95] sky130_fd_sc_hd__buf_2
Xoutput750 net750 vssd vssd vccd vccd la_data_in_mprj[96] sky130_fd_sc_hd__buf_2
Xoutput751 net751 vssd vssd vccd vccd la_data_in_mprj[97] sky130_fd_sc_hd__buf_2
Xoutput752 net752 vssd vssd vccd vccd la_data_in_mprj[98] sky130_fd_sc_hd__buf_2
Xoutput753 net753 vssd vssd vccd vccd la_data_in_mprj[99] sky130_fd_sc_hd__buf_2
Xoutput754 net754 vssd vssd vccd vccd la_data_in_mprj[9] sky130_fd_sc_hd__buf_2
Xoutput755 net755 vssd vssd vccd vccd mprj_ack_i_core sky130_fd_sc_hd__buf_2
Xoutput756 net756 vssd vssd vccd vccd mprj_dat_i_core[0] sky130_fd_sc_hd__buf_2
Xoutput757 net757 vssd vssd vccd vccd mprj_dat_i_core[10] sky130_fd_sc_hd__buf_2
Xoutput758 net758 vssd vssd vccd vccd mprj_dat_i_core[11] sky130_fd_sc_hd__buf_2
Xoutput759 net759 vssd vssd vccd vccd mprj_dat_i_core[12] sky130_fd_sc_hd__buf_2
Xoutput760 net760 vssd vssd vccd vccd mprj_dat_i_core[13] sky130_fd_sc_hd__buf_2
Xoutput761 net761 vssd vssd vccd vccd mprj_dat_i_core[14] sky130_fd_sc_hd__buf_2
Xoutput762 net762 vssd vssd vccd vccd mprj_dat_i_core[15] sky130_fd_sc_hd__buf_2
Xoutput763 net763 vssd vssd vccd vccd mprj_dat_i_core[16] sky130_fd_sc_hd__buf_2
Xoutput764 net764 vssd vssd vccd vccd mprj_dat_i_core[17] sky130_fd_sc_hd__buf_2
Xoutput765 net765 vssd vssd vccd vccd mprj_dat_i_core[18] sky130_fd_sc_hd__buf_2
Xoutput766 net766 vssd vssd vccd vccd mprj_dat_i_core[19] sky130_fd_sc_hd__buf_2
Xoutput767 net767 vssd vssd vccd vccd mprj_dat_i_core[1] sky130_fd_sc_hd__buf_2
Xoutput768 net768 vssd vssd vccd vccd mprj_dat_i_core[20] sky130_fd_sc_hd__buf_2
Xoutput769 net769 vssd vssd vccd vccd mprj_dat_i_core[21] sky130_fd_sc_hd__buf_2
Xoutput770 net770 vssd vssd vccd vccd mprj_dat_i_core[22] sky130_fd_sc_hd__buf_2
Xoutput771 net771 vssd vssd vccd vccd mprj_dat_i_core[23] sky130_fd_sc_hd__buf_2
Xoutput772 net772 vssd vssd vccd vccd mprj_dat_i_core[24] sky130_fd_sc_hd__buf_2
Xoutput773 net773 vssd vssd vccd vccd mprj_dat_i_core[25] sky130_fd_sc_hd__buf_2
Xoutput774 net774 vssd vssd vccd vccd mprj_dat_i_core[26] sky130_fd_sc_hd__buf_2
Xoutput775 net775 vssd vssd vccd vccd mprj_dat_i_core[27] sky130_fd_sc_hd__buf_2
Xoutput776 net776 vssd vssd vccd vccd mprj_dat_i_core[28] sky130_fd_sc_hd__buf_2
Xoutput777 net777 vssd vssd vccd vccd mprj_dat_i_core[29] sky130_fd_sc_hd__buf_2
Xoutput778 net778 vssd vssd vccd vccd mprj_dat_i_core[2] sky130_fd_sc_hd__buf_2
Xoutput779 net779 vssd vssd vccd vccd mprj_dat_i_core[30] sky130_fd_sc_hd__buf_2
Xoutput780 net780 vssd vssd vccd vccd mprj_dat_i_core[31] sky130_fd_sc_hd__buf_2
Xoutput781 net781 vssd vssd vccd vccd mprj_dat_i_core[3] sky130_fd_sc_hd__buf_2
Xoutput782 net782 vssd vssd vccd vccd mprj_dat_i_core[4] sky130_fd_sc_hd__buf_2
Xoutput783 net783 vssd vssd vccd vccd mprj_dat_i_core[5] sky130_fd_sc_hd__buf_2
Xoutput784 net784 vssd vssd vccd vccd mprj_dat_i_core[6] sky130_fd_sc_hd__buf_2
Xoutput785 net785 vssd vssd vccd vccd mprj_dat_i_core[7] sky130_fd_sc_hd__buf_2
Xoutput786 net786 vssd vssd vccd vccd mprj_dat_i_core[8] sky130_fd_sc_hd__buf_2
Xoutput787 net787 vssd vssd vccd vccd mprj_dat_i_core[9] sky130_fd_sc_hd__buf_2
Xoutput788 net788 vssd vssd vccd vccd user1_vcc_powergood sky130_fd_sc_hd__buf_2
Xoutput789 net789 vssd vssd vccd vccd user1_vdd_powergood sky130_fd_sc_hd__buf_2
Xoutput790 net790 vssd vssd vccd vccd user2_vcc_powergood sky130_fd_sc_hd__buf_2
Xoutput791 net791 vssd vssd vccd vccd user2_vdd_powergood sky130_fd_sc_hd__buf_2
Xoutput792 net792 vssd vssd vccd vccd user_irq[0] sky130_fd_sc_hd__buf_2
Xoutput793 net793 vssd vssd vccd vccd user_irq[1] sky130_fd_sc_hd__buf_2
Xoutput794 net794 vssd vssd vccd vccd user_irq[2] sky130_fd_sc_hd__buf_2
Xpowergood_check mprj2_vdd_logic1 mprj_vdd_logic1 vccd vssd vdda1 vssa1 vdda2 vssa2 mgmt_protect_hv
X\user_irq_buffers[0]  \user_irq_bar[0]\ vssd vssd vccd vccd net792 sky130_fd_sc_hd__clkinv_4
X\user_irq_buffers[1]  \user_irq_bar[1]\ vssd vssd vccd vccd net793 sky130_fd_sc_hd__clkinv_4
X\user_irq_buffers[2]  \user_irq_bar[2]\ vssd vssd vccd vccd net794 sky130_fd_sc_hd__clkinv_4
X\user_irq_ena_buf[0]  net624 \mprj_logic1[458]\ vssd vssd vccd vccd \user_irq_enable[0]\ sky130_fd_sc_hd__and2_1
X\user_irq_ena_buf[1]  net625 \mprj_logic1[459]\ vssd vssd vccd vccd \user_irq_enable[1]\ sky130_fd_sc_hd__and2_1
X\user_irq_ena_buf[2]  net626 \mprj_logic1[460]\ vssd vssd vccd vccd \user_irq_enable[2]\ sky130_fd_sc_hd__and2_1
X\user_irq_gates[0]  net621 \user_irq_enable[0]\ vssd vssd vccd vccd \user_irq_bar[0]\ sky130_fd_sc_hd__nand2_1
X\user_irq_gates[1]  net622 \user_irq_enable[1]\ vssd vssd vccd vccd \user_irq_bar[1]\ sky130_fd_sc_hd__nand2_1
X\user_irq_gates[2]  net623 \user_irq_enable[2]\ vssd vssd vccd vccd \user_irq_bar[2]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_buffers[0]  \la_data_in_mprj_bar[0]\ vssd vssd vccd vccd net627 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[100]  \la_data_in_mprj_bar[100]\ vssd vssd vccd vccd net628 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[101]  \la_data_in_mprj_bar[101]\ vssd vssd vccd vccd net629 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[102]  \la_data_in_mprj_bar[102]\ vssd vssd vccd vccd net630 sky130_fd_sc_hd__inv_2
X\user_to_mprj_in_buffers[103]  \la_data_in_mprj_bar[103]\ vssd vssd vccd vccd net631 sky130_fd_sc_hd__inv_2
X\user_to_mprj_in_buffers[104]  \la_data_in_mprj_bar[104]\ vssd vssd vccd vccd net632 sky130_fd_sc_hd__inv_2
X\user_to_mprj_in_buffers[105]  \la_data_in_mprj_bar[105]\ vssd vssd vccd vccd net633 sky130_fd_sc_hd__inv_2
X\user_to_mprj_in_buffers[106]  \la_data_in_mprj_bar[106]\ vssd vssd vccd vccd net634 sky130_fd_sc_hd__inv_2
X\user_to_mprj_in_buffers[107]  \la_data_in_mprj_bar[107]\ vssd vssd vccd vccd net635 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[108]  \la_data_in_mprj_bar[108]\ vssd vssd vccd vccd net636 sky130_fd_sc_hd__inv_2
X\user_to_mprj_in_buffers[109]  \la_data_in_mprj_bar[109]\ vssd vssd vccd vccd net637 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[10]  \la_data_in_mprj_bar[10]\ vssd vssd vccd vccd net638 sky130_fd_sc_hd__inv_6
X\user_to_mprj_in_buffers[110]  \la_data_in_mprj_bar[110]\ vssd vssd vccd vccd net639 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[111]  \la_data_in_mprj_bar[111]\ vssd vssd vccd vccd net640 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[112]  \la_data_in_mprj_bar[112]\ vssd vssd vccd vccd net641 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[113]  \la_data_in_mprj_bar[113]\ vssd vssd vccd vccd net642 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[114]  \la_data_in_mprj_bar[114]\ vssd vssd vccd vccd net643 sky130_fd_sc_hd__inv_2
X\user_to_mprj_in_buffers[115]  \la_data_in_mprj_bar[115]\ vssd vssd vccd vccd net644 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[116]  \la_data_in_mprj_bar[116]\ vssd vssd vccd vccd net645 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[117]  \la_data_in_mprj_bar[117]\ vssd vssd vccd vccd net646 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[118]  \la_data_in_mprj_bar[118]\ vssd vssd vccd vccd net647 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[119]  \la_data_in_mprj_bar[119]\ vssd vssd vccd vccd net648 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[11]  \la_data_in_mprj_bar[11]\ vssd vssd vccd vccd net649 sky130_fd_sc_hd__inv_6
X\user_to_mprj_in_buffers[120]  \la_data_in_mprj_bar[120]\ vssd vssd vccd vccd net650 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[121]  \la_data_in_mprj_bar[121]\ vssd vssd vccd vccd net651 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[122]  \la_data_in_mprj_bar[122]\ vssd vssd vccd vccd net652 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[123]  \la_data_in_mprj_bar[123]\ vssd vssd vccd vccd net653 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[124]  \la_data_in_mprj_bar[124]\ vssd vssd vccd vccd net654 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[125]  \la_data_in_mprj_bar[125]\ vssd vssd vccd vccd net655 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[126]  \la_data_in_mprj_bar[126]\ vssd vssd vccd vccd net656 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[127]  \la_data_in_mprj_bar[127]\ vssd vssd vccd vccd net657 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[12]  \la_data_in_mprj_bar[12]\ vssd vssd vccd vccd net658 sky130_fd_sc_hd__clkinv_8
X\user_to_mprj_in_buffers[13]  \la_data_in_mprj_bar[13]\ vssd vssd vccd vccd net659 sky130_fd_sc_hd__inv_2
X\user_to_mprj_in_buffers[14]  \la_data_in_mprj_bar[14]\ vssd vssd vccd vccd net660 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[15]  \la_data_in_mprj_bar[15]\ vssd vssd vccd vccd net661 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[16]  \la_data_in_mprj_bar[16]\ vssd vssd vccd vccd net662 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[17]  \la_data_in_mprj_bar[17]\ vssd vssd vccd vccd net663 sky130_fd_sc_hd__inv_2
X\user_to_mprj_in_buffers[18]  \la_data_in_mprj_bar[18]\ vssd vssd vccd vccd net664 sky130_fd_sc_hd__inv_2
X\user_to_mprj_in_buffers[19]  \la_data_in_mprj_bar[19]\ vssd vssd vccd vccd net665 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[1]  \la_data_in_mprj_bar[1]\ vssd vssd vccd vccd net666 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[20]  \la_data_in_mprj_bar[20]\ vssd vssd vccd vccd net667 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[21]  \la_data_in_mprj_bar[21]\ vssd vssd vccd vccd net668 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[22]  \la_data_in_mprj_bar[22]\ vssd vssd vccd vccd net669 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[23]  \la_data_in_mprj_bar[23]\ vssd vssd vccd vccd net670 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[24]  \la_data_in_mprj_bar[24]\ vssd vssd vccd vccd net671 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[25]  \la_data_in_mprj_bar[25]\ vssd vssd vccd vccd net672 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[26]  \la_data_in_mprj_bar[26]\ vssd vssd vccd vccd net673 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[27]  \la_data_in_mprj_bar[27]\ vssd vssd vccd vccd net674 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[28]  \la_data_in_mprj_bar[28]\ vssd vssd vccd vccd net675 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[29]  \la_data_in_mprj_bar[29]\ vssd vssd vccd vccd net676 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[2]  \la_data_in_mprj_bar[2]\ vssd vssd vccd vccd net677 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[30]  \la_data_in_mprj_bar[30]\ vssd vssd vccd vccd net678 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[31]  \la_data_in_mprj_bar[31]\ vssd vssd vccd vccd net679 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[32]  \la_data_in_mprj_bar[32]\ vssd vssd vccd vccd net680 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[33]  \la_data_in_mprj_bar[33]\ vssd vssd vccd vccd net681 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[34]  \la_data_in_mprj_bar[34]\ vssd vssd vccd vccd net682 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[35]  \la_data_in_mprj_bar[35]\ vssd vssd vccd vccd net683 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[36]  \la_data_in_mprj_bar[36]\ vssd vssd vccd vccd net684 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[37]  \la_data_in_mprj_bar[37]\ vssd vssd vccd vccd net685 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[38]  \la_data_in_mprj_bar[38]\ vssd vssd vccd vccd net686 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[39]  \la_data_in_mprj_bar[39]\ vssd vssd vccd vccd net687 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[3]  \la_data_in_mprj_bar[3]\ vssd vssd vccd vccd net688 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[40]  \la_data_in_mprj_bar[40]\ vssd vssd vccd vccd net689 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[41]  \la_data_in_mprj_bar[41]\ vssd vssd vccd vccd net690 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[42]  \la_data_in_mprj_bar[42]\ vssd vssd vccd vccd net691 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[43]  \la_data_in_mprj_bar[43]\ vssd vssd vccd vccd net692 sky130_fd_sc_hd__inv_2
X\user_to_mprj_in_buffers[44]  \la_data_in_mprj_bar[44]\ vssd vssd vccd vccd net693 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[45]  \la_data_in_mprj_bar[45]\ vssd vssd vccd vccd net694 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[46]  \la_data_in_mprj_bar[46]\ vssd vssd vccd vccd net695 sky130_fd_sc_hd__inv_2
X\user_to_mprj_in_buffers[47]  \la_data_in_mprj_bar[47]\ vssd vssd vccd vccd net696 sky130_fd_sc_hd__inv_2
X\user_to_mprj_in_buffers[48]  \la_data_in_mprj_bar[48]\ vssd vssd vccd vccd net697 sky130_fd_sc_hd__inv_2
X\user_to_mprj_in_buffers[49]  \la_data_in_mprj_bar[49]\ vssd vssd vccd vccd net698 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[4]  \la_data_in_mprj_bar[4]\ vssd vssd vccd vccd net699 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[50]  \la_data_in_mprj_bar[50]\ vssd vssd vccd vccd net700 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[51]  \la_data_in_mprj_bar[51]\ vssd vssd vccd vccd net701 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[52]  \la_data_in_mprj_bar[52]\ vssd vssd vccd vccd net702 sky130_fd_sc_hd__inv_2
X\user_to_mprj_in_buffers[53]  \la_data_in_mprj_bar[53]\ vssd vssd vccd vccd net703 sky130_fd_sc_hd__inv_2
X\user_to_mprj_in_buffers[54]  \la_data_in_mprj_bar[54]\ vssd vssd vccd vccd net704 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[55]  \la_data_in_mprj_bar[55]\ vssd vssd vccd vccd net705 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[56]  \la_data_in_mprj_bar[56]\ vssd vssd vccd vccd net706 sky130_fd_sc_hd__inv_2
X\user_to_mprj_in_buffers[57]  \la_data_in_mprj_bar[57]\ vssd vssd vccd vccd net707 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[58]  \la_data_in_mprj_bar[58]\ vssd vssd vccd vccd net708 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[59]  \la_data_in_mprj_bar[59]\ vssd vssd vccd vccd net709 sky130_fd_sc_hd__inv_2
X\user_to_mprj_in_buffers[5]  \la_data_in_mprj_bar[5]\ vssd vssd vccd vccd net710 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[60]  \la_data_in_mprj_bar[60]\ vssd vssd vccd vccd net711 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[61]  \la_data_in_mprj_bar[61]\ vssd vssd vccd vccd net712 sky130_fd_sc_hd__clkinv_2
X\user_to_mprj_in_buffers[62]  \la_data_in_mprj_bar[62]\ vssd vssd vccd vccd net713 sky130_fd_sc_hd__inv_2
X\user_to_mprj_in_buffers[63]  \la_data_in_mprj_bar[63]\ vssd vssd vccd vccd net714 sky130_fd_sc_hd__inv_2
X\user_to_mprj_in_buffers[64]  \la_data_in_mprj_bar[64]\ vssd vssd vccd vccd net715 sky130_fd_sc_hd__inv_2
X\user_to_mprj_in_buffers[65]  \la_data_in_mprj_bar[65]\ vssd vssd vccd vccd net716 sky130_fd_sc_hd__clkinv_2
X\user_to_mprj_in_buffers[66]  \la_data_in_mprj_bar[66]\ vssd vssd vccd vccd net717 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[67]  \la_data_in_mprj_bar[67]\ vssd vssd vccd vccd net718 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[68]  \la_data_in_mprj_bar[68]\ vssd vssd vccd vccd net719 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[69]  \la_data_in_mprj_bar[69]\ vssd vssd vccd vccd net720 sky130_fd_sc_hd__inv_2
X\user_to_mprj_in_buffers[6]  \la_data_in_mprj_bar[6]\ vssd vssd vccd vccd net721 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[70]  \la_data_in_mprj_bar[70]\ vssd vssd vccd vccd net722 sky130_fd_sc_hd__inv_2
X\user_to_mprj_in_buffers[71]  \la_data_in_mprj_bar[71]\ vssd vssd vccd vccd net723 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[72]  \la_data_in_mprj_bar[72]\ vssd vssd vccd vccd net724 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[73]  \la_data_in_mprj_bar[73]\ vssd vssd vccd vccd net725 sky130_fd_sc_hd__inv_2
X\user_to_mprj_in_buffers[74]  \la_data_in_mprj_bar[74]\ vssd vssd vccd vccd net726 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[75]  \la_data_in_mprj_bar[75]\ vssd vssd vccd vccd net727 sky130_fd_sc_hd__inv_2
X\user_to_mprj_in_buffers[76]  \la_data_in_mprj_bar[76]\ vssd vssd vccd vccd net728 sky130_fd_sc_hd__inv_2
X\user_to_mprj_in_buffers[77]  \la_data_in_mprj_bar[77]\ vssd vssd vccd vccd net729 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[78]  \la_data_in_mprj_bar[78]\ vssd vssd vccd vccd net730 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[79]  \la_data_in_mprj_bar[79]\ vssd vssd vccd vccd net731 sky130_fd_sc_hd__inv_2
X\user_to_mprj_in_buffers[7]  \la_data_in_mprj_bar[7]\ vssd vssd vccd vccd net732 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[80]  \la_data_in_mprj_bar[80]\ vssd vssd vccd vccd net733 sky130_fd_sc_hd__inv_2
X\user_to_mprj_in_buffers[81]  \la_data_in_mprj_bar[81]\ vssd vssd vccd vccd net734 sky130_fd_sc_hd__inv_2
X\user_to_mprj_in_buffers[82]  \la_data_in_mprj_bar[82]\ vssd vssd vccd vccd net735 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[83]  \la_data_in_mprj_bar[83]\ vssd vssd vccd vccd net736 sky130_fd_sc_hd__inv_2
X\user_to_mprj_in_buffers[84]  \la_data_in_mprj_bar[84]\ vssd vssd vccd vccd net737 sky130_fd_sc_hd__inv_2
X\user_to_mprj_in_buffers[85]  \la_data_in_mprj_bar[85]\ vssd vssd vccd vccd net738 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[86]  \la_data_in_mprj_bar[86]\ vssd vssd vccd vccd net739 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[87]  \la_data_in_mprj_bar[87]\ vssd vssd vccd vccd net740 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[88]  \la_data_in_mprj_bar[88]\ vssd vssd vccd vccd net741 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[89]  \la_data_in_mprj_bar[89]\ vssd vssd vccd vccd net742 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[8]  \la_data_in_mprj_bar[8]\ vssd vssd vccd vccd net743 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[90]  \la_data_in_mprj_bar[90]\ vssd vssd vccd vccd net744 sky130_fd_sc_hd__inv_2
X\user_to_mprj_in_buffers[91]  \la_data_in_mprj_bar[91]\ vssd vssd vccd vccd net745 sky130_fd_sc_hd__inv_2
X\user_to_mprj_in_buffers[92]  \la_data_in_mprj_bar[92]\ vssd vssd vccd vccd net746 sky130_fd_sc_hd__inv_2
X\user_to_mprj_in_buffers[93]  \la_data_in_mprj_bar[93]\ vssd vssd vccd vccd net747 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[94]  \la_data_in_mprj_bar[94]\ vssd vssd vccd vccd net748 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[95]  \la_data_in_mprj_bar[95]\ vssd vssd vccd vccd net749 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[96]  \la_data_in_mprj_bar[96]\ vssd vssd vccd vccd net750 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[97]  \la_data_in_mprj_bar[97]\ vssd vssd vccd vccd net751 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[98]  \la_data_in_mprj_bar[98]\ vssd vssd vccd vccd net752 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[99]  \la_data_in_mprj_bar[99]\ vssd vssd vccd vccd net753 sky130_fd_sc_hd__clkinv_4
X\user_to_mprj_in_buffers[9]  \la_data_in_mprj_bar[9]\ vssd vssd vccd vccd net754 sky130_fd_sc_hd__inv_6
X\user_to_mprj_in_ena_buf[0]  net260 \mprj_logic1[330]\ vssd vssd vccd vccd \la_data_in_enable[0]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[100]  net261 \mprj_logic1[430]\ vssd vssd vccd vccd \la_data_in_enable[100]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[101]  net262 \mprj_logic1[431]\ vssd vssd vccd vccd \la_data_in_enable[101]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[102]  net263 \mprj_logic1[432]\ vssd vssd vccd vccd \la_data_in_enable[102]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[103]  net264 \mprj_logic1[433]\ vssd vssd vccd vccd \la_data_in_enable[103]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[104]  net265 \mprj_logic1[434]\ vssd vssd vccd vccd \la_data_in_enable[104]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[105]  net266 \mprj_logic1[435]\ vssd vssd vccd vccd \la_data_in_enable[105]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[106]  net267 \mprj_logic1[436]\ vssd vssd vccd vccd \la_data_in_enable[106]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[107]  net268 \mprj_logic1[437]\ vssd vssd vccd vccd \la_data_in_enable[107]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[108]  net269 \mprj_logic1[438]\ vssd vssd vccd vccd \la_data_in_enable[108]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[109]  net270 \mprj_logic1[439]\ vssd vssd vccd vccd \la_data_in_enable[109]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[10]  net271 \mprj_logic1[340]\ vssd vssd vccd vccd \la_data_in_enable[10]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[110]  net272 \mprj_logic1[440]\ vssd vssd vccd vccd \la_data_in_enable[110]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[111]  net273 \mprj_logic1[441]\ vssd vssd vccd vccd \la_data_in_enable[111]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[112]  net274 \mprj_logic1[442]\ vssd vssd vccd vccd \la_data_in_enable[112]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[113]  net275 \mprj_logic1[443]\ vssd vssd vccd vccd \la_data_in_enable[113]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[114]  net276 \mprj_logic1[444]\ vssd vssd vccd vccd \la_data_in_enable[114]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[115]  net277 \mprj_logic1[445]\ vssd vssd vccd vccd \la_data_in_enable[115]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[116]  net278 \mprj_logic1[446]\ vssd vssd vccd vccd \la_data_in_enable[116]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[117]  net279 \mprj_logic1[447]\ vssd vssd vccd vccd \la_data_in_enable[117]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[118]  net280 \mprj_logic1[448]\ vssd vssd vccd vccd \la_data_in_enable[118]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[119]  net281 \mprj_logic1[449]\ vssd vssd vccd vccd \la_data_in_enable[119]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[11]  net282 \mprj_logic1[341]\ vssd vssd vccd vccd \la_data_in_enable[11]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[120]  net283 \mprj_logic1[450]\ vssd vssd vccd vccd \la_data_in_enable[120]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[121]  net284 \mprj_logic1[451]\ vssd vssd vccd vccd \la_data_in_enable[121]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[122]  net285 \mprj_logic1[452]\ vssd vssd vccd vccd \la_data_in_enable[122]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[123]  net286 \mprj_logic1[453]\ vssd vssd vccd vccd \la_data_in_enable[123]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[124]  net287 \mprj_logic1[454]\ vssd vssd vccd vccd \la_data_in_enable[124]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[125]  net288 \mprj_logic1[455]\ vssd vssd vccd vccd \la_data_in_enable[125]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[126]  net289 \mprj_logic1[456]\ vssd vssd vccd vccd \la_data_in_enable[126]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[127]  net290 \mprj_logic1[457]\ vssd vssd vccd vccd \la_data_in_enable[127]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[12]  net291 \mprj_logic1[342]\ vssd vssd vccd vccd \la_data_in_enable[12]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[13]  net292 \mprj_logic1[343]\ vssd vssd vccd vccd \la_data_in_enable[13]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[14]  net293 \mprj_logic1[344]\ vssd vssd vccd vccd \la_data_in_enable[14]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[15]  net294 \mprj_logic1[345]\ vssd vssd vccd vccd \la_data_in_enable[15]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[16]  net295 \mprj_logic1[346]\ vssd vssd vccd vccd \la_data_in_enable[16]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[17]  net296 \mprj_logic1[347]\ vssd vssd vccd vccd \la_data_in_enable[17]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[18]  net297 \mprj_logic1[348]\ vssd vssd vccd vccd \la_data_in_enable[18]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[19]  net298 \mprj_logic1[349]\ vssd vssd vccd vccd \la_data_in_enable[19]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[1]  net299 \mprj_logic1[331]\ vssd vssd vccd vccd \la_data_in_enable[1]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[20]  net300 \mprj_logic1[350]\ vssd vssd vccd vccd \la_data_in_enable[20]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[21]  net301 \mprj_logic1[351]\ vssd vssd vccd vccd \la_data_in_enable[21]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[22]  net302 \mprj_logic1[352]\ vssd vssd vccd vccd \la_data_in_enable[22]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[23]  net303 \mprj_logic1[353]\ vssd vssd vccd vccd \la_data_in_enable[23]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[24]  net304 \mprj_logic1[354]\ vssd vssd vccd vccd \la_data_in_enable[24]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[25]  net305 \mprj_logic1[355]\ vssd vssd vccd vccd \la_data_in_enable[25]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[26]  net306 \mprj_logic1[356]\ vssd vssd vccd vccd \la_data_in_enable[26]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[27]  net307 \mprj_logic1[357]\ vssd vssd vccd vccd \la_data_in_enable[27]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[28]  net308 \mprj_logic1[358]\ vssd vssd vccd vccd \la_data_in_enable[28]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[29]  net309 \mprj_logic1[359]\ vssd vssd vccd vccd \la_data_in_enable[29]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[2]  net310 \mprj_logic1[332]\ vssd vssd vccd vccd \la_data_in_enable[2]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[30]  net311 \mprj_logic1[360]\ vssd vssd vccd vccd \la_data_in_enable[30]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[31]  net312 \mprj_logic1[361]\ vssd vssd vccd vccd \la_data_in_enable[31]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[32]  net313 \mprj_logic1[362]\ vssd vssd vccd vccd \la_data_in_enable[32]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[33]  net314 \mprj_logic1[363]\ vssd vssd vccd vccd \la_data_in_enable[33]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[34]  net315 \mprj_logic1[364]\ vssd vssd vccd vccd \la_data_in_enable[34]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[35]  net316 \mprj_logic1[365]\ vssd vssd vccd vccd \la_data_in_enable[35]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[36]  net317 \mprj_logic1[366]\ vssd vssd vccd vccd \la_data_in_enable[36]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[37]  net318 \mprj_logic1[367]\ vssd vssd vccd vccd \la_data_in_enable[37]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[38]  net319 \mprj_logic1[368]\ vssd vssd vccd vccd \la_data_in_enable[38]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[39]  net320 \mprj_logic1[369]\ vssd vssd vccd vccd \la_data_in_enable[39]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[3]  net321 \mprj_logic1[333]\ vssd vssd vccd vccd \la_data_in_enable[3]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[40]  net322 \mprj_logic1[370]\ vssd vssd vccd vccd \la_data_in_enable[40]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[41]  net323 \mprj_logic1[371]\ vssd vssd vccd vccd \la_data_in_enable[41]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[42]  net324 \mprj_logic1[372]\ vssd vssd vccd vccd \la_data_in_enable[42]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[43]  net325 \mprj_logic1[373]\ vssd vssd vccd vccd \la_data_in_enable[43]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[44]  net326 \mprj_logic1[374]\ vssd vssd vccd vccd \la_data_in_enable[44]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[45]  net327 \mprj_logic1[375]\ vssd vssd vccd vccd \la_data_in_enable[45]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[46]  net328 \mprj_logic1[376]\ vssd vssd vccd vccd \la_data_in_enable[46]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[47]  net329 \mprj_logic1[377]\ vssd vssd vccd vccd \la_data_in_enable[47]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[48]  net330 \mprj_logic1[378]\ vssd vssd vccd vccd \la_data_in_enable[48]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[49]  net331 \mprj_logic1[379]\ vssd vssd vccd vccd \la_data_in_enable[49]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[4]  net332 \mprj_logic1[334]\ vssd vssd vccd vccd \la_data_in_enable[4]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[50]  net333 \mprj_logic1[380]\ vssd vssd vccd vccd \la_data_in_enable[50]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[51]  net334 \mprj_logic1[381]\ vssd vssd vccd vccd \la_data_in_enable[51]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[52]  net335 \mprj_logic1[382]\ vssd vssd vccd vccd \la_data_in_enable[52]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[53]  net336 \mprj_logic1[383]\ vssd vssd vccd vccd \la_data_in_enable[53]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[54]  net337 \mprj_logic1[384]\ vssd vssd vccd vccd \la_data_in_enable[54]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[55]  net338 \mprj_logic1[385]\ vssd vssd vccd vccd \la_data_in_enable[55]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[56]  net339 \mprj_logic1[386]\ vssd vssd vccd vccd \la_data_in_enable[56]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[57]  net340 \mprj_logic1[387]\ vssd vssd vccd vccd \la_data_in_enable[57]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[58]  net341 \mprj_logic1[388]\ vssd vssd vccd vccd \la_data_in_enable[58]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[59]  net342 \mprj_logic1[389]\ vssd vssd vccd vccd \la_data_in_enable[59]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[5]  net343 \mprj_logic1[335]\ vssd vssd vccd vccd \la_data_in_enable[5]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[60]  net344 \mprj_logic1[390]\ vssd vssd vccd vccd \la_data_in_enable[60]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[61]  net345 \mprj_logic1[391]\ vssd vssd vccd vccd \la_data_in_enable[61]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[62]  net346 \mprj_logic1[392]\ vssd vssd vccd vccd \la_data_in_enable[62]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[63]  net347 \mprj_logic1[393]\ vssd vssd vccd vccd \la_data_in_enable[63]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[64]  net348 \mprj_logic1[394]\ vssd vssd vccd vccd \la_data_in_enable[64]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[65]  net349 \mprj_logic1[395]\ vssd vssd vccd vccd \la_data_in_enable[65]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[66]  net350 \mprj_logic1[396]\ vssd vssd vccd vccd \la_data_in_enable[66]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[67]  net351 \mprj_logic1[397]\ vssd vssd vccd vccd \la_data_in_enable[67]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[68]  net352 \mprj_logic1[398]\ vssd vssd vccd vccd \la_data_in_enable[68]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[69]  net353 \mprj_logic1[399]\ vssd vssd vccd vccd \la_data_in_enable[69]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[6]  net354 \mprj_logic1[336]\ vssd vssd vccd vccd \la_data_in_enable[6]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[70]  net355 \mprj_logic1[400]\ vssd vssd vccd vccd \la_data_in_enable[70]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[71]  net356 \mprj_logic1[401]\ vssd vssd vccd vccd \la_data_in_enable[71]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[72]  net357 \mprj_logic1[402]\ vssd vssd vccd vccd \la_data_in_enable[72]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[73]  net358 \mprj_logic1[403]\ vssd vssd vccd vccd \la_data_in_enable[73]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[74]  net359 \mprj_logic1[404]\ vssd vssd vccd vccd \la_data_in_enable[74]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[75]  net360 \mprj_logic1[405]\ vssd vssd vccd vccd \la_data_in_enable[75]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[76]  net361 \mprj_logic1[406]\ vssd vssd vccd vccd \la_data_in_enable[76]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[77]  net362 \mprj_logic1[407]\ vssd vssd vccd vccd \la_data_in_enable[77]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[78]  net363 \mprj_logic1[408]\ vssd vssd vccd vccd \la_data_in_enable[78]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[79]  net364 \mprj_logic1[409]\ vssd vssd vccd vccd \la_data_in_enable[79]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[7]  net365 \mprj_logic1[337]\ vssd vssd vccd vccd \la_data_in_enable[7]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[80]  net366 \mprj_logic1[410]\ vssd vssd vccd vccd \la_data_in_enable[80]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[81]  net367 \mprj_logic1[411]\ vssd vssd vccd vccd \la_data_in_enable[81]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[82]  net368 \mprj_logic1[412]\ vssd vssd vccd vccd \la_data_in_enable[82]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[83]  net369 \mprj_logic1[413]\ vssd vssd vccd vccd \la_data_in_enable[83]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[84]  net370 \mprj_logic1[414]\ vssd vssd vccd vccd \la_data_in_enable[84]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[85]  net371 \mprj_logic1[415]\ vssd vssd vccd vccd \la_data_in_enable[85]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[86]  net372 \mprj_logic1[416]\ vssd vssd vccd vccd \la_data_in_enable[86]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[87]  net373 \mprj_logic1[417]\ vssd vssd vccd vccd \la_data_in_enable[87]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[88]  net374 \mprj_logic1[418]\ vssd vssd vccd vccd \la_data_in_enable[88]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[89]  net375 \mprj_logic1[419]\ vssd vssd vccd vccd \la_data_in_enable[89]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[8]  net376 \mprj_logic1[338]\ vssd vssd vccd vccd \la_data_in_enable[8]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[90]  net377 \mprj_logic1[420]\ vssd vssd vccd vccd \la_data_in_enable[90]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[91]  net378 \mprj_logic1[421]\ vssd vssd vccd vccd \la_data_in_enable[91]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[92]  net379 \mprj_logic1[422]\ vssd vssd vccd vccd \la_data_in_enable[92]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[93]  net380 \mprj_logic1[423]\ vssd vssd vccd vccd \la_data_in_enable[93]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[94]  net381 \mprj_logic1[424]\ vssd vssd vccd vccd \la_data_in_enable[94]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[95]  net382 \mprj_logic1[425]\ vssd vssd vccd vccd \la_data_in_enable[95]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[96]  net383 \mprj_logic1[426]\ vssd vssd vccd vccd \la_data_in_enable[96]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[97]  net384 \mprj_logic1[427]\ vssd vssd vccd vccd \la_data_in_enable[97]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[98]  net385 \mprj_logic1[428]\ vssd vssd vccd vccd \la_data_in_enable[98]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[99]  net386 \mprj_logic1[429]\ vssd vssd vccd vccd \la_data_in_enable[99]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_ena_buf[9]  net387 \mprj_logic1[339]\ vssd vssd vccd vccd \la_data_in_enable[9]\ sky130_fd_sc_hd__and2_1
X\user_to_mprj_in_gates[0]  net4 \la_data_in_enable[0]\ vssd vssd vccd vccd \la_data_in_mprj_bar[0]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[100]  net5 \la_data_in_enable[100]\ vssd vssd vccd vccd \la_data_in_mprj_bar[100]\ sky130_fd_sc_hd__nand2_2
X\user_to_mprj_in_gates[101]  net6 \la_data_in_enable[101]\ vssd vssd vccd vccd \la_data_in_mprj_bar[101]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[102]  net7 \la_data_in_enable[102]\ vssd vssd vccd vccd \la_data_in_mprj_bar[102]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[103]  net8 \la_data_in_enable[103]\ vssd vssd vccd vccd \la_data_in_mprj_bar[103]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[104]  net9 \la_data_in_enable[104]\ vssd vssd vccd vccd \la_data_in_mprj_bar[104]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[105]  net10 \la_data_in_enable[105]\ vssd vssd vccd vccd \la_data_in_mprj_bar[105]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[106]  net11 \la_data_in_enable[106]\ vssd vssd vccd vccd \la_data_in_mprj_bar[106]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[107]  net12 \la_data_in_enable[107]\ vssd vssd vccd vccd \la_data_in_mprj_bar[107]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[108]  net13 \la_data_in_enable[108]\ vssd vssd vccd vccd \la_data_in_mprj_bar[108]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[109]  net14 \la_data_in_enable[109]\ vssd vssd vccd vccd \la_data_in_mprj_bar[109]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[10]  net15 \la_data_in_enable[10]\ vssd vssd vccd vccd \la_data_in_mprj_bar[10]\ sky130_fd_sc_hd__nand2_2
X\user_to_mprj_in_gates[110]  net16 \la_data_in_enable[110]\ vssd vssd vccd vccd \la_data_in_mprj_bar[110]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[111]  net17 \la_data_in_enable[111]\ vssd vssd vccd vccd \la_data_in_mprj_bar[111]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[112]  net18 \la_data_in_enable[112]\ vssd vssd vccd vccd \la_data_in_mprj_bar[112]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[113]  net19 \la_data_in_enable[113]\ vssd vssd vccd vccd \la_data_in_mprj_bar[113]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[114]  net20 \la_data_in_enable[114]\ vssd vssd vccd vccd \la_data_in_mprj_bar[114]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[115]  net21 \la_data_in_enable[115]\ vssd vssd vccd vccd \la_data_in_mprj_bar[115]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[116]  net22 \la_data_in_enable[116]\ vssd vssd vccd vccd \la_data_in_mprj_bar[116]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[117]  net23 \la_data_in_enable[117]\ vssd vssd vccd vccd \la_data_in_mprj_bar[117]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[118]  net24 \la_data_in_enable[118]\ vssd vssd vccd vccd \la_data_in_mprj_bar[118]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[119]  net25 \la_data_in_enable[119]\ vssd vssd vccd vccd \la_data_in_mprj_bar[119]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[11]  net26 \la_data_in_enable[11]\ vssd vssd vccd vccd \la_data_in_mprj_bar[11]\ sky130_fd_sc_hd__nand2_2
X\user_to_mprj_in_gates[120]  net27 \la_data_in_enable[120]\ vssd vssd vccd vccd \la_data_in_mprj_bar[120]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[121]  net28 \la_data_in_enable[121]\ vssd vssd vccd vccd \la_data_in_mprj_bar[121]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[122]  net29 \la_data_in_enable[122]\ vssd vssd vccd vccd \la_data_in_mprj_bar[122]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[123]  net30 \la_data_in_enable[123]\ vssd vssd vccd vccd \la_data_in_mprj_bar[123]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[124]  net31 \la_data_in_enable[124]\ vssd vssd vccd vccd \la_data_in_mprj_bar[124]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[125]  net32 \la_data_in_enable[125]\ vssd vssd vccd vccd \la_data_in_mprj_bar[125]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[126]  net33 \la_data_in_enable[126]\ vssd vssd vccd vccd \la_data_in_mprj_bar[126]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[127]  net34 \la_data_in_enable[127]\ vssd vssd vccd vccd \la_data_in_mprj_bar[127]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[12]  net35 \la_data_in_enable[12]\ vssd vssd vccd vccd \la_data_in_mprj_bar[12]\ sky130_fd_sc_hd__nand2_2
X\user_to_mprj_in_gates[13]  net36 \la_data_in_enable[13]\ vssd vssd vccd vccd \la_data_in_mprj_bar[13]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[14]  net37 \la_data_in_enable[14]\ vssd vssd vccd vccd \la_data_in_mprj_bar[14]\ sky130_fd_sc_hd__nand2_2
X\user_to_mprj_in_gates[15]  net38 \la_data_in_enable[15]\ vssd vssd vccd vccd \la_data_in_mprj_bar[15]\ sky130_fd_sc_hd__nand2_2
X\user_to_mprj_in_gates[16]  net39 \la_data_in_enable[16]\ vssd vssd vccd vccd \la_data_in_mprj_bar[16]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[17]  net40 \la_data_in_enable[17]\ vssd vssd vccd vccd \la_data_in_mprj_bar[17]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[18]  net41 \la_data_in_enable[18]\ vssd vssd vccd vccd \la_data_in_mprj_bar[18]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[19]  net42 \la_data_in_enable[19]\ vssd vssd vccd vccd \la_data_in_mprj_bar[19]\ sky130_fd_sc_hd__nand2_2
X\user_to_mprj_in_gates[1]  net43 \la_data_in_enable[1]\ vssd vssd vccd vccd \la_data_in_mprj_bar[1]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[20]  net44 \la_data_in_enable[20]\ vssd vssd vccd vccd \la_data_in_mprj_bar[20]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[21]  net45 \la_data_in_enable[21]\ vssd vssd vccd vccd \la_data_in_mprj_bar[21]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[22]  net46 \la_data_in_enable[22]\ vssd vssd vccd vccd \la_data_in_mprj_bar[22]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[23]  net47 \la_data_in_enable[23]\ vssd vssd vccd vccd \la_data_in_mprj_bar[23]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[24]  net48 \la_data_in_enable[24]\ vssd vssd vccd vccd \la_data_in_mprj_bar[24]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[25]  net49 \la_data_in_enable[25]\ vssd vssd vccd vccd \la_data_in_mprj_bar[25]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[26]  net50 \la_data_in_enable[26]\ vssd vssd vccd vccd \la_data_in_mprj_bar[26]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[27]  net51 \la_data_in_enable[27]\ vssd vssd vccd vccd \la_data_in_mprj_bar[27]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[28]  net52 \la_data_in_enable[28]\ vssd vssd vccd vccd \la_data_in_mprj_bar[28]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[29]  net53 \la_data_in_enable[29]\ vssd vssd vccd vccd \la_data_in_mprj_bar[29]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[2]  net54 \la_data_in_enable[2]\ vssd vssd vccd vccd \la_data_in_mprj_bar[2]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[30]  net55 \la_data_in_enable[30]\ vssd vssd vccd vccd \la_data_in_mprj_bar[30]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[31]  net56 \la_data_in_enable[31]\ vssd vssd vccd vccd \la_data_in_mprj_bar[31]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[32]  net57 \la_data_in_enable[32]\ vssd vssd vccd vccd \la_data_in_mprj_bar[32]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[33]  net58 \la_data_in_enable[33]\ vssd vssd vccd vccd \la_data_in_mprj_bar[33]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[34]  net59 \la_data_in_enable[34]\ vssd vssd vccd vccd \la_data_in_mprj_bar[34]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[35]  net60 \la_data_in_enable[35]\ vssd vssd vccd vccd \la_data_in_mprj_bar[35]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[36]  net61 \la_data_in_enable[36]\ vssd vssd vccd vccd \la_data_in_mprj_bar[36]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[37]  net62 \la_data_in_enable[37]\ vssd vssd vccd vccd \la_data_in_mprj_bar[37]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[38]  net63 \la_data_in_enable[38]\ vssd vssd vccd vccd \la_data_in_mprj_bar[38]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[39]  net64 \la_data_in_enable[39]\ vssd vssd vccd vccd \la_data_in_mprj_bar[39]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[3]  net65 \la_data_in_enable[3]\ vssd vssd vccd vccd \la_data_in_mprj_bar[3]\ sky130_fd_sc_hd__nand2_2
X\user_to_mprj_in_gates[40]  net66 \la_data_in_enable[40]\ vssd vssd vccd vccd \la_data_in_mprj_bar[40]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[41]  net67 \la_data_in_enable[41]\ vssd vssd vccd vccd \la_data_in_mprj_bar[41]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[42]  net68 \la_data_in_enable[42]\ vssd vssd vccd vccd \la_data_in_mprj_bar[42]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[43]  net69 \la_data_in_enable[43]\ vssd vssd vccd vccd \la_data_in_mprj_bar[43]\ sky130_fd_sc_hd__nand2_2
X\user_to_mprj_in_gates[44]  net70 \la_data_in_enable[44]\ vssd vssd vccd vccd \la_data_in_mprj_bar[44]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[45]  net71 \la_data_in_enable[45]\ vssd vssd vccd vccd \la_data_in_mprj_bar[45]\ sky130_fd_sc_hd__nand2_2
X\user_to_mprj_in_gates[46]  net72 \la_data_in_enable[46]\ vssd vssd vccd vccd \la_data_in_mprj_bar[46]\ sky130_fd_sc_hd__nand2_2
X\user_to_mprj_in_gates[47]  net73 \la_data_in_enable[47]\ vssd vssd vccd vccd \la_data_in_mprj_bar[47]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[48]  net74 \la_data_in_enable[48]\ vssd vssd vccd vccd \la_data_in_mprj_bar[48]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[49]  net75 \la_data_in_enable[49]\ vssd vssd vccd vccd \la_data_in_mprj_bar[49]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[4]  net76 \la_data_in_enable[4]\ vssd vssd vccd vccd \la_data_in_mprj_bar[4]\ sky130_fd_sc_hd__nand2_4
X\user_to_mprj_in_gates[50]  net77 \la_data_in_enable[50]\ vssd vssd vccd vccd \la_data_in_mprj_bar[50]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[51]  net78 \la_data_in_enable[51]\ vssd vssd vccd vccd \la_data_in_mprj_bar[51]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[52]  net79 \la_data_in_enable[52]\ vssd vssd vccd vccd \la_data_in_mprj_bar[52]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[53]  net80 \la_data_in_enable[53]\ vssd vssd vccd vccd \la_data_in_mprj_bar[53]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[54]  net81 \la_data_in_enable[54]\ vssd vssd vccd vccd \la_data_in_mprj_bar[54]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[55]  net82 \la_data_in_enable[55]\ vssd vssd vccd vccd \la_data_in_mprj_bar[55]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[56]  net83 \la_data_in_enable[56]\ vssd vssd vccd vccd \la_data_in_mprj_bar[56]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[57]  net84 \la_data_in_enable[57]\ vssd vssd vccd vccd \la_data_in_mprj_bar[57]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[58]  net85 \la_data_in_enable[58]\ vssd vssd vccd vccd \la_data_in_mprj_bar[58]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[59]  net86 \la_data_in_enable[59]\ vssd vssd vccd vccd \la_data_in_mprj_bar[59]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[5]  net87 \la_data_in_enable[5]\ vssd vssd vccd vccd \la_data_in_mprj_bar[5]\ sky130_fd_sc_hd__nand2_4
X\user_to_mprj_in_gates[60]  net88 \la_data_in_enable[60]\ vssd vssd vccd vccd \la_data_in_mprj_bar[60]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[61]  net89 \la_data_in_enable[61]\ vssd vssd vccd vccd \la_data_in_mprj_bar[61]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[62]  net90 \la_data_in_enable[62]\ vssd vssd vccd vccd \la_data_in_mprj_bar[62]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[63]  net91 \la_data_in_enable[63]\ vssd vssd vccd vccd \la_data_in_mprj_bar[63]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[64]  net92 \la_data_in_enable[64]\ vssd vssd vccd vccd \la_data_in_mprj_bar[64]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[65]  net93 \la_data_in_enable[65]\ vssd vssd vccd vccd \la_data_in_mprj_bar[65]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[66]  net94 \la_data_in_enable[66]\ vssd vssd vccd vccd \la_data_in_mprj_bar[66]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[67]  net95 \la_data_in_enable[67]\ vssd vssd vccd vccd \la_data_in_mprj_bar[67]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[68]  net96 \la_data_in_enable[68]\ vssd vssd vccd vccd \la_data_in_mprj_bar[68]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[69]  net97 \la_data_in_enable[69]\ vssd vssd vccd vccd \la_data_in_mprj_bar[69]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[6]  net98 \la_data_in_enable[6]\ vssd vssd vccd vccd \la_data_in_mprj_bar[6]\ sky130_fd_sc_hd__nand2_4
X\user_to_mprj_in_gates[70]  net99 \la_data_in_enable[70]\ vssd vssd vccd vccd \la_data_in_mprj_bar[70]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[71]  net100 \la_data_in_enable[71]\ vssd vssd vccd vccd \la_data_in_mprj_bar[71]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[72]  net101 \la_data_in_enable[72]\ vssd vssd vccd vccd \la_data_in_mprj_bar[72]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[73]  net102 \la_data_in_enable[73]\ vssd vssd vccd vccd \la_data_in_mprj_bar[73]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[74]  net103 \la_data_in_enable[74]\ vssd vssd vccd vccd \la_data_in_mprj_bar[74]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[75]  net104 \la_data_in_enable[75]\ vssd vssd vccd vccd \la_data_in_mprj_bar[75]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[76]  net105 \la_data_in_enable[76]\ vssd vssd vccd vccd \la_data_in_mprj_bar[76]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[77]  net106 \la_data_in_enable[77]\ vssd vssd vccd vccd \la_data_in_mprj_bar[77]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[78]  net107 \la_data_in_enable[78]\ vssd vssd vccd vccd \la_data_in_mprj_bar[78]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[79]  net108 \la_data_in_enable[79]\ vssd vssd vccd vccd \la_data_in_mprj_bar[79]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[7]  net109 \la_data_in_enable[7]\ vssd vssd vccd vccd \la_data_in_mprj_bar[7]\ sky130_fd_sc_hd__nand2_4
X\user_to_mprj_in_gates[80]  net110 \la_data_in_enable[80]\ vssd vssd vccd vccd \la_data_in_mprj_bar[80]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[81]  net111 \la_data_in_enable[81]\ vssd vssd vccd vccd \la_data_in_mprj_bar[81]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[82]  net112 \la_data_in_enable[82]\ vssd vssd vccd vccd \la_data_in_mprj_bar[82]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[83]  net113 \la_data_in_enable[83]\ vssd vssd vccd vccd \la_data_in_mprj_bar[83]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[84]  net114 \la_data_in_enable[84]\ vssd vssd vccd vccd \la_data_in_mprj_bar[84]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[85]  net115 \la_data_in_enable[85]\ vssd vssd vccd vccd \la_data_in_mprj_bar[85]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[86]  net116 \la_data_in_enable[86]\ vssd vssd vccd vccd \la_data_in_mprj_bar[86]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[87]  net117 \la_data_in_enable[87]\ vssd vssd vccd vccd \la_data_in_mprj_bar[87]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[88]  net118 \la_data_in_enable[88]\ vssd vssd vccd vccd \la_data_in_mprj_bar[88]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[89]  net119 \la_data_in_enable[89]\ vssd vssd vccd vccd \la_data_in_mprj_bar[89]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[8]  net120 \la_data_in_enable[8]\ vssd vssd vccd vccd \la_data_in_mprj_bar[8]\ sky130_fd_sc_hd__nand2_4
X\user_to_mprj_in_gates[90]  net121 \la_data_in_enable[90]\ vssd vssd vccd vccd \la_data_in_mprj_bar[90]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[91]  net122 \la_data_in_enable[91]\ vssd vssd vccd vccd \la_data_in_mprj_bar[91]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[92]  net123 \la_data_in_enable[92]\ vssd vssd vccd vccd \la_data_in_mprj_bar[92]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[93]  net124 \la_data_in_enable[93]\ vssd vssd vccd vccd \la_data_in_mprj_bar[93]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[94]  net125 \la_data_in_enable[94]\ vssd vssd vccd vccd \la_data_in_mprj_bar[94]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[95]  net126 \la_data_in_enable[95]\ vssd vssd vccd vccd \la_data_in_mprj_bar[95]\ sky130_fd_sc_hd__nand2_2
X\user_to_mprj_in_gates[96]  net127 \la_data_in_enable[96]\ vssd vssd vccd vccd \la_data_in_mprj_bar[96]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[97]  net128 \la_data_in_enable[97]\ vssd vssd vccd vccd \la_data_in_mprj_bar[97]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[98]  net129 \la_data_in_enable[98]\ vssd vssd vccd vccd \la_data_in_mprj_bar[98]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[99]  net130 \la_data_in_enable[99]\ vssd vssd vccd vccd \la_data_in_mprj_bar[99]\ sky130_fd_sc_hd__nand2_1
X\user_to_mprj_in_gates[9]  net131 \la_data_in_enable[9]\ vssd vssd vccd vccd \la_data_in_mprj_bar[9]\ sky130_fd_sc_hd__nand2_4
X\user_to_mprj_oen_buffers[0]  _201_ \mprj_logic1[202]\ vssd vssd vccd vccd la_oenb_core[0] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[100]  _202_ \mprj_logic1[302]\ vssd vssd vccd vccd la_oenb_core[100] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[101]  _203_ \mprj_logic1[303]\ vssd vssd vccd vccd la_oenb_core[101] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[102]  _204_ \mprj_logic1[304]\ vssd vssd vccd vccd la_oenb_core[102] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[103]  _205_ \mprj_logic1[305]\ vssd vssd vccd vccd la_oenb_core[103] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[104]  _206_ \mprj_logic1[306]\ vssd vssd vccd vccd la_oenb_core[104] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[105]  _207_ \mprj_logic1[307]\ vssd vssd vccd vccd la_oenb_core[105] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[106]  _208_ \mprj_logic1[308]\ vssd vssd vccd vccd la_oenb_core[106] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[107]  _209_ \mprj_logic1[309]\ vssd vssd vccd vccd la_oenb_core[107] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[108]  _210_ \mprj_logic1[310]\ vssd vssd vccd vccd la_oenb_core[108] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[109]  _211_ \mprj_logic1[311]\ vssd vssd vccd vccd la_oenb_core[109] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[10]  _212_ \mprj_logic1[212]\ vssd vssd vccd vccd la_oenb_core[10] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[110]  _213_ \mprj_logic1[312]\ vssd vssd vccd vccd la_oenb_core[110] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[111]  _214_ \mprj_logic1[313]\ vssd vssd vccd vccd la_oenb_core[111] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[112]  _215_ \mprj_logic1[314]\ vssd vssd vccd vccd la_oenb_core[112] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[113]  _216_ \mprj_logic1[315]\ vssd vssd vccd vccd la_oenb_core[113] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[114]  _217_ \mprj_logic1[316]\ vssd vssd vccd vccd la_oenb_core[114] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[115]  _218_ \mprj_logic1[317]\ vssd vssd vccd vccd la_oenb_core[115] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[116]  _219_ \mprj_logic1[318]\ vssd vssd vccd vccd la_oenb_core[116] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[117]  _220_ \mprj_logic1[319]\ vssd vssd vccd vccd la_oenb_core[117] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[118]  _221_ \mprj_logic1[320]\ vssd vssd vccd vccd la_oenb_core[118] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[119]  _222_ \mprj_logic1[321]\ vssd vssd vccd vccd la_oenb_core[119] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[11]  _223_ \mprj_logic1[213]\ vssd vssd vccd vccd la_oenb_core[11] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[120]  _224_ \mprj_logic1[322]\ vssd vssd vccd vccd la_oenb_core[120] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[121]  _225_ \mprj_logic1[323]\ vssd vssd vccd vccd la_oenb_core[121] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[122]  _226_ \mprj_logic1[324]\ vssd vssd vccd vccd la_oenb_core[122] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[123]  _227_ \mprj_logic1[325]\ vssd vssd vccd vccd la_oenb_core[123] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[124]  _228_ \mprj_logic1[326]\ vssd vssd vccd vccd la_oenb_core[124] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[125]  _229_ \mprj_logic1[327]\ vssd vssd vccd vccd la_oenb_core[125] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[126]  _230_ \mprj_logic1[328]\ vssd vssd vccd vccd la_oenb_core[126] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[127]  _231_ \mprj_logic1[329]\ vssd vssd vccd vccd la_oenb_core[127] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[12]  _232_ \mprj_logic1[214]\ vssd vssd vccd vccd la_oenb_core[12] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[13]  _233_ \mprj_logic1[215]\ vssd vssd vccd vccd la_oenb_core[13] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[14]  _234_ \mprj_logic1[216]\ vssd vssd vccd vccd la_oenb_core[14] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[15]  _235_ \mprj_logic1[217]\ vssd vssd vccd vccd la_oenb_core[15] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[16]  _236_ \mprj_logic1[218]\ vssd vssd vccd vccd la_oenb_core[16] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[17]  _237_ \mprj_logic1[219]\ vssd vssd vccd vccd la_oenb_core[17] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[18]  _238_ \mprj_logic1[220]\ vssd vssd vccd vccd la_oenb_core[18] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[19]  _239_ \mprj_logic1[221]\ vssd vssd vccd vccd la_oenb_core[19] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[1]  _240_ \mprj_logic1[203]\ vssd vssd vccd vccd la_oenb_core[1] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[20]  _241_ \mprj_logic1[222]\ vssd vssd vccd vccd la_oenb_core[20] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[21]  _242_ \mprj_logic1[223]\ vssd vssd vccd vccd la_oenb_core[21] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[22]  _243_ \mprj_logic1[224]\ vssd vssd vccd vccd la_oenb_core[22] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[23]  _244_ \mprj_logic1[225]\ vssd vssd vccd vccd la_oenb_core[23] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[24]  _245_ \mprj_logic1[226]\ vssd vssd vccd vccd la_oenb_core[24] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[25]  _246_ \mprj_logic1[227]\ vssd vssd vccd vccd la_oenb_core[25] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[26]  _247_ \mprj_logic1[228]\ vssd vssd vccd vccd la_oenb_core[26] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[27]  _248_ \mprj_logic1[229]\ vssd vssd vccd vccd la_oenb_core[27] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[28]  _249_ \mprj_logic1[230]\ vssd vssd vccd vccd la_oenb_core[28] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[29]  _250_ \mprj_logic1[231]\ vssd vssd vccd vccd la_oenb_core[29] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[2]  _251_ \mprj_logic1[204]\ vssd vssd vccd vccd la_oenb_core[2] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[30]  _252_ \mprj_logic1[232]\ vssd vssd vccd vccd la_oenb_core[30] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[31]  _253_ \mprj_logic1[233]\ vssd vssd vccd vccd la_oenb_core[31] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[32]  _254_ \mprj_logic1[234]\ vssd vssd vccd vccd la_oenb_core[32] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[33]  _255_ \mprj_logic1[235]\ vssd vssd vccd vccd la_oenb_core[33] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[34]  _256_ \mprj_logic1[236]\ vssd vssd vccd vccd la_oenb_core[34] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[35]  _257_ \mprj_logic1[237]\ vssd vssd vccd vccd la_oenb_core[35] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[36]  _258_ \mprj_logic1[238]\ vssd vssd vccd vccd la_oenb_core[36] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[37]  _259_ \mprj_logic1[239]\ vssd vssd vccd vccd la_oenb_core[37] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[38]  _260_ \mprj_logic1[240]\ vssd vssd vccd vccd la_oenb_core[38] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[39]  _261_ \mprj_logic1[241]\ vssd vssd vccd vccd la_oenb_core[39] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[3]  _262_ \mprj_logic1[205]\ vssd vssd vccd vccd la_oenb_core[3] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[40]  _263_ \mprj_logic1[242]\ vssd vssd vccd vccd la_oenb_core[40] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[41]  _264_ \mprj_logic1[243]\ vssd vssd vccd vccd la_oenb_core[41] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[42]  _265_ \mprj_logic1[244]\ vssd vssd vccd vccd la_oenb_core[42] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[43]  _266_ \mprj_logic1[245]\ vssd vssd vccd vccd la_oenb_core[43] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[44]  _267_ \mprj_logic1[246]\ vssd vssd vccd vccd la_oenb_core[44] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[45]  _268_ \mprj_logic1[247]\ vssd vssd vccd vccd la_oenb_core[45] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[46]  _269_ \mprj_logic1[248]\ vssd vssd vccd vccd la_oenb_core[46] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[47]  _270_ \mprj_logic1[249]\ vssd vssd vccd vccd la_oenb_core[47] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[48]  _271_ \mprj_logic1[250]\ vssd vssd vccd vccd la_oenb_core[48] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[49]  _272_ \mprj_logic1[251]\ vssd vssd vccd vccd la_oenb_core[49] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[4]  _273_ \mprj_logic1[206]\ vssd vssd vccd vccd la_oenb_core[4] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[50]  _274_ \mprj_logic1[252]\ vssd vssd vccd vccd la_oenb_core[50] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[51]  _275_ \mprj_logic1[253]\ vssd vssd vccd vccd la_oenb_core[51] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[52]  _276_ \mprj_logic1[254]\ vssd vssd vccd vccd la_oenb_core[52] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[53]  _277_ \mprj_logic1[255]\ vssd vssd vccd vccd la_oenb_core[53] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[54]  _278_ \mprj_logic1[256]\ vssd vssd vccd vccd la_oenb_core[54] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[55]  _279_ \mprj_logic1[257]\ vssd vssd vccd vccd la_oenb_core[55] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[56]  _280_ \mprj_logic1[258]\ vssd vssd vccd vccd la_oenb_core[56] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[57]  _281_ \mprj_logic1[259]\ vssd vssd vccd vccd la_oenb_core[57] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[58]  _282_ \mprj_logic1[260]\ vssd vssd vccd vccd la_oenb_core[58] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[59]  _283_ \mprj_logic1[261]\ vssd vssd vccd vccd la_oenb_core[59] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[5]  _284_ \mprj_logic1[207]\ vssd vssd vccd vccd la_oenb_core[5] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[60]  _285_ \mprj_logic1[262]\ vssd vssd vccd vccd la_oenb_core[60] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[61]  _286_ \mprj_logic1[263]\ vssd vssd vccd vccd la_oenb_core[61] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[62]  _287_ \mprj_logic1[264]\ vssd vssd vccd vccd la_oenb_core[62] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[63]  _288_ \mprj_logic1[265]\ vssd vssd vccd vccd la_oenb_core[63] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[64]  _289_ \mprj_logic1[266]\ vssd vssd vccd vccd la_oenb_core[64] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[65]  _290_ \mprj_logic1[267]\ vssd vssd vccd vccd la_oenb_core[65] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[66]  _291_ \mprj_logic1[268]\ vssd vssd vccd vccd la_oenb_core[66] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[67]  _292_ \mprj_logic1[269]\ vssd vssd vccd vccd la_oenb_core[67] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[68]  _293_ \mprj_logic1[270]\ vssd vssd vccd vccd la_oenb_core[68] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[69]  _294_ \mprj_logic1[271]\ vssd vssd vccd vccd la_oenb_core[69] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[6]  _295_ \mprj_logic1[208]\ vssd vssd vccd vccd la_oenb_core[6] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[70]  _296_ \mprj_logic1[272]\ vssd vssd vccd vccd la_oenb_core[70] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[71]  _297_ \mprj_logic1[273]\ vssd vssd vccd vccd la_oenb_core[71] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[72]  _298_ \mprj_logic1[274]\ vssd vssd vccd vccd la_oenb_core[72] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[73]  _299_ \mprj_logic1[275]\ vssd vssd vccd vccd la_oenb_core[73] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[74]  _300_ \mprj_logic1[276]\ vssd vssd vccd vccd la_oenb_core[74] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[75]  _301_ \mprj_logic1[277]\ vssd vssd vccd vccd la_oenb_core[75] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[76]  _302_ \mprj_logic1[278]\ vssd vssd vccd vccd la_oenb_core[76] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[77]  _303_ \mprj_logic1[279]\ vssd vssd vccd vccd la_oenb_core[77] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[78]  _304_ \mprj_logic1[280]\ vssd vssd vccd vccd la_oenb_core[78] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[79]  _305_ \mprj_logic1[281]\ vssd vssd vccd vccd la_oenb_core[79] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[7]  _306_ \mprj_logic1[209]\ vssd vssd vccd vccd la_oenb_core[7] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[80]  _307_ \mprj_logic1[282]\ vssd vssd vccd vccd la_oenb_core[80] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[81]  _308_ \mprj_logic1[283]\ vssd vssd vccd vccd la_oenb_core[81] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[82]  _309_ \mprj_logic1[284]\ vssd vssd vccd vccd la_oenb_core[82] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[83]  _310_ \mprj_logic1[285]\ vssd vssd vccd vccd la_oenb_core[83] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[84]  _311_ \mprj_logic1[286]\ vssd vssd vccd vccd la_oenb_core[84] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[85]  _312_ \mprj_logic1[287]\ vssd vssd vccd vccd la_oenb_core[85] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[86]  _313_ \mprj_logic1[288]\ vssd vssd vccd vccd la_oenb_core[86] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[87]  _314_ \mprj_logic1[289]\ vssd vssd vccd vccd la_oenb_core[87] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[88]  _315_ \mprj_logic1[290]\ vssd vssd vccd vccd la_oenb_core[88] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[89]  _316_ \mprj_logic1[291]\ vssd vssd vccd vccd la_oenb_core[89] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[8]  _317_ \mprj_logic1[210]\ vssd vssd vccd vccd la_oenb_core[8] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[90]  _318_ \mprj_logic1[292]\ vssd vssd vccd vccd la_oenb_core[90] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[91]  _319_ \mprj_logic1[293]\ vssd vssd vccd vccd la_oenb_core[91] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[92]  _320_ \mprj_logic1[294]\ vssd vssd vccd vccd la_oenb_core[92] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[93]  _321_ \mprj_logic1[295]\ vssd vssd vccd vccd la_oenb_core[93] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[94]  _322_ \mprj_logic1[296]\ vssd vssd vccd vccd la_oenb_core[94] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[95]  _323_ \mprj_logic1[297]\ vssd vssd vccd vccd la_oenb_core[95] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[96]  _324_ \mprj_logic1[298]\ vssd vssd vccd vccd la_oenb_core[96] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[97]  _325_ \mprj_logic1[299]\ vssd vssd vccd vccd la_oenb_core[97] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[98]  _326_ \mprj_logic1[300]\ vssd vssd vccd vccd la_oenb_core[98] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[99]  _327_ \mprj_logic1[301]\ vssd vssd vccd vccd la_oenb_core[99] sky130_fd_sc_hd__einvp_8
X\user_to_mprj_oen_buffers[9]  _328_ \mprj_logic1[211]\ vssd vssd vccd vccd la_oenb_core[9] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_wb_ena_buf net614 \mprj_logic1[462]\ vssd vssd vccd vccd wb_in_enable sky130_fd_sc_hd__and2_4
Xuser_wb_ack_buffer mprj_ack_i_core_bar vssd vssd vccd vccd net755 sky130_fd_sc_hd__clkinv_8
Xuser_wb_ack_gate net516 wb_in_enable vssd vssd vccd vccd mprj_ack_i_core_bar sky130_fd_sc_hd__nand2_4
X\user_wb_dat_buffers[0]  \mprj_dat_i_core_bar[0]\ vssd vssd vccd vccd net756 sky130_fd_sc_hd__clkinv_8
X\user_wb_dat_buffers[10]  \mprj_dat_i_core_bar[10]\ vssd vssd vccd vccd net757 sky130_fd_sc_hd__clkinv_8
X\user_wb_dat_buffers[11]  \mprj_dat_i_core_bar[11]\ vssd vssd vccd vccd net758 sky130_fd_sc_hd__clkinv_8
X\user_wb_dat_buffers[12]  \mprj_dat_i_core_bar[12]\ vssd vssd vccd vccd net759 sky130_fd_sc_hd__clkinv_8
X\user_wb_dat_buffers[13]  \mprj_dat_i_core_bar[13]\ vssd vssd vccd vccd net760 sky130_fd_sc_hd__clkinv_8
X\user_wb_dat_buffers[14]  \mprj_dat_i_core_bar[14]\ vssd vssd vccd vccd net761 sky130_fd_sc_hd__clkinv_8
X\user_wb_dat_buffers[15]  \mprj_dat_i_core_bar[15]\ vssd vssd vccd vccd net762 sky130_fd_sc_hd__clkinv_4
X\user_wb_dat_buffers[16]  \mprj_dat_i_core_bar[16]\ vssd vssd vccd vccd net763 sky130_fd_sc_hd__clkinv_4
X\user_wb_dat_buffers[17]  \mprj_dat_i_core_bar[17]\ vssd vssd vccd vccd net764 sky130_fd_sc_hd__clkinv_4
X\user_wb_dat_buffers[18]  \mprj_dat_i_core_bar[18]\ vssd vssd vccd vccd net765 sky130_fd_sc_hd__inv_6
X\user_wb_dat_buffers[19]  \mprj_dat_i_core_bar[19]\ vssd vssd vccd vccd net766 sky130_fd_sc_hd__clkinv_8
X\user_wb_dat_buffers[1]  \mprj_dat_i_core_bar[1]\ vssd vssd vccd vccd net767 sky130_fd_sc_hd__clkinv_8
X\user_wb_dat_buffers[20]  \mprj_dat_i_core_bar[20]\ vssd vssd vccd vccd net768 sky130_fd_sc_hd__clkinv_8
X\user_wb_dat_buffers[21]  \mprj_dat_i_core_bar[21]\ vssd vssd vccd vccd net769 sky130_fd_sc_hd__clkinv_8
X\user_wb_dat_buffers[22]  \mprj_dat_i_core_bar[22]\ vssd vssd vccd vccd net770 sky130_fd_sc_hd__clkinv_8
X\user_wb_dat_buffers[23]  \mprj_dat_i_core_bar[23]\ vssd vssd vccd vccd net771 sky130_fd_sc_hd__inv_6
X\user_wb_dat_buffers[24]  \mprj_dat_i_core_bar[24]\ vssd vssd vccd vccd net772 sky130_fd_sc_hd__clkinv_8
X\user_wb_dat_buffers[25]  \mprj_dat_i_core_bar[25]\ vssd vssd vccd vccd net773 sky130_fd_sc_hd__inv_6
X\user_wb_dat_buffers[26]  \mprj_dat_i_core_bar[26]\ vssd vssd vccd vccd net774 sky130_fd_sc_hd__clkinv_8
X\user_wb_dat_buffers[27]  \mprj_dat_i_core_bar[27]\ vssd vssd vccd vccd net775 sky130_fd_sc_hd__clkinv_8
X\user_wb_dat_buffers[28]  \mprj_dat_i_core_bar[28]\ vssd vssd vccd vccd net776 sky130_fd_sc_hd__clkinv_8
X\user_wb_dat_buffers[29]  \mprj_dat_i_core_bar[29]\ vssd vssd vccd vccd net777 sky130_fd_sc_hd__clkinv_8
X\user_wb_dat_buffers[2]  \mprj_dat_i_core_bar[2]\ vssd vssd vccd vccd net778 sky130_fd_sc_hd__clkinv_8
X\user_wb_dat_buffers[30]  \mprj_dat_i_core_bar[30]\ vssd vssd vccd vccd net779 sky130_fd_sc_hd__clkinv_8
X\user_wb_dat_buffers[31]  \mprj_dat_i_core_bar[31]\ vssd vssd vccd vccd net780 sky130_fd_sc_hd__inv_6
X\user_wb_dat_buffers[3]  \mprj_dat_i_core_bar[3]\ vssd vssd vccd vccd net781 sky130_fd_sc_hd__clkinv_8
X\user_wb_dat_buffers[4]  \mprj_dat_i_core_bar[4]\ vssd vssd vccd vccd net782 sky130_fd_sc_hd__clkinv_8
X\user_wb_dat_buffers[5]  \mprj_dat_i_core_bar[5]\ vssd vssd vccd vccd net783 sky130_fd_sc_hd__clkinv_8
X\user_wb_dat_buffers[6]  \mprj_dat_i_core_bar[6]\ vssd vssd vccd vccd net784 sky130_fd_sc_hd__clkinv_8
X\user_wb_dat_buffers[7]  \mprj_dat_i_core_bar[7]\ vssd vssd vccd vccd net785 sky130_fd_sc_hd__clkinv_8
X\user_wb_dat_buffers[8]  \mprj_dat_i_core_bar[8]\ vssd vssd vccd vccd net786 sky130_fd_sc_hd__clkinv_8
X\user_wb_dat_buffers[9]  \mprj_dat_i_core_bar[9]\ vssd vssd vccd vccd net787 sky130_fd_sc_hd__clkinv_8
X\user_wb_dat_gates[0]  net550 wb_in_enable vssd vssd vccd vccd \mprj_dat_i_core_bar[0]\ sky130_fd_sc_hd__nand2_4
X\user_wb_dat_gates[10]  net551 wb_in_enable vssd vssd vccd vccd \mprj_dat_i_core_bar[10]\ sky130_fd_sc_hd__nand2_4
X\user_wb_dat_gates[11]  net552 wb_in_enable vssd vssd vccd vccd \mprj_dat_i_core_bar[11]\ sky130_fd_sc_hd__nand2_4
X\user_wb_dat_gates[12]  net553 wb_in_enable vssd vssd vccd vccd \mprj_dat_i_core_bar[12]\ sky130_fd_sc_hd__nand2_4
X\user_wb_dat_gates[13]  net554 wb_in_enable vssd vssd vccd vccd \mprj_dat_i_core_bar[13]\ sky130_fd_sc_hd__nand2_4
X\user_wb_dat_gates[14]  net555 wb_in_enable vssd vssd vccd vccd \mprj_dat_i_core_bar[14]\ sky130_fd_sc_hd__nand2_4
X\user_wb_dat_gates[15]  net556 wb_in_enable vssd vssd vccd vccd \mprj_dat_i_core_bar[15]\ sky130_fd_sc_hd__nand2_4
X\user_wb_dat_gates[16]  net557 wb_in_enable vssd vssd vccd vccd \mprj_dat_i_core_bar[16]\ sky130_fd_sc_hd__nand2_8
X\user_wb_dat_gates[17]  net558 wb_in_enable vssd vssd vccd vccd \mprj_dat_i_core_bar[17]\ sky130_fd_sc_hd__nand2_4
X\user_wb_dat_gates[18]  net559 wb_in_enable vssd vssd vccd vccd \mprj_dat_i_core_bar[18]\ sky130_fd_sc_hd__nand2_4
X\user_wb_dat_gates[19]  net560 wb_in_enable vssd vssd vccd vccd \mprj_dat_i_core_bar[19]\ sky130_fd_sc_hd__nand2_4
X\user_wb_dat_gates[1]  net561 wb_in_enable vssd vssd vccd vccd \mprj_dat_i_core_bar[1]\ sky130_fd_sc_hd__nand2_8
X\user_wb_dat_gates[20]  net562 wb_in_enable vssd vssd vccd vccd \mprj_dat_i_core_bar[20]\ sky130_fd_sc_hd__nand2_4
X\user_wb_dat_gates[21]  net563 wb_in_enable vssd vssd vccd vccd \mprj_dat_i_core_bar[21]\ sky130_fd_sc_hd__nand2_2
X\user_wb_dat_gates[22]  net564 wb_in_enable vssd vssd vccd vccd \mprj_dat_i_core_bar[22]\ sky130_fd_sc_hd__nand2_2
X\user_wb_dat_gates[23]  net565 wb_in_enable vssd vssd vccd vccd \mprj_dat_i_core_bar[23]\ sky130_fd_sc_hd__nand2_2
X\user_wb_dat_gates[24]  net566 wb_in_enable vssd vssd vccd vccd \mprj_dat_i_core_bar[24]\ sky130_fd_sc_hd__nand2_2
X\user_wb_dat_gates[25]  net567 wb_in_enable vssd vssd vccd vccd \mprj_dat_i_core_bar[25]\ sky130_fd_sc_hd__nand2_2
X\user_wb_dat_gates[26]  net568 wb_in_enable vssd vssd vccd vccd \mprj_dat_i_core_bar[26]\ sky130_fd_sc_hd__nand2_4
X\user_wb_dat_gates[27]  net569 wb_in_enable vssd vssd vccd vccd \mprj_dat_i_core_bar[27]\ sky130_fd_sc_hd__nand2_2
X\user_wb_dat_gates[28]  net570 wb_in_enable vssd vssd vccd vccd \mprj_dat_i_core_bar[28]\ sky130_fd_sc_hd__nand2_2
X\user_wb_dat_gates[29]  net571 wb_in_enable vssd vssd vccd vccd \mprj_dat_i_core_bar[29]\ sky130_fd_sc_hd__nand2_2
X\user_wb_dat_gates[2]  net572 wb_in_enable vssd vssd vccd vccd \mprj_dat_i_core_bar[2]\ sky130_fd_sc_hd__nand2_8
X\user_wb_dat_gates[30]  net573 wb_in_enable vssd vssd vccd vccd \mprj_dat_i_core_bar[30]\ sky130_fd_sc_hd__nand2_2
X\user_wb_dat_gates[31]  net574 wb_in_enable vssd vssd vccd vccd \mprj_dat_i_core_bar[31]\ sky130_fd_sc_hd__nand2_2
X\user_wb_dat_gates[3]  net575 wb_in_enable vssd vssd vccd vccd \mprj_dat_i_core_bar[3]\ sky130_fd_sc_hd__nand2_4
X\user_wb_dat_gates[4]  net576 wb_in_enable vssd vssd vccd vccd \mprj_dat_i_core_bar[4]\ sky130_fd_sc_hd__nand2_4
X\user_wb_dat_gates[5]  net577 wb_in_enable vssd vssd vccd vccd \mprj_dat_i_core_bar[5]\ sky130_fd_sc_hd__nand2_4
X\user_wb_dat_gates[6]  net578 wb_in_enable vssd vssd vccd vccd \mprj_dat_i_core_bar[6]\ sky130_fd_sc_hd__nand2_4
X\user_wb_dat_gates[7]  net579 wb_in_enable vssd vssd vccd vccd \mprj_dat_i_core_bar[7]\ sky130_fd_sc_hd__nand2_8
X\user_wb_dat_gates[8]  net580 wb_in_enable vssd vssd vccd vccd \mprj_dat_i_core_bar[8]\ sky130_fd_sc_hd__nand2_4
X\user_wb_dat_gates[9]  net581 wb_in_enable vssd vssd vccd vccd \mprj_dat_i_core_bar[9]\ sky130_fd_sc_hd__nand2_4

.ends
.end
