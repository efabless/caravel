VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mprj_vias
  CLASS BLOCK ;
  FOREIGN mprj_vias ;
  ORIGIN 0.000 0.000 ;
  SIZE 0 BY 0 ;
END mprj_vias
END LIBRARY

