* NGSPICE file created from housekeeping.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtn_1 abstract view
.subckt sky130_fd_sc_hd__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_1 abstract view
.subckt sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_1 abstract view
.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

.subckt housekeeping VGND VPWR debug_in debug_mode debug_oeb debug_out irq[0] irq[1]
+ irq[2] mask_rev_in[0] mask_rev_in[10] mask_rev_in[11] mask_rev_in[12] mask_rev_in[13]
+ mask_rev_in[14] mask_rev_in[15] mask_rev_in[16] mask_rev_in[17] mask_rev_in[18]
+ mask_rev_in[19] mask_rev_in[1] mask_rev_in[20] mask_rev_in[21] mask_rev_in[22] mask_rev_in[23]
+ mask_rev_in[24] mask_rev_in[25] mask_rev_in[26] mask_rev_in[27] mask_rev_in[28]
+ mask_rev_in[29] mask_rev_in[2] mask_rev_in[30] mask_rev_in[31] mask_rev_in[3] mask_rev_in[4]
+ mask_rev_in[5] mask_rev_in[6] mask_rev_in[7] mask_rev_in[8] mask_rev_in[9] mgmt_gpio_in[0]
+ mgmt_gpio_in[10] mgmt_gpio_in[11] mgmt_gpio_in[12] mgmt_gpio_in[13] mgmt_gpio_in[14]
+ mgmt_gpio_in[15] mgmt_gpio_in[16] mgmt_gpio_in[17] mgmt_gpio_in[18] mgmt_gpio_in[19]
+ mgmt_gpio_in[1] mgmt_gpio_in[20] mgmt_gpio_in[21] mgmt_gpio_in[22] mgmt_gpio_in[23]
+ mgmt_gpio_in[24] mgmt_gpio_in[25] mgmt_gpio_in[26] mgmt_gpio_in[27] mgmt_gpio_in[28]
+ mgmt_gpio_in[29] mgmt_gpio_in[2] mgmt_gpio_in[30] mgmt_gpio_in[31] mgmt_gpio_in[32]
+ mgmt_gpio_in[33] mgmt_gpio_in[34] mgmt_gpio_in[35] mgmt_gpio_in[36] mgmt_gpio_in[37]
+ mgmt_gpio_in[3] mgmt_gpio_in[4] mgmt_gpio_in[5] mgmt_gpio_in[6] mgmt_gpio_in[7]
+ mgmt_gpio_in[8] mgmt_gpio_in[9] mgmt_gpio_oeb[0] mgmt_gpio_oeb[10] mgmt_gpio_oeb[11]
+ mgmt_gpio_oeb[12] mgmt_gpio_oeb[13] mgmt_gpio_oeb[14] mgmt_gpio_oeb[15] mgmt_gpio_oeb[16]
+ mgmt_gpio_oeb[17] mgmt_gpio_oeb[18] mgmt_gpio_oeb[19] mgmt_gpio_oeb[1] mgmt_gpio_oeb[20]
+ mgmt_gpio_oeb[21] mgmt_gpio_oeb[22] mgmt_gpio_oeb[23] mgmt_gpio_oeb[24] mgmt_gpio_oeb[25]
+ mgmt_gpio_oeb[26] mgmt_gpio_oeb[27] mgmt_gpio_oeb[28] mgmt_gpio_oeb[29] mgmt_gpio_oeb[2]
+ mgmt_gpio_oeb[30] mgmt_gpio_oeb[31] mgmt_gpio_oeb[32] mgmt_gpio_oeb[33] mgmt_gpio_oeb[34]
+ mgmt_gpio_oeb[35] mgmt_gpio_oeb[36] mgmt_gpio_oeb[37] mgmt_gpio_oeb[3] mgmt_gpio_oeb[4]
+ mgmt_gpio_oeb[5] mgmt_gpio_oeb[6] mgmt_gpio_oeb[7] mgmt_gpio_oeb[8] mgmt_gpio_oeb[9]
+ mgmt_gpio_out[0] mgmt_gpio_out[10] mgmt_gpio_out[11] mgmt_gpio_out[12] mgmt_gpio_out[13]
+ mgmt_gpio_out[14] mgmt_gpio_out[15] mgmt_gpio_out[16] mgmt_gpio_out[17] mgmt_gpio_out[18]
+ mgmt_gpio_out[19] mgmt_gpio_out[1] mgmt_gpio_out[20] mgmt_gpio_out[21] mgmt_gpio_out[22]
+ mgmt_gpio_out[23] mgmt_gpio_out[24] mgmt_gpio_out[25] mgmt_gpio_out[26] mgmt_gpio_out[27]
+ mgmt_gpio_out[28] mgmt_gpio_out[29] mgmt_gpio_out[2] mgmt_gpio_out[30] mgmt_gpio_out[31]
+ mgmt_gpio_out[32] mgmt_gpio_out[33] mgmt_gpio_out[34] mgmt_gpio_out[35] mgmt_gpio_out[36]
+ mgmt_gpio_out[37] mgmt_gpio_out[3] mgmt_gpio_out[4] mgmt_gpio_out[5] mgmt_gpio_out[6]
+ mgmt_gpio_out[7] mgmt_gpio_out[8] mgmt_gpio_out[9] pad_flash_clk pad_flash_clk_oeb
+ pad_flash_csb pad_flash_csb_oeb pad_flash_io0_di pad_flash_io0_do pad_flash_io0_ieb
+ pad_flash_io0_oeb pad_flash_io1_di pad_flash_io1_do pad_flash_io1_ieb pad_flash_io1_oeb
+ pll90_sel[0] pll90_sel[1] pll90_sel[2] pll_bypass pll_dco_ena pll_div[0] pll_div[1]
+ pll_div[2] pll_div[3] pll_div[4] pll_ena pll_sel[0] pll_sel[1] pll_sel[2] pll_trim[0]
+ pll_trim[10] pll_trim[11] pll_trim[12] pll_trim[13] pll_trim[14] pll_trim[15] pll_trim[16]
+ pll_trim[17] pll_trim[18] pll_trim[19] pll_trim[1] pll_trim[20] pll_trim[21] pll_trim[22]
+ pll_trim[23] pll_trim[24] pll_trim[25] pll_trim[2] pll_trim[3] pll_trim[4] pll_trim[5]
+ pll_trim[6] pll_trim[7] pll_trim[8] pll_trim[9] porb pwr_ctrl_out[0] pwr_ctrl_out[1]
+ pwr_ctrl_out[2] pwr_ctrl_out[3] qspi_enabled reset ser_rx ser_tx serial_clock serial_data_1
+ serial_data_2 serial_load serial_resetn spi_csb spi_enabled spi_sck spi_sdi spi_sdo
+ spi_sdoenb spimemio_flash_clk spimemio_flash_csb spimemio_flash_io0_di spimemio_flash_io0_do
+ spimemio_flash_io0_oeb spimemio_flash_io1_di spimemio_flash_io1_do spimemio_flash_io1_oeb
+ spimemio_flash_io2_di spimemio_flash_io2_do spimemio_flash_io2_oeb spimemio_flash_io3_di
+ spimemio_flash_io3_do spimemio_flash_io3_oeb trap uart_enabled user_clock usr1_vcc_pwrgood
+ usr1_vdd_pwrgood usr2_vcc_pwrgood usr2_vdd_pwrgood wb_ack_o wb_adr_i[0] wb_adr_i[10]
+ wb_adr_i[11] wb_adr_i[12] wb_adr_i[13] wb_adr_i[14] wb_adr_i[15] wb_adr_i[16] wb_adr_i[17]
+ wb_adr_i[18] wb_adr_i[19] wb_adr_i[1] wb_adr_i[20] wb_adr_i[21] wb_adr_i[22] wb_adr_i[23]
+ wb_adr_i[24] wb_adr_i[25] wb_adr_i[26] wb_adr_i[27] wb_adr_i[28] wb_adr_i[29] wb_adr_i[2]
+ wb_adr_i[30] wb_adr_i[31] wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6] wb_adr_i[7]
+ wb_adr_i[8] wb_adr_i[9] wb_clk_i wb_cyc_i wb_dat_i[0] wb_dat_i[10] wb_dat_i[11]
+ wb_dat_i[12] wb_dat_i[13] wb_dat_i[14] wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18]
+ wb_dat_i[19] wb_dat_i[1] wb_dat_i[20] wb_dat_i[21] wb_dat_i[22] wb_dat_i[23] wb_dat_i[24]
+ wb_dat_i[25] wb_dat_i[26] wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[2] wb_dat_i[30]
+ wb_dat_i[31] wb_dat_i[3] wb_dat_i[4] wb_dat_i[5] wb_dat_i[6] wb_dat_i[7] wb_dat_i[8]
+ wb_dat_i[9] wb_dat_o[0] wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13] wb_dat_o[14]
+ wb_dat_o[15] wb_dat_o[16] wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[1] wb_dat_o[20]
+ wb_dat_o[21] wb_dat_o[22] wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26] wb_dat_o[27]
+ wb_dat_o[28] wb_dat_o[29] wb_dat_o[2] wb_dat_o[30] wb_dat_o[31] wb_dat_o[3] wb_dat_o[4]
+ wb_dat_o[5] wb_dat_o[6] wb_dat_o[7] wb_dat_o[8] wb_dat_o[9] wb_rstn_i wb_sel_i[0]
+ wb_sel_i[1] wb_sel_i[2] wb_sel_i[3] wb_stb_i wb_we_i
XFILLER_39_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6914_ _7123_/CLK _6914_/D _6407_/A VGND VGND VPWR VPWR _6914_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6845_ _7068_/CLK _6845_/D fanout505/X VGND VGND VPWR VPWR _6845_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6776_ _7200_/CLK _6776_/D _6348_/B VGND VGND VPWR VPWR _6776_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_168_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3988_ hold486/X _6397_/A0 _3991_/S VGND VGND VPWR VPWR _3988_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5727_ _7019_/Q _5663_/X _5678_/X _7067_/Q _5726_/X VGND VGND VPWR VPWR _5728_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_109_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5658_ _7151_/Q _7150_/Q VGND VGND VPWR VPWR _5706_/C sky130_fd_sc_hd__and2_2
X_4609_ _5036_/A _4609_/B _4794_/A VGND VGND VPWR VPWR _5095_/A sky130_fd_sc_hd__nor3_2
XFILLER_190_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5589_ _6562_/Q _5648_/C _7143_/Q VGND VGND VPWR VPWR _5589_/X sky130_fd_sc_hd__a21o_1
XFILLER_151_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold340 _5324_/X VGND VGND VPWR VPWR _6907_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold351 _6883_/Q VGND VGND VPWR VPWR hold351/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold362 _4179_/X VGND VGND VPWR VPWR _6638_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 _7112_/Q VGND VGND VPWR VPWR hold373/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 _4256_/X VGND VGND VPWR VPWR _6709_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold395 _7073_/Q VGND VGND VPWR VPWR hold395/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1040 _4074_/X VGND VGND VPWR VPWR _6555_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1051 _6898_/Q VGND VGND VPWR VPWR _5314_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1062 _4277_/X VGND VGND VPWR VPWR _6726_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1073 _6930_/Q VGND VGND VPWR VPWR _5350_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1084 _5269_/X VGND VGND VPWR VPWR _6858_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_202 _5681_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1095 _5581_/X VGND VGND VPWR VPWR _7135_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_213 _7169_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_224 _5376_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_235 _5555_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_246 _5677_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_257 _5581_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4960_ _4960_/A _4960_/B _4959_/X VGND VGND VPWR VPWR _4961_/B sky130_fd_sc_hd__or3b_1
XFILLER_17_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3911_ _6346_/A _3888_/B _3191_/Y VGND VGND VPWR VPWR _3911_/Y sky130_fd_sc_hd__o21ai_1
X_4891_ _4516_/B _4871_/Y _4880_/X _4890_/X VGND VGND VPWR VPWR _4891_/X sky130_fd_sc_hd__a211o_1
XFILLER_149_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6630_ _7193_/CLK _6630_/D VGND VGND VPWR VPWR _6630_/Q sky130_fd_sc_hd__dfxtp_1
X_3842_ _6456_/Q _3794_/B _6458_/Q VGND VGND VPWR VPWR _3842_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6561_ _7033_/CLK _6561_/D fanout504/X VGND VGND VPWR VPWR _6561_/Q sky130_fd_sc_hd__dfrtp_4
X_3773_ _7066_/Q _5502_/A _4028_/A _6521_/Q VGND VGND VPWR VPWR _3773_/X sky130_fd_sc_hd__a22o_1
XFILLER_192_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5512_ _5536_/A1 _5512_/A1 _5519_/S VGND VGND VPWR VPWR _5512_/X sky130_fd_sc_hd__mux2_1
X_6492_ _6759_/CLK _6492_/D fanout488/X VGND VGND VPWR VPWR _6492_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_172_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5443_ _5584_/A0 hold429/X _5447_/S VGND VGND VPWR VPWR _5443_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5374_ _5569_/A0 hold319/X _5375_/S VGND VGND VPWR VPWR _5374_/X sky130_fd_sc_hd__mux2_1
X_7113_ _7135_/CLK _7113_/D fanout519/X VGND VGND VPWR VPWR _7113_/Q sky130_fd_sc_hd__dfrtp_1
X_4325_ _4325_/A0 _5212_/C _4329_/S VGND VGND VPWR VPWR _4325_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7044_ _7137_/CLK _7044_/D fanout501/X VGND VGND VPWR VPWR _7044_/Q sky130_fd_sc_hd__dfrtp_4
X_4256_ hold383/X _5533_/A1 _4257_/S VGND VGND VPWR VPWR _4256_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3207_ _7061_/Q VGND VGND VPWR VPWR _3207_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4187_ _4187_/A0 _3410_/X _4188_/S VGND VGND VPWR VPWR _6645_/D sky130_fd_sc_hd__mux2_1
XFILLER_27_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6828_ _7138_/CLK _6828_/D fanout520/X VGND VGND VPWR VPWR _6828_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6759_ _6759_/CLK _6759_/D fanout489/X VGND VGND VPWR VPWR _6759_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_109_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold170 _4157_/X VGND VGND VPWR VPWR _6619_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold181 _6624_/Q VGND VGND VPWR VPWR hold181/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 _5215_/X VGND VGND VPWR VPWR _6813_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_120_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4110_ hold127/X hold173/X _4110_/S VGND VGND VPWR VPWR _4110_/X sky130_fd_sc_hd__mux2_1
X_5090_ _5090_/A _5090_/B _5089_/X VGND VGND VPWR VPWR _5170_/B sky130_fd_sc_hd__or3b_1
X_4041_ _5476_/A0 _4041_/A1 _4045_/S VGND VGND VPWR VPWR _4041_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5992_ _6033_/A _6020_/C _6040_/C VGND VGND VPWR VPWR _5992_/X sky130_fd_sc_hd__and3_4
XFILLER_24_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4943_ _4395_/Y _5060_/B _4833_/Y VGND VGND VPWR VPWR _5053_/B sky130_fd_sc_hd__a21o_1
XFILLER_17_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4874_ _5001_/A _4931_/B _5001_/C VGND VGND VPWR VPWR _4897_/C sky130_fd_sc_hd__and3_1
XFILLER_177_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6613_ _6708_/CLK _6613_/D _6432_/A VGND VGND VPWR VPWR _6613_/Q sky130_fd_sc_hd__dfrtp_4
X_3825_ _3824_/X _3825_/A1 _3833_/S VGND VGND VPWR VPWR _6466_/D sky130_fd_sc_hd__mux2_1
XFILLER_193_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6544_ _3945_/A1 _6544_/D _6432_/X VGND VGND VPWR VPWR hold72/A sky130_fd_sc_hd__dfrtp_4
XFILLER_158_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3756_ _7103_/Q _5544_/A _4104_/A input61/X _3739_/X VGND VGND VPWR VPWR _3760_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_5_0_csclk clkbuf_3_5_0_csclk/A VGND VGND VPWR VPWR _6882_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_145_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6475_ _6760_/CLK _6475_/D fanout490/X VGND VGND VPWR VPWR _6475_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_145_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3687_ _6995_/Q _3300_/Y _4022_/A _6517_/Q _3686_/X VGND VGND VPWR VPWR _3688_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_106_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5426_ _5558_/A0 hold187/X _5429_/S VGND VGND VPWR VPWR _5426_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput220 _6546_/Q VGND VGND VPWR VPWR mgmt_gpio_out[16] sky130_fd_sc_hd__buf_12
Xoutput231 _6828_/Q VGND VGND VPWR VPWR mgmt_gpio_out[26] sky130_fd_sc_hd__buf_12
Xoutput242 _3919_/X VGND VGND VPWR VPWR mgmt_gpio_out[36] sky130_fd_sc_hd__buf_12
Xoutput253 _3943_/X VGND VGND VPWR VPWR pad_flash_csb sky130_fd_sc_hd__buf_12
XFILLER_133_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput264 _6806_/Q VGND VGND VPWR VPWR pll_bypass sky130_fd_sc_hd__buf_12
X_5357_ _5552_/A0 hold504/X _5357_/S VGND VGND VPWR VPWR _5357_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput275 _6490_/Q VGND VGND VPWR VPWR pll_trim[0] sky130_fd_sc_hd__buf_12
XFILLER_87_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput286 _6491_/Q VGND VGND VPWR VPWR pll_trim[1] sky130_fd_sc_hd__buf_12
Xoutput297 _6496_/Q VGND VGND VPWR VPWR pll_trim[6] sky130_fd_sc_hd__buf_12
X_4308_ _5531_/A1 hold948/X _4311_/S VGND VGND VPWR VPWR _4308_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5288_ hold9/X _5288_/A1 hold32/X VGND VGND VPWR VPWR hold33/A sky130_fd_sc_hd__mux2_1
XFILLER_59_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7027_ _7078_/CLK _7027_/D fanout515/X VGND VGND VPWR VPWR _7027_/Q sky130_fd_sc_hd__dfstp_1
X_4239_ _5549_/A0 hold377/X hold59/X VGND VGND VPWR VPWR _4239_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout491 fanout527/X VGND VGND VPWR VPWR fanout491/X sky130_fd_sc_hd__buf_6
XFILLER_171_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3610_ _6618_/Q _4153_/A _4141_/A _6608_/Q VGND VGND VPWR VPWR _3610_/X sky130_fd_sc_hd__a22o_1
XFILLER_159_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4590_ _5076_/B _4694_/B VGND VGND VPWR VPWR _4598_/B sky130_fd_sc_hd__nor2_1
X_3541_ _3541_/A _3541_/B _3541_/C _3541_/D VGND VGND VPWR VPWR _3542_/D sky130_fd_sc_hd__or4_1
XFILLER_190_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold906 hold906/A VGND VGND VPWR VPWR hold906/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold917 _3980_/X VGND VGND VPWR VPWR _6480_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold928 _6851_/Q VGND VGND VPWR VPWR hold928/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold939 _5437_/X VGND VGND VPWR VPWR _7008_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6260_ _6666_/Q wire412/X _6016_/X hold89/A VGND VGND VPWR VPWR _6260_/X sky130_fd_sc_hd__a22o_1
X_3472_ _3731_/A _3538_/B VGND VGND VPWR VPWR _3472_/Y sky130_fd_sc_hd__nor2_1
X_5211_ _6393_/A0 _5211_/A1 _5211_/S VGND VGND VPWR VPWR _5211_/X sky130_fd_sc_hd__mux2_1
X_6191_ _7080_/Q _5994_/X _6030_/X _7000_/Q _6190_/X VGND VGND VPWR VPWR _6192_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_170_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5142_ _5142_/A _5142_/B _5141_/X VGND VGND VPWR VPWR _5172_/C sky130_fd_sc_hd__or3b_1
XFILLER_111_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1606 _6691_/Q VGND VGND VPWR VPWR _3888_/A sky130_fd_sc_hd__dlygate4sd3_1
X_5073_ _5095_/A _5073_/B _5072_/X VGND VGND VPWR VPWR _5155_/B sky130_fd_sc_hd__or3b_1
X_4024_ _4024_/A0 _6394_/A0 _4027_/S VGND VGND VPWR VPWR _4024_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5975_ _7157_/Q _7158_/Q VGND VGND VPWR VPWR _6021_/A sky130_fd_sc_hd__or2_4
X_4926_ _4926_/A _4992_/B VGND VGND VPWR VPWR _5031_/C sky130_fd_sc_hd__nand2_1
XFILLER_21_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4857_ _4857_/A _4857_/B _4857_/C _4857_/D VGND VGND VPWR VPWR _4857_/X sky130_fd_sc_hd__and4_1
XFILLER_165_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3808_ hold16/A _3823_/B VGND VGND VPWR VPWR _3821_/S sky130_fd_sc_hd__and2_1
XFILLER_165_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4788_ _5003_/A _4802_/A _5076_/B _4679_/B VGND VGND VPWR VPWR _4985_/C sky130_fd_sc_hd__o22ai_1
X_6527_ _7207_/CLK _6527_/D fanout484/X VGND VGND VPWR VPWR _6527_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_118_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3739_ _6890_/Q _5304_/A _5571_/A _7127_/Q VGND VGND VPWR VPWR _3739_/X sky130_fd_sc_hd__a22o_1
X_6458_ _3945_/A1 _6458_/D _6413_/X VGND VGND VPWR VPWR _6458_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_134_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5409_ _5586_/A0 _5409_/A1 _5411_/S VGND VGND VPWR VPWR _5409_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6389_ _6699_/Q _6389_/A2 _6388_/X VGND VGND VPWR VPWR _6389_/X sky130_fd_sc_hd__a21o_1
XFILLER_87_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5760_ _7069_/Q _5678_/X _5682_/X _7085_/Q _5759_/X VGND VGND VPWR VPWR _5771_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_15_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4711_ _4814_/A _5023_/B _4839_/B _4689_/X _4710_/X VGND VGND VPWR VPWR _4713_/C
+ sky130_fd_sc_hd__o311a_1
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5691_ _5960_/B _5691_/B VGND VGND VPWR VPWR _5691_/Y sky130_fd_sc_hd__nand2_8
XFILLER_147_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4642_ _4642_/A _4642_/B _4642_/C _4642_/D VGND VGND VPWR VPWR _4642_/X sky130_fd_sc_hd__and4_1
XFILLER_163_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4573_ _4484_/B _4573_/B VGND VGND VPWR VPWR _4981_/C sky130_fd_sc_hd__nand2b_2
Xmax_cap400 _6023_/B VGND VGND VPWR VPWR _6308_/A2 sky130_fd_sc_hd__buf_8
XFILLER_162_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap411 _6022_/C VGND VGND VPWR VPWR _6336_/A2 sky130_fd_sc_hd__buf_12
Xhold703 _6689_/Q VGND VGND VPWR VPWR hold703/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold714 _4323_/X VGND VGND VPWR VPWR _6765_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap422 _5661_/X VGND VGND VPWR VPWR _5846_/A2 sky130_fd_sc_hd__buf_8
X_6312_ _6689_/Q _6024_/A _6040_/X _6529_/Q VGND VGND VPWR VPWR _6312_/X sky130_fd_sc_hd__a22o_1
Xmax_cap433 _4228_/Y VGND VGND VPWR VPWR _6390_/A2 sky130_fd_sc_hd__clkbuf_2
X_3524_ _3524_/A _3524_/B _3524_/C _3524_/D VGND VGND VPWR VPWR _3542_/C sky130_fd_sc_hd__or4_2
Xhold725 _6481_/Q VGND VGND VPWR VPWR hold725/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold736 _5417_/X VGND VGND VPWR VPWR _6990_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold747 _6534_/Q VGND VGND VPWR VPWR hold747/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold758 _5519_/X VGND VGND VPWR VPWR _7081_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6243_ _6596_/Q _6046_/B _6232_/X _6242_/X _6318_/S VGND VGND VPWR VPWR _6243_/X
+ sky130_fd_sc_hd__o221a_1
Xhold769 _6902_/Q VGND VGND VPWR VPWR hold769/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_170_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3455_ hold57/X _3495_/A VGND VGND VPWR VPWR _4040_/A sky130_fd_sc_hd__nor2_4
XFILLER_115_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6174_ _6904_/Q _6022_/B _6199_/B1 _6872_/Q VGND VGND VPWR VPWR _6174_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3386_ _6952_/Q _5367_/A _5562_/A _7125_/Q _3381_/X VGND VGND VPWR VPWR _3392_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_57_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5125_ _5125_/A _5125_/B VGND VGND VPWR VPWR _5128_/C sky130_fd_sc_hd__nor2_1
Xhold1403 _6683_/Q VGND VGND VPWR VPWR _4237_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1414 _7192_/Q VGND VGND VPWR VPWR hold1414/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1425 _6642_/Q VGND VGND VPWR VPWR _4184_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1436 _7189_/Q VGND VGND VPWR VPWR _6349_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1447 _5359_/X VGND VGND VPWR VPWR _6938_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5056_ _5023_/A _4694_/B _4950_/B _4887_/C VGND VGND VPWR VPWR _5056_/X sky130_fd_sc_hd__o211a_1
Xhold1458 _6778_/Q VGND VGND VPWR VPWR _5034_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1469 _3449_/X VGND VGND VPWR VPWR _6788_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4007_ _5586_/A0 _4007_/A1 _4009_/S VGND VGND VPWR VPWR _4007_/X sky130_fd_sc_hd__mux2_1
XTAP_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_1_wb_clk_i clkbuf_1_0_1_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_2_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_80_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5958_ _6725_/Q _5702_/X _5706_/X _7094_/Q VGND VGND VPWR VPWR _5958_/X sky130_fd_sc_hd__a22o_1
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4909_ _4915_/C VGND VGND VPWR VPWR _4909_/Y sky130_fd_sc_hd__inv_2
X_5889_ _6722_/Q _5702_/X _5706_/X _7091_/Q VGND VGND VPWR VPWR _5889_/X sky130_fd_sc_hd__a22o_1
XFILLER_187_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_2_2_0_csclk clkbuf_2_3_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_5_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_181_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold30 hold30/A VGND VGND VPWR VPWR hold30/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 hold41/A VGND VGND VPWR VPWR hold41/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold52 hold52/A VGND VGND VPWR VPWR hold52/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold63 hold63/A VGND VGND VPWR VPWR hold63/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 hold74/A VGND VGND VPWR VPWR hold74/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 hold85/A VGND VGND VPWR VPWR hold85/X sky130_fd_sc_hd__buf_6
Xhold96 hold96/A VGND VGND VPWR VPWR hold96/X sky130_fd_sc_hd__buf_6
XFILLER_29_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_5 _5268_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3240_ _4621_/B VGND VGND VPWR VPWR _4610_/A sky130_fd_sc_hd__clkinv_2
XFILLER_100_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6930_ _7130_/CLK _6930_/D fanout519/X VGND VGND VPWR VPWR _6930_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_35_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6861_ _7110_/CLK _6861_/D fanout507/X VGND VGND VPWR VPWR _6861_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_6_csclk _7018_/CLK VGND VGND VPWR VPWR _6755_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_34_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5812_ _6895_/Q _5655_/X _5688_/X _6863_/Q _5811_/X VGND VGND VPWR VPWR _5813_/D
+ sky130_fd_sc_hd__a221o_1
X_6792_ _7209_/CLK _6792_/D fanout484/X VGND VGND VPWR VPWR _6792_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5743_ _6972_/Q _5960_/B VGND VGND VPWR VPWR _5743_/X sky130_fd_sc_hd__or2_1
XFILLER_148_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5674_ _6930_/Q _5670_/X _5673_/X VGND VGND VPWR VPWR _5681_/C sky130_fd_sc_hd__a21o_1
X_4625_ _5021_/B _4679_/B VGND VGND VPWR VPWR _5177_/A sky130_fd_sc_hd__nor2_1
XFILLER_148_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold500 _7110_/Q VGND VGND VPWR VPWR hold500/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold511 _5267_/X VGND VGND VPWR VPWR _6857_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4556_ _4556_/A VGND VGND VPWR VPWR _4783_/A sky130_fd_sc_hd__inv_2
Xhold522 _7210_/Q VGND VGND VPWR VPWR hold522/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold533 _5301_/X VGND VGND VPWR VPWR _6887_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3507_ _3726_/B _3507_/B VGND VGND VPWR VPWR _4034_/A sky130_fd_sc_hd__nor2_4
Xhold544 _6853_/Q VGND VGND VPWR VPWR hold544/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 _5312_/X VGND VGND VPWR VPWR _6897_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold566 _5204_/X VGND VGND VPWR VPWR _6806_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4487_ _4759_/A _4846_/D VGND VGND VPWR VPWR _4530_/B sky130_fd_sc_hd__nand2_2
Xhold577 _6719_/Q VGND VGND VPWR VPWR hold577/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold588 _5346_/X VGND VGND VPWR VPWR _6927_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6226_ _6521_/Q _5994_/X _5998_/Y _6761_/Q _6223_/X VGND VGND VPWR VPWR _6232_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3438_ _6895_/Q _5304_/A _5502_/A _7071_/Q _3425_/X VGND VGND VPWR VPWR _3446_/B
+ sky130_fd_sc_hd__a221o_1
Xhold599 _7079_/Q VGND VGND VPWR VPWR hold599/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6157_ _7140_/Q _6308_/A2 _6338_/B1 _7100_/Q _6147_/X VGND VGND VPWR VPWR _6157_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3369_ _6889_/Q _3318_/Y _5358_/A _6945_/Q VGND VGND VPWR VPWR _3369_/X sky130_fd_sc_hd__a22o_1
Xhold1200 _5556_/X VGND VGND VPWR VPWR _7113_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1211 _6793_/Q VGND VGND VPWR VPWR _5188_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5108_ _5108_/A _5108_/B VGND VGND VPWR VPWR _5109_/D sky130_fd_sc_hd__nor2_1
Xhold1222 _6616_/Q VGND VGND VPWR VPWR _4154_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1233 _5377_/X VGND VGND VPWR VPWR _6954_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6088_ _7060_/Q _6205_/B1 _6206_/B1 _6980_/Q VGND VGND VPWR VPWR _6088_/X sky130_fd_sc_hd__a22o_1
Xhold1244 _6970_/Q VGND VGND VPWR VPWR _5395_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1255 _4160_/X VGND VGND VPWR VPWR _6621_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1266 _5521_/X VGND VGND VPWR VPWR _7082_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1277 _6511_/Q VGND VGND VPWR VPWR _4017_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5039_ _5039_/A _5039_/B _5038_/X VGND VGND VPWR VPWR _5039_/X sky130_fd_sc_hd__or3b_1
XTAP_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1288 _3968_/X VGND VGND VPWR VPWR _6474_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1299 _6482_/Q VGND VGND VPWR VPWR _3984_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_578 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput120 wb_adr_i[29] VGND VGND VPWR VPWR input120/X sky130_fd_sc_hd__clkbuf_1
Xinput131 wb_cyc_i VGND VGND VPWR VPWR input131/X sky130_fd_sc_hd__clkbuf_1
XFILLER_163_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput142 wb_dat_i[19] VGND VGND VPWR VPWR _6372_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput153 wb_dat_i[29] VGND VGND VPWR VPWR _6379_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput164 wb_rstn_i VGND VGND VPWR VPWR input164/X sky130_fd_sc_hd__clkbuf_4
XFILLER_48_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4410_ _4433_/C _4436_/B VGND VGND VPWR VPWR _5001_/A sky130_fd_sc_hd__and2b_1
XFILLER_184_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5390_ _5567_/A0 hold765/X _5393_/S VGND VGND VPWR VPWR _5390_/X sky130_fd_sc_hd__mux2_1
X_4341_ _4605_/A _4621_/B VGND VGND VPWR VPWR _4341_/X sky130_fd_sc_hd__and2_2
XFILLER_113_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7060_ _7075_/CLK _7060_/D fanout515/X VGND VGND VPWR VPWR _7060_/Q sky130_fd_sc_hd__dfrtp_4
X_4272_ hold297/X _5459_/A0 _4275_/S VGND VGND VPWR VPWR _4272_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6011_ _7002_/Q _6006_/Y _6007_/Y _7103_/Q _6010_/X VGND VGND VPWR VPWR _6012_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_140_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3223_ _6933_/Q VGND VGND VPWR VPWR _3223_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6913_ _7138_/CLK _6913_/D fanout524/X VGND VGND VPWR VPWR _6913_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6844_ _7110_/CLK _6844_/D fanout505/X VGND VGND VPWR VPWR _6844_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6775_ _6986_/CLK _6775_/D fanout491/X VGND VGND VPWR VPWR _6775_/Q sky130_fd_sc_hd__dfrtp_4
X_3987_ hold591/X _6396_/A0 _3991_/S VGND VGND VPWR VPWR _3987_/X sky130_fd_sc_hd__mux2_1
X_5726_ _6947_/Q _5666_/X _5688_/X _6859_/Q VGND VGND VPWR VPWR _5726_/X sky130_fd_sc_hd__a22o_1
XFILLER_109_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5657_ _6890_/Q _5655_/X _5656_/X _6994_/Q VGND VGND VPWR VPWR _5657_/X sky130_fd_sc_hd__a22o_1
XFILLER_136_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4608_ _4792_/A _4797_/A _4607_/X VGND VGND VPWR VPWR _4644_/B sky130_fd_sc_hd__a21o_1
XFILLER_184_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5588_ hold40/X _5588_/A1 hold70/X VGND VGND VPWR VPWR hold71/A sky130_fd_sc_hd__mux2_1
Xhold330 _4123_/X VGND VGND VPWR VPWR _6590_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_163_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold341 _7027_/Q VGND VGND VPWR VPWR hold341/X sky130_fd_sc_hd__dlygate4sd3_1
X_4539_ _4819_/C _4971_/B VGND VGND VPWR VPWR _4553_/B sky130_fd_sc_hd__and2_1
Xhold352 _5297_/X VGND VGND VPWR VPWR _6883_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold363 _6669_/Q VGND VGND VPWR VPWR hold363/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 _5555_/X VGND VGND VPWR VPWR _7112_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold385 _6658_/Q VGND VGND VPWR VPWR hold385/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold396 _5510_/X VGND VGND VPWR VPWR _7073_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6209_ _7118_/Q _6322_/B1 _6030_/X _7001_/Q _6208_/X VGND VGND VPWR VPWR _6217_/B
+ sky130_fd_sc_hd__a221o_1
X_7189_ _7193_/CLK _7189_/D VGND VGND VPWR VPWR _7189_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1030 _5554_/X VGND VGND VPWR VPWR _7111_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1041 _6498_/Q VGND VGND VPWR VPWR _4002_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1052 _5314_/X VGND VGND VPWR VPWR _6898_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1063 _7026_/Q VGND VGND VPWR VPWR _5458_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1074 _5350_/X VGND VGND VPWR VPWR _6930_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1085 hold1453/X VGND VGND VPWR VPWR _5494_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_203 _5699_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1096 _6538_/Q VGND VGND VPWR VPWR _4049_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_214 _3957_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_225 _6027_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_236 _5581_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_247 _5685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_258 _3937_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_71_csclk _6753_/CLK VGND VGND VPWR VPWR _6825_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_64_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3910_ _3906_/X _3908_/Y _6565_/Q _3896_/B VGND VGND VPWR VPWR _6565_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_32_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4890_ _5174_/A _4890_/B _4890_/C _4890_/D VGND VGND VPWR VPWR _4890_/X sky130_fd_sc_hd__or4_1
X_3841_ _3913_/B1 _3795_/Y _6459_/Q VGND VGND VPWR VPWR _3841_/X sky130_fd_sc_hd__a21o_1
XFILLER_60_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3772_ _6793_/Q _5187_/A _3767_/X _3769_/X _3771_/X VGND VGND VPWR VPWR _3789_/B
+ sky130_fd_sc_hd__a2111o_1
X_6560_ _6664_/CLK _6560_/D _6426_/A VGND VGND VPWR VPWR _6560_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_9_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5511_ _5511_/A _5535_/B VGND VGND VPWR VPWR _5519_/S sky130_fd_sc_hd__nand2_8
X_6491_ _6759_/CLK _6491_/D fanout488/X VGND VGND VPWR VPWR _6491_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_118_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5442_ _5583_/A0 hold245/X _5447_/S VGND VGND VPWR VPWR _5442_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5373_ _5550_/A0 hold569/X _5375_/S VGND VGND VPWR VPWR _5373_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_24_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7129_/CLK sky130_fd_sc_hd__clkbuf_16
X_7112_ _7137_/CLK _7112_/D fanout501/X VGND VGND VPWR VPWR _7112_/Q sky130_fd_sc_hd__dfstp_1
X_4324_ _4324_/A _5535_/B VGND VGND VPWR VPWR _4329_/S sky130_fd_sc_hd__and2_2
XFILLER_160_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7043_ _7043_/CLK _7043_/D fanout514/X VGND VGND VPWR VPWR _7043_/Q sky130_fd_sc_hd__dfstp_1
X_4255_ hold829/X _4327_/A1 _4257_/S VGND VGND VPWR VPWR _4255_/X sky130_fd_sc_hd__mux2_1
X_3206_ _7069_/Q VGND VGND VPWR VPWR _3206_/Y sky130_fd_sc_hd__inv_2
X_4186_ _4186_/A0 _3447_/X _4188_/S VGND VGND VPWR VPWR _6644_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_39_csclk _6931_/CLK VGND VGND VPWR VPWR _7079_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_95_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_1_0_csclk clkbuf_3_1_0_csclk/A VGND VGND VPWR VPWR _7018_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_82_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6827_ _7136_/CLK _6827_/D fanout520/X VGND VGND VPWR VPWR _6827_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6758_ _6760_/CLK _6758_/D fanout490/X VGND VGND VPWR VPWR _6758_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_149_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5709_ _6842_/Q _5691_/Y _5708_/X _5681_/X _5650_/Y VGND VGND VPWR VPWR _5709_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_148_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6689_ _7094_/CLK _6689_/D fanout494/X VGND VGND VPWR VPWR _6689_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_109_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold160 _5515_/X VGND VGND VPWR VPWR _7077_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold171 _7131_/Q VGND VGND VPWR VPWR hold171/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold182 _4163_/X VGND VGND VPWR VPWR _6624_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold193 hold193/A VGND VGND VPWR VPWR hold193/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_120_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4040_ _4040_/A _4330_/B VGND VGND VPWR VPWR _4045_/S sky130_fd_sc_hd__nand2_2
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5991_ _6019_/A _6039_/C _6030_/C VGND VGND VPWR VPWR _6029_/B sky130_fd_sc_hd__and3b_2
XFILLER_91_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4942_ _4942_/A _5023_/B VGND VGND VPWR VPWR _5060_/B sky130_fd_sc_hd__nand2_1
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4873_ _5050_/A _5050_/B VGND VGND VPWR VPWR _4873_/Y sky130_fd_sc_hd__nand2_1
XFILLER_178_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6612_ _6664_/CLK _6612_/D _6426_/A VGND VGND VPWR VPWR _6612_/Q sky130_fd_sc_hd__dfrtp_1
X_3824_ hold64/A hold72/A _3816_/Y _3823_/X VGND VGND VPWR VPWR _3824_/X sky130_fd_sc_hd__a22o_1
XFILLER_177_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6543_ _3945_/A1 _6543_/D _6431_/X VGND VGND VPWR VPWR _6543_/Q sky130_fd_sc_hd__dfrtp_4
X_3755_ _3755_/A _3755_/B _3755_/C _3755_/D VGND VGND VPWR VPWR _3790_/B sky130_fd_sc_hd__or4_1
XFILLER_192_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3686_ _7003_/Q _5430_/A _4034_/A _6527_/Q VGND VGND VPWR VPWR _3686_/X sky130_fd_sc_hd__a22o_1
X_6474_ _6825_/CLK _6474_/D fanout490/X VGND VGND VPWR VPWR _6474_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_145_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5425_ _5539_/A1 hold279/X _5429_/S VGND VGND VPWR VPWR _5425_/X sky130_fd_sc_hd__mux2_1
Xoutput210 _3227_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[7] sky130_fd_sc_hd__buf_12
Xoutput221 _6547_/Q VGND VGND VPWR VPWR mgmt_gpio_out[17] sky130_fd_sc_hd__buf_12
XFILLER_133_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput232 _6829_/Q VGND VGND VPWR VPWR mgmt_gpio_out[27] sky130_fd_sc_hd__buf_12
Xoutput243 _3918_/X VGND VGND VPWR VPWR mgmt_gpio_out[37] sky130_fd_sc_hd__buf_12
Xoutput254 _3944_/Y VGND VGND VPWR VPWR pad_flash_csb_oeb sky130_fd_sc_hd__buf_12
X_5356_ _5578_/A0 hold832/X _5357_/S VGND VGND VPWR VPWR _5356_/X sky130_fd_sc_hd__mux2_1
Xoutput265 _6792_/Q VGND VGND VPWR VPWR pll_dco_ena sky130_fd_sc_hd__buf_12
Xoutput276 _6484_/Q VGND VGND VPWR VPWR pll_trim[10] sky130_fd_sc_hd__buf_12
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput287 _6478_/Q VGND VGND VPWR VPWR pll_trim[20] sky130_fd_sc_hd__buf_12
X_4307_ _5212_/C hold960/X _4311_/S VGND VGND VPWR VPWR _4307_/X sky130_fd_sc_hd__mux2_1
Xoutput298 _6497_/Q VGND VGND VPWR VPWR pll_trim[7] sky130_fd_sc_hd__buf_12
X_5287_ hold565/X hold775/X hold32/X VGND VGND VPWR VPWR _5287_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7026_ _7074_/CLK _7026_/D fanout501/X VGND VGND VPWR VPWR _7026_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_87_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4238_ hold36/X _4238_/A1 hold59/X VGND VGND VPWR VPWR hold60/A sky130_fd_sc_hd__mux2_1
XFILLER_28_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4169_ _4169_/A0 _3601_/X _4173_/S VGND VGND VPWR VPWR _6629_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire359 _6094_/A VGND VGND VPWR VPWR _6292_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_136_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout470 _5581_/A0 VGND VGND VPWR VPWR _5521_/A0 sky130_fd_sc_hd__buf_6
XFILLER_59_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout481 _6440_/B VGND VGND VPWR VPWR _6441_/B sky130_fd_sc_hd__buf_4
XFILLER_120_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout492 _6432_/A VGND VGND VPWR VPWR _6433_/A sky130_fd_sc_hd__buf_4
XFILLER_65_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3540_ input30/X _3304_/Y _3751_/A2 _3961_/B _3539_/X VGND VGND VPWR VPWR _3541_/D
+ sky130_fd_sc_hd__a221o_2
Xhold907 _5587_/X VGND VGND VPWR VPWR _7141_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold918 _6834_/Q VGND VGND VPWR VPWR hold918/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3471_ _3476_/A _3471_/B VGND VGND VPWR VPWR _3471_/Y sky130_fd_sc_hd__nor2_4
Xhold929 _5261_/X VGND VGND VPWR VPWR _6851_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5210_ _5210_/A _6392_/B VGND VGND VPWR VPWR _5211_/S sky130_fd_sc_hd__nand2_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6190_ _6952_/Q _6024_/A _6009_/X _6976_/Q VGND VGND VPWR VPWR _6190_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5141_ _4872_/A _4728_/Y _4916_/A _4618_/C VGND VGND VPWR VPWR _5141_/X sky130_fd_sc_hd__o211a_1
XFILLER_69_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5072_ _4645_/X _4665_/B _4668_/X _4693_/A VGND VGND VPWR VPWR _5072_/X sky130_fd_sc_hd__a31o_1
Xhold1607 _6839_/Q VGND VGND VPWR VPWR hold441/A sky130_fd_sc_hd__dlygate4sd3_1
X_4023_ _4023_/A0 _6393_/A0 _4027_/S VGND VGND VPWR VPWR _4023_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5974_ _7157_/Q _7158_/Q VGND VGND VPWR VPWR _6020_/C sky130_fd_sc_hd__nor2_4
XFILLER_80_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4925_ _5095_/A _4925_/B _4924_/Y VGND VGND VPWR VPWR _4925_/X sky130_fd_sc_hd__or3b_1
XFILLER_100_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4856_ _4759_/A _4395_/Y _4502_/A _4833_/Y VGND VGND VPWR VPWR _4857_/D sky130_fd_sc_hd__a211oi_1
XFILLER_178_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3807_ hold64/A hold53/A hold25/A VGND VGND VPWR VPWR _3823_/B sky130_fd_sc_hd__and3_1
XFILLER_119_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4787_ _5076_/B _4689_/B _4770_/C VGND VGND VPWR VPWR _4982_/B sky130_fd_sc_hd__o21bai_2
XFILLER_119_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6526_ _7207_/CLK _6526_/D fanout484/X VGND VGND VPWR VPWR _6526_/Q sky130_fd_sc_hd__dfrtp_2
X_3738_ _6858_/Q _5268_/A _5340_/A _6922_/Q VGND VGND VPWR VPWR _3738_/X sky130_fd_sc_hd__a22o_1
XFILLER_109_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6457_ _3927_/A1 _6457_/D _6412_/X VGND VGND VPWR VPWR _6457_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_161_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3669_ _3669_/A _3669_/B _3669_/C _3669_/D VGND VGND VPWR VPWR _3723_/A sky130_fd_sc_hd__or4_1
XFILLER_118_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5408_ _5549_/A0 hold637/X _5411_/S VGND VGND VPWR VPWR _5408_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6388_ _6700_/Q _6357_/A _6358_/B _6698_/Q VGND VGND VPWR VPWR _6388_/X sky130_fd_sc_hd__a22o_1
X_5339_ _5579_/A0 hold506/X _5339_/S VGND VGND VPWR VPWR _5339_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_554 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7009_ _7080_/CLK _7009_/D fanout502/X VGND VGND VPWR VPWR _7009_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_75_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_719 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4710_ _4832_/B _4677_/B _4689_/B _5076_/A _4709_/X VGND VGND VPWR VPWR _4710_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_30_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5690_ _5938_/B _5705_/B _5703_/B VGND VGND VPWR VPWR _5690_/X sky130_fd_sc_hd__and3_4
XFILLER_147_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4641_ _4639_/A _4639_/B _4689_/B _5076_/B _4640_/X VGND VGND VPWR VPWR _4642_/D
+ sky130_fd_sc_hd__o221a_1
X_4572_ _5021_/A _4981_/B _4571_/X VGND VGND VPWR VPWR _4572_/Y sky130_fd_sc_hd__o21ai_1
Xmax_cap401 _5980_/Y VGND VGND VPWR VPWR _6027_/A sky130_fd_sc_hd__buf_12
XFILLER_116_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold704 _4244_/X VGND VGND VPWR VPWR _6689_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6311_ _6673_/Q _6340_/A2 wire394/X _6637_/Q _6310_/X VGND VGND VPWR VPWR _6315_/B
+ sky130_fd_sc_hd__a221o_1
Xmax_cap423 _5642_/X VGND VGND VPWR VPWR _6323_/A2 sky130_fd_sc_hd__buf_12
Xhold715 _6520_/Q VGND VGND VPWR VPWR hold715/X sky130_fd_sc_hd__dlygate4sd3_1
X_3523_ _6502_/Q _3778_/A2 _5295_/A _6886_/Q _3522_/X VGND VGND VPWR VPWR _3524_/D
+ sky130_fd_sc_hd__a221o_1
Xhold726 _3982_/X VGND VGND VPWR VPWR _6481_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold737 _6505_/Q VGND VGND VPWR VPWR hold737/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold748 _4044_/X VGND VGND VPWR VPWR _6534_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6242_ _6292_/A _6242_/B _6242_/C _6242_/D VGND VGND VPWR VPWR _6242_/X sky130_fd_sc_hd__or4_1
Xhold759 _6614_/Q VGND VGND VPWR VPWR hold759/X sky130_fd_sc_hd__dlygate4sd3_1
X_3454_ _3528_/B hold49/X VGND VGND VPWR VPWR _4240_/A sky130_fd_sc_hd__nor2_4
Xmax_cap478 _4732_/A VGND VGND VPWR VPWR _4999_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_130_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3385_ _7080_/Q _5511_/A _5430_/A _7008_/Q VGND VGND VPWR VPWR _3385_/X sky130_fd_sc_hd__a22o_1
X_6173_ _6968_/Q _6025_/D _6212_/B1 _7048_/Q _6172_/X VGND VGND VPWR VPWR _6180_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_97_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5124_ _5124_/A _5124_/B _5124_/C _4708_/B VGND VGND VPWR VPWR _5125_/B sky130_fd_sc_hd__or4b_1
Xhold1404 _7195_/Q VGND VGND VPWR VPWR hold1404/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1415 _7196_/Q VGND VGND VPWR VPWR _6356_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1426 _6630_/Q VGND VGND VPWR VPWR _4170_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1437 _6779_/Q VGND VGND VPWR VPWR _3258_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5055_ _5126_/B _5162_/B _5126_/C _5162_/C VGND VGND VPWR VPWR _5067_/B sky130_fd_sc_hd__or4_1
XFILLER_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1448 _6708_/Q VGND VGND VPWR VPWR hold829/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1459 _5222_/X VGND VGND VPWR VPWR hold968/A sky130_fd_sc_hd__dlygate4sd3_1
X_4006_ hold85/X hold167/X _4009_/S VGND VGND VPWR VPWR _4006_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5957_ _5957_/A _5957_/B _5957_/C _5957_/D VGND VGND VPWR VPWR _5957_/X sky130_fd_sc_hd__or4_1
X_4908_ _4832_/B _5108_/A _5021_/B _4677_/B VGND VGND VPWR VPWR _4915_/C sky130_fd_sc_hd__o22ai_1
XFILLER_21_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5888_ _6517_/Q _5966_/B1 _5887_/X VGND VGND VPWR VPWR _5891_/C sky130_fd_sc_hd__a21o_1
XFILLER_178_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4839_ _4839_/A _4839_/B VGND VGND VPWR VPWR _5127_/B sky130_fd_sc_hd__nor2_1
XFILLER_138_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6509_ _6708_/CLK _6509_/D _6432_/A VGND VGND VPWR VPWR _6509_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_134_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold20 hold20/A VGND VGND VPWR VPWR hold20/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold31 hold31/A VGND VGND VPWR VPWR hold31/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold42 hold42/A VGND VGND VPWR VPWR hold42/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 hold53/A VGND VGND VPWR VPWR hold53/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold64 hold64/A VGND VGND VPWR VPWR hold64/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 hold75/A VGND VGND VPWR VPWR hold75/X sky130_fd_sc_hd__buf_6
Xhold86 hold86/A VGND VGND VPWR VPWR hold86/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 hold97/A VGND VGND VPWR VPWR hold97/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_6 _4120_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6860_ _7136_/CLK _6860_/D fanout520/X VGND VGND VPWR VPWR _6860_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_35_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5811_ _6919_/Q _5677_/X _5694_/X _7079_/Q VGND VGND VPWR VPWR _5811_/X sky130_fd_sc_hd__a22o_1
XFILLER_62_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6791_ _7209_/CLK _6791_/D fanout484/X VGND VGND VPWR VPWR _6791_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5742_ _7012_/Q _5686_/X _5966_/B1 _7036_/Q _5741_/X VGND VGND VPWR VPWR _5750_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_50_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5673_ _7058_/Q _5671_/X _5955_/A2 _6922_/Q VGND VGND VPWR VPWR _5673_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4624_ _4814_/A _4639_/B VGND VGND VPWR VPWR _4679_/B sky130_fd_sc_hd__or2_4
XFILLER_163_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold501 _5552_/X VGND VGND VPWR VPWR _7110_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4555_ _4802_/B _4802_/C VGND VGND VPWR VPWR _4556_/A sky130_fd_sc_hd__nor2_1
Xhold512 _6985_/Q VGND VGND VPWR VPWR hold512/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 _6396_/X VGND VGND VPWR VPWR _7210_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold534 _6796_/Q VGND VGND VPWR VPWR hold534/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3506_ _6862_/Q _5268_/A _4153_/A _6620_/Q _3505_/X VGND VGND VPWR VPWR _3515_/B
+ sky130_fd_sc_hd__a221o_1
Xhold545 _5263_/X VGND VGND VPWR VPWR _6853_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold556 _7005_/Q VGND VGND VPWR VPWR hold556/X sky130_fd_sc_hd__dlygate4sd3_1
X_4486_ _4996_/A _4942_/A VGND VGND VPWR VPWR _5065_/A sky130_fd_sc_hd__nor2_1
Xhold567 _6865_/Q VGND VGND VPWR VPWR hold567/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 _4268_/X VGND VGND VPWR VPWR _6719_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6225_ _6611_/Q _6023_/C _6020_/X _6706_/Q VGND VGND VPWR VPWR _6241_/B sky130_fd_sc_hd__a22o_1
Xhold589 _6863_/Q VGND VGND VPWR VPWR hold589/X sky130_fd_sc_hd__dlygate4sd3_1
X_3437_ _6959_/Q _3320_/Y _4083_/S _3957_/A _3436_/X VGND VGND VPWR VPWR _3446_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_106_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3368_ _7065_/Q _5493_/A _5259_/A _6857_/Q _3346_/X VGND VGND VPWR VPWR _3371_/C
+ sky130_fd_sc_hd__a221o_1
X_6156_ _6156_/A _6156_/B _6156_/C _6156_/D VGND VGND VPWR VPWR _6156_/X sky130_fd_sc_hd__or4_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1201 _6762_/Q VGND VGND VPWR VPWR _4320_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1212 _5188_/X VGND VGND VPWR VPWR _6793_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5107_ _5107_/A _5107_/B _5107_/C _4676_/X VGND VGND VPWR VPWR _5178_/B sky130_fd_sc_hd__or4b_1
Xhold1223 _4154_/X VGND VGND VPWR VPWR _6616_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1234 _6811_/Q VGND VGND VPWR VPWR _5211_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6087_ _6988_/Q _6203_/A2 _6336_/A2 _6956_/Q _6086_/X VGND VGND VPWR VPWR _6094_/B
+ sky130_fd_sc_hd__a221o_1
X_3299_ _3299_/A _3299_/B VGND VGND VPWR VPWR _3340_/B sky130_fd_sc_hd__nand2_8
Xhold1245 _5395_/X VGND VGND VPWR VPWR _6970_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1256 _6914_/Q VGND VGND VPWR VPWR _5332_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1267 _6601_/Q VGND VGND VPWR VPWR _4136_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1278 _4017_/X VGND VGND VPWR VPWR _6511_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5038_ _4396_/X _4668_/X _4836_/Y _4453_/A VGND VGND VPWR VPWR _5038_/X sky130_fd_sc_hd__a31o_1
Xhold1289 _7090_/Q VGND VGND VPWR VPWR _5530_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6989_ _7140_/CLK _6989_/D fanout523/X VGND VGND VPWR VPWR _6989_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput110 wb_adr_i[1] VGND VGND VPWR VPWR _4846_/A sky130_fd_sc_hd__buf_6
Xinput121 wb_adr_i[2] VGND VGND VPWR VPWR _4951_/A sky130_fd_sc_hd__clkbuf_2
Xinput132 wb_dat_i[0] VGND VGND VPWR VPWR _6363_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput143 wb_dat_i[1] VGND VGND VPWR VPWR _6367_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_49_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput154 wb_dat_i[2] VGND VGND VPWR VPWR _6370_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput165 wb_sel_i[0] VGND VGND VPWR VPWR _6360_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4340_ _4348_/A _4348_/B _4348_/C VGND VGND VPWR VPWR _4404_/B sky130_fd_sc_hd__and3_1
XFILLER_125_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4271_ _4271_/A0 _5521_/A0 _4275_/S VGND VGND VPWR VPWR _4271_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6010_ _6866_/Q _6023_/C _6009_/X _6970_/Q VGND VGND VPWR VPWR _6010_/X sky130_fd_sc_hd__a22o_1
X_3222_ _6941_/Q VGND VGND VPWR VPWR _3222_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6912_ _7134_/CLK hold3/X fanout524/X VGND VGND VPWR VPWR _6912_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6843_ _7012_/CLK _6843_/D fanout505/X VGND VGND VPWR VPWR _6843_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_62_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6774_ _6825_/CLK _6774_/D fanout498/X VGND VGND VPWR VPWR _6774_/Q sky130_fd_sc_hd__dfrtp_4
X_3986_ _3986_/A0 _6395_/A0 _3991_/S VGND VGND VPWR VPWR _3986_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5725_ _6995_/Q _5656_/X _5661_/X _6883_/Q _5724_/X VGND VGND VPWR VPWR _5728_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5656_ _7152_/Q _5706_/B _5703_/B VGND VGND VPWR VPWR _5656_/X sky130_fd_sc_hd__and3_4
XFILLER_191_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4607_ _4981_/C _4846_/C _4993_/A _4607_/D VGND VGND VPWR VPWR _4607_/X sky130_fd_sc_hd__and4b_1
X_5587_ _5587_/A0 hold906/X hold70/X VGND VGND VPWR VPWR _5587_/X sky130_fd_sc_hd__mux2_1
Xhold320 _5374_/X VGND VGND VPWR VPWR _6952_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold331 _6809_/Q VGND VGND VPWR VPWR hold331/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4538_ _4570_/B _4538_/B VGND VGND VPWR VPWR _5036_/A sky130_fd_sc_hd__nand2_8
XFILLER_190_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold342 _5459_/X VGND VGND VPWR VPWR _7027_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold353 _6859_/Q VGND VGND VPWR VPWR hold353/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold364 _4215_/X VGND VGND VPWR VPWR _6669_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold375 _6913_/Q VGND VGND VPWR VPWR hold375/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold386 _4202_/X VGND VGND VPWR VPWR _6658_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4469_ _4474_/A _4832_/B VGND VGND VPWR VPWR _4839_/A sky130_fd_sc_hd__or2_1
Xhold397 _6881_/Q VGND VGND VPWR VPWR hold397/X sky130_fd_sc_hd__dlygate4sd3_1
X_6208_ _7142_/Q _6308_/A2 _6338_/B1 _7102_/Q _6197_/X VGND VGND VPWR VPWR _6208_/X
+ sky130_fd_sc_hd__a221o_1
X_7188_ _7200_/CLK _7188_/D _6348_/B VGND VGND VPWR VPWR _7188_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_58_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6139_ _6862_/Q _6025_/A _6027_/D _6886_/Q _6138_/X VGND VGND VPWR VPWR _6142_/C
+ sky130_fd_sc_hd__a221o_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1020 _5319_/X VGND VGND VPWR VPWR _6903_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1031 _6890_/Q VGND VGND VPWR VPWR _5305_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1042 _4002_/X VGND VGND VPWR VPWR _6498_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_133_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1053 _6924_/Q VGND VGND VPWR VPWR _5343_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1064 _5458_/X VGND VGND VPWR VPWR _7026_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1075 _6978_/Q VGND VGND VPWR VPWR _5404_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1086 _6537_/Q VGND VGND VPWR VPWR _4048_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1097 _4049_/X VGND VGND VPWR VPWR _6538_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_204 _5982_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_215 _7214_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_226 wire394/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_237 _5581_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_248 _5693_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_259 hold36/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_5_csclk _7018_/CLK VGND VGND VPWR VPWR _7094_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_150_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3840_ _6460_/Q _6445_/Q _3840_/S VGND VGND VPWR VPWR _6460_/D sky130_fd_sc_hd__mux2_1
XFILLER_32_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3771_ _7058_/Q _3329_/Y _4040_/A _6531_/Q _3770_/X VGND VGND VPWR VPWR _3771_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_158_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5510_ _5579_/A0 hold395/X _5510_/S VGND VGND VPWR VPWR _5510_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6490_ _6759_/CLK _6490_/D fanout488/X VGND VGND VPWR VPWR _6490_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_9_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5441_ _5573_/A0 hold797/X _5447_/S VGND VGND VPWR VPWR _5441_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5372_ _5549_/A0 hold657/X _5375_/S VGND VGND VPWR VPWR _5372_/X sky130_fd_sc_hd__mux2_1
X_7111_ _7123_/CLK _7111_/D fanout527/X VGND VGND VPWR VPWR _7111_/Q sky130_fd_sc_hd__dfstp_1
X_4323_ hold713/X _6397_/A0 _4323_/S VGND VGND VPWR VPWR _4323_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7042_ _7042_/CLK _7042_/D fanout497/X VGND VGND VPWR VPWR _7042_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_101_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4254_ hold942/X _5531_/A1 _4257_/S VGND VGND VPWR VPWR _4254_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3205_ _7077_/Q VGND VGND VPWR VPWR _3205_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4185_ _6643_/Q _4185_/A1 _4188_/S VGND VGND VPWR VPWR _6643_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6826_ _7136_/CLK _6826_/D fanout520/X VGND VGND VPWR VPWR _6826_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_51_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6757_ _6759_/CLK _6757_/D fanout488/X VGND VGND VPWR VPWR _6757_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_149_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3969_ hold4/X hold7/X _3971_/S VGND VGND VPWR VPWR hold8/A sky130_fd_sc_hd__mux2_8
XFILLER_50_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5708_ _5708_/A _5708_/B _5708_/C _5708_/D VGND VGND VPWR VPWR _5708_/X sky130_fd_sc_hd__or4_1
XFILLER_109_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6688_ _7094_/CLK _6688_/D fanout496/X VGND VGND VPWR VPWR _6688_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_148_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5639_ _5634_/Y _5638_/Y _5643_/B VGND VGND VPWR VPWR _7157_/D sky130_fd_sc_hd__a21oi_1
XFILLER_164_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold150 _6739_/Q VGND VGND VPWR VPWR hold150/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 _6861_/Q VGND VGND VPWR VPWR hold161/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 _5576_/X VGND VGND VPWR VPWR _7131_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold183 _6961_/Q VGND VGND VPWR VPWR hold183/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 _4126_/X VGND VGND VPWR VPWR _6593_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5990_ _7050_/Q _5988_/X _6022_/B _6898_/Q VGND VGND VPWR VPWR _5990_/X sky130_fd_sc_hd__a22o_1
XFILLER_64_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4941_ _4459_/B _4446_/Y _4843_/B _4940_/Y VGND VGND VPWR VPWR _5126_/C sky130_fd_sc_hd__a211o_1
X_4872_ _4872_/A _4872_/B VGND VGND VPWR VPWR _4894_/C sky130_fd_sc_hd__nor2_1
XFILLER_178_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6611_ _6664_/CLK _6611_/D _6426_/A VGND VGND VPWR VPWR _6611_/Q sky130_fd_sc_hd__dfrtp_2
X_3823_ hold16/A _3823_/B VGND VGND VPWR VPWR _3823_/X sky130_fd_sc_hd__or2_1
X_6542_ _3945_/A1 _6542_/D _6430_/X VGND VGND VPWR VPWR _6542_/Q sky130_fd_sc_hd__dfrtp_1
X_3754_ _6946_/Q _5367_/A _4252_/A _6706_/Q _3738_/X VGND VGND VPWR VPWR _3755_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_158_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6473_ _3945_/A1 _6473_/D _6428_/X VGND VGND VPWR VPWR _6473_/Q sky130_fd_sc_hd__dfrtp_2
X_3685_ _7027_/Q _3326_/Y _4153_/A _6617_/Q _3684_/X VGND VGND VPWR VPWR _3688_/C
+ sky130_fd_sc_hd__a221o_2
X_5424_ _5583_/A0 hold239/X _5429_/S VGND VGND VPWR VPWR _5424_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput200 _3202_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[32] sky130_fd_sc_hd__buf_12
Xoutput211 _3226_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[8] sky130_fd_sc_hd__buf_12
Xoutput222 _6548_/Q VGND VGND VPWR VPWR mgmt_gpio_out[18] sky130_fd_sc_hd__buf_12
Xoutput233 _6830_/Q VGND VGND VPWR VPWR mgmt_gpio_out[28] sky130_fd_sc_hd__buf_12
Xoutput244 _6557_/Q VGND VGND VPWR VPWR mgmt_gpio_out[3] sky130_fd_sc_hd__buf_12
XFILLER_160_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5355_ _5586_/A0 hold989/X _5357_/S VGND VGND VPWR VPWR _5355_/X sky130_fd_sc_hd__mux2_1
Xoutput255 _3951_/X VGND VGND VPWR VPWR pad_flash_io0_do sky130_fd_sc_hd__buf_12
Xoutput266 _6793_/Q VGND VGND VPWR VPWR pll_div[0] sky130_fd_sc_hd__buf_12
Xoutput277 _6485_/Q VGND VGND VPWR VPWR pll_trim[11] sky130_fd_sc_hd__buf_12
X_4306_ _4306_/A _6392_/B VGND VGND VPWR VPWR _4311_/S sky130_fd_sc_hd__nand2_4
Xoutput288 _6479_/Q VGND VGND VPWR VPWR pll_trim[21] sky130_fd_sc_hd__buf_12
XFILLER_160_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput299 _6482_/Q VGND VGND VPWR VPWR pll_trim[8] sky130_fd_sc_hd__buf_12
XFILLER_99_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5286_ hold31/X _5313_/B VGND VGND VPWR VPWR hold32/A sky130_fd_sc_hd__nand2_4
XFILLER_141_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7025_ _7110_/CLK _7025_/D fanout507/X VGND VGND VPWR VPWR _7025_/Q sky130_fd_sc_hd__dfrtp_1
X_4237_ hold44/X _4237_/A1 hold59/X VGND VGND VPWR VPWR hold63/A sky130_fd_sc_hd__mux2_1
XFILLER_101_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4168_ _4168_/A0 _3660_/X _4173_/S VGND VGND VPWR VPWR _6628_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4099_ hold840/X _4098_/X _4103_/S VGND VGND VPWR VPWR _4099_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6809_ _7033_/CLK _6809_/D fanout503/X VGND VGND VPWR VPWR _6809_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_11_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_70_csclk _6753_/CLK VGND VGND VPWR VPWR _6986_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_124_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout460 hold43/X VGND VGND VPWR VPWR hold44/A sky130_fd_sc_hd__buf_4
XFILLER_93_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout471 hold565/X VGND VGND VPWR VPWR _5581_/A0 sky130_fd_sc_hd__buf_8
Xfanout482 _6407_/B VGND VGND VPWR VPWR _6440_/B sky130_fd_sc_hd__buf_4
XFILLER_46_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout493 fanout496/X VGND VGND VPWR VPWR _6432_/A sky130_fd_sc_hd__buf_6
XFILLER_58_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_23_csclk _6820_/CLK VGND VGND VPWR VPWR _7075_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_38_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7055_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold908 _6687_/Q VGND VGND VPWR VPWR hold908/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold919 _5242_/X VGND VGND VPWR VPWR _6834_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3470_ _6926_/Q _5340_/A _5322_/A _6910_/Q _3469_/X VGND VGND VPWR VPWR _3484_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5140_ _5140_/A _5140_/B _5119_/Y VGND VGND VPWR VPWR _5172_/B sky130_fd_sc_hd__or3b_1
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1608 _7156_/Q VGND VGND VPWR VPWR _5636_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5071_ _6362_/A _5112_/C _5071_/C VGND VGND VPWR VPWR _5156_/A sky130_fd_sc_hd__or3_1
XFILLER_96_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4022_ _4022_/A _4330_/B VGND VGND VPWR VPWR _4027_/S sky130_fd_sc_hd__and2_2
XFILLER_84_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5973_ _6019_/A _6006_/B VGND VGND VPWR VPWR _6023_/A sky130_fd_sc_hd__nor2_2
XFILLER_64_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4924_ _4924_/A _4924_/B VGND VGND VPWR VPWR _4924_/Y sky130_fd_sc_hd__nor2_1
XFILLER_178_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4855_ _4461_/B _5021_/B _4707_/B _4784_/A _4837_/X VGND VGND VPWR VPWR _4857_/C
+ sky130_fd_sc_hd__o221a_1
X_3806_ _6541_/Q _3806_/B VGND VGND VPWR VPWR _3833_/S sky130_fd_sc_hd__nand2b_4
XFILLER_166_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4786_ _4485_/A _4971_/A _4598_/B VGND VGND VPWR VPWR _4786_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_165_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6525_ _6708_/CLK _6525_/D _6441_/A VGND VGND VPWR VPWR _6525_/Q sky130_fd_sc_hd__dfrtp_4
X_3737_ _6665_/Q _4210_/A _4159_/A _6621_/Q VGND VGND VPWR VPWR _3737_/X sky130_fd_sc_hd__a22o_2
XFILLER_118_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6456_ _3927_/A1 _6456_/D _6411_/X VGND VGND VPWR VPWR _6456_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3668_ _7136_/Q hold69/A hold77/A _7043_/Q _3667_/X VGND VGND VPWR VPWR _3669_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_133_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5407_ _5557_/A0 hold603/X _5411_/S VGND VGND VPWR VPWR _5407_/X sky130_fd_sc_hd__mux2_1
X_6387_ _6387_/A1 _4230_/X _6362_/A _3191_/Y VGND VGND VPWR VPWR _7205_/D sky130_fd_sc_hd__o211a_2
X_3599_ _7085_/Q _5520_/A _4330_/A _6774_/Q _3598_/X VGND VGND VPWR VPWR _3600_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_88_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5338_ _5578_/A0 hold809/X _5339_/S VGND VGND VPWR VPWR _5338_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5269_ _5536_/A1 _5269_/A1 _5276_/S VGND VGND VPWR VPWR _5269_/X sky130_fd_sc_hd__mux2_1
X_7008_ _7080_/CLK _7008_/D fanout502/X VGND VGND VPWR VPWR _7008_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4640_ _4677_/B _5108_/A _5076_/B VGND VGND VPWR VPWR _4640_/X sky130_fd_sc_hd__a21o_1
XFILLER_30_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4571_ _4569_/B _4784_/A _4568_/X _4484_/A VGND VGND VPWR VPWR _4571_/X sky130_fd_sc_hd__o211a_1
XFILLER_190_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap402 _6022_/A VGND VGND VPWR VPWR _6320_/B1 sky130_fd_sc_hd__buf_8
X_6310_ _6668_/Q wire412/X _6016_/X _6684_/Q VGND VGND VPWR VPWR _6310_/X sky130_fd_sc_hd__a22o_1
Xmax_cap413 _6023_/C VGND VGND VPWR VPWR _6199_/B1 sky130_fd_sc_hd__buf_8
X_3522_ _7086_/Q _5520_/A _3329_/Y _7062_/Q VGND VGND VPWR VPWR _3522_/X sky130_fd_sc_hd__a22o_1
Xhold705 _6974_/Q VGND VGND VPWR VPWR hold705/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold716 _4027_/X VGND VGND VPWR VPWR _6520_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold727 _6704_/Q VGND VGND VPWR VPWR hold727/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold738 _4009_/X VGND VGND VPWR VPWR _6505_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6241_ _6241_/A _6241_/B _6241_/C _6241_/D VGND VGND VPWR VPWR _6242_/D sky130_fd_sc_hd__or4_1
Xhold749 _6758_/Q VGND VGND VPWR VPWR hold749/X sky130_fd_sc_hd__dlygate4sd3_1
X_3453_ _6902_/Q hold22/A _5529_/A _7094_/Q _3452_/X VGND VGND VPWR VPWR _3468_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_170_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap479 _4376_/B VGND VGND VPWR VPWR _4466_/B sky130_fd_sc_hd__clkbuf_2
X_6172_ _7056_/Q _5988_/X _6024_/D _6944_/Q VGND VGND VPWR VPWR _6172_/X sky130_fd_sc_hd__a22o_1
X_3384_ _6984_/Q _3341_/Y _3983_/A _6488_/Q VGND VGND VPWR VPWR _3384_/X sky130_fd_sc_hd__a22o_1
XFILLER_97_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5123_ _5123_/A _5123_/B _5123_/C VGND VGND VPWR VPWR _5123_/X sky130_fd_sc_hd__and3_1
Xhold1405 _6633_/Q VGND VGND VPWR VPWR hold1405/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1416 _6491_/Q VGND VGND VPWR VPWR hold1416/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1427 _6628_/Q VGND VGND VPWR VPWR _4168_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1438 _3299_/A VGND VGND VPWR VPWR _3303_/A sky130_fd_sc_hd__dlygate4sd3_1
X_5054_ _5054_/A _5054_/B VGND VGND VPWR VPWR _5162_/C sky130_fd_sc_hd__nand2_1
Xhold1449 _4255_/X VGND VGND VPWR VPWR _6708_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4005_ _5584_/A0 hold490/X _4009_/S VGND VGND VPWR VPWR _4005_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5956_ _6755_/Q _5664_/X _5670_/X _6679_/Q _5955_/X VGND VGND VPWR VPWR _5957_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4907_ _4984_/A _4983_/A _4986_/A _5079_/A VGND VGND VPWR VPWR _4915_/B sky130_fd_sc_hd__or4_1
XFILLER_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5887_ _6772_/Q _5663_/X _5667_/X _6617_/Q VGND VGND VPWR VPWR _5887_/X sky130_fd_sc_hd__a22o_1
XFILLER_138_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4838_ _4951_/B _4838_/B VGND VGND VPWR VPWR _4868_/A sky130_fd_sc_hd__and2_1
XFILLER_138_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4769_ _4446_/Y _4870_/B _4741_/X _5134_/A _4768_/X VGND VGND VPWR VPWR _4770_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_107_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6508_ _6664_/CLK _6508_/D _6426_/A VGND VGND VPWR VPWR _6508_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_193_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6439_ _6441_/A _6440_/B VGND VGND VPWR VPWR _6439_/X sky130_fd_sc_hd__and2_1
XFILLER_162_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold10 hold10/A VGND VGND VPWR VPWR hold10/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 hold21/A VGND VGND VPWR VPWR hold21/X sky130_fd_sc_hd__buf_8
XFILLER_102_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold32 hold32/A VGND VGND VPWR VPWR hold32/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 hold62/X VGND VGND VPWR VPWR hold43/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold54 hold54/A VGND VGND VPWR VPWR hold54/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 hold65/A VGND VGND VPWR VPWR hold65/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 hold76/A VGND VGND VPWR VPWR hold76/X sky130_fd_sc_hd__buf_8
XFILLER_188_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold87 hold87/A VGND VGND VPWR VPWR hold87/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold98 hold98/A VGND VGND VPWR VPWR hold98/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_7 hold22/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5810_ _6903_/Q _5693_/X _5703_/X _6855_/Q _5809_/X VGND VGND VPWR VPWR _5813_/C
+ sky130_fd_sc_hd__a221o_1
X_6790_ _3945_/A1 _6790_/D _6441_/X VGND VGND VPWR VPWR _6790_/Q sky130_fd_sc_hd__dfrtn_1
X_5741_ _6964_/Q _5675_/X _5702_/X _6980_/Q VGND VGND VPWR VPWR _5741_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5672_ _5938_/B _5699_/B _5699_/C VGND VGND VPWR VPWR _5672_/X sky130_fd_sc_hd__and3_4
XFILLER_187_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4623_ _4784_/B _4639_/B VGND VGND VPWR VPWR _4627_/C sky130_fd_sc_hd__nor2_1
XFILLER_148_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4554_ _4792_/A _4792_/C _4792_/B VGND VGND VPWR VPWR _4802_/C sky130_fd_sc_hd__o21bai_1
Xhold502 _6759_/Q VGND VGND VPWR VPWR hold502/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold513 _5411_/X VGND VGND VPWR VPWR _6985_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold524 _6889_/Q VGND VGND VPWR VPWR hold524/X sky130_fd_sc_hd__dlygate4sd3_1
X_3505_ _6659_/Q _4198_/A _4147_/A _6615_/Q VGND VGND VPWR VPWR _3505_/X sky130_fd_sc_hd__a22o_1
Xhold535 _5191_/X VGND VGND VPWR VPWR _6796_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 _6604_/Q VGND VGND VPWR VPWR hold546/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4485_ _4485_/A _4657_/C VGND VGND VPWR VPWR _4887_/C sky130_fd_sc_hd__nand2_1
XFILLER_116_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold557 _5434_/X VGND VGND VPWR VPWR _7005_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold568 _5276_/X VGND VGND VPWR VPWR _6865_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6224_ _6536_/Q _5988_/X _6022_/B _6655_/Q VGND VGND VPWR VPWR _6241_/A sky130_fd_sc_hd__a22o_1
Xhold579 _6750_/Q VGND VGND VPWR VPWR hold579/X sky130_fd_sc_hd__dlygate4sd3_1
X_3436_ _6943_/Q _5358_/A _5571_/A _7132_/Q VGND VGND VPWR VPWR _3436_/X sky130_fd_sc_hd__a22o_1
XFILLER_131_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6155_ _6975_/Q _6009_/X _6206_/B1 _6983_/Q _6154_/X VGND VGND VPWR VPWR _6156_/D
+ sky130_fd_sc_hd__a221o_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3367_ _7001_/Q _3300_/Y _5466_/A _7041_/Q _3345_/X VGND VGND VPWR VPWR _3371_/B
+ sky130_fd_sc_hd__a221o_2
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1202 _4320_/X VGND VGND VPWR VPWR _6762_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5106_ _5106_/A _5106_/B _5106_/C _5105_/X VGND VGND VPWR VPWR _5156_/C sky130_fd_sc_hd__or4b_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1213 _6533_/Q VGND VGND VPWR VPWR _4043_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6086_ _6972_/Q _6009_/X _6030_/X _6996_/Q VGND VGND VPWR VPWR _6086_/X sky130_fd_sc_hd__a22o_1
Xhold1224 _6866_/Q VGND VGND VPWR VPWR _5278_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_3298_ _3526_/A _3476_/A VGND VGND VPWR VPWR _3298_/Y sky130_fd_sc_hd__nor2_8
Xhold1235 _5211_/X VGND VGND VPWR VPWR _6811_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1246 _6721_/Q VGND VGND VPWR VPWR _4271_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1257 _5332_/X VGND VGND VPWR VPWR _6914_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5037_ _4485_/A _5035_/Y _5036_/Y _4876_/A VGND VGND VPWR VPWR _5136_/A sky130_fd_sc_hd__a22o_1
Xhold1268 _4136_/X VGND VGND VPWR VPWR _6601_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1279 _6665_/Q VGND VGND VPWR VPWR _4211_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6988_ _7137_/CLK _6988_/D fanout501/X VGND VGND VPWR VPWR _6988_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_15_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5939_ _6668_/Q _5677_/X _5689_/X _5938_/X VGND VGND VPWR VPWR _5939_/X sky130_fd_sc_hd__a22o_1
XFILLER_15_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput100 wb_adr_i[10] VGND VGND VPWR VPWR _4339_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput111 wb_adr_i[20] VGND VGND VPWR VPWR _4654_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_49_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput122 wb_adr_i[30] VGND VGND VPWR VPWR _3884_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_88_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput133 wb_dat_i[10] VGND VGND VPWR VPWR _6369_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput144 wb_dat_i[20] VGND VGND VPWR VPWR _6375_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput155 wb_dat_i[30] VGND VGND VPWR VPWR _6381_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput166 wb_sel_i[1] VGND VGND VPWR VPWR _6389_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_102_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_731 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4270_ _4270_/A _5580_/B VGND VGND VPWR VPWR _4275_/S sky130_fd_sc_hd__and2_2
XFILLER_113_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3221_ _6949_/Q VGND VGND VPWR VPWR _3221_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6911_ _7126_/CLK _6911_/D fanout524/X VGND VGND VPWR VPWR _6911_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_63_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6842_ _7068_/CLK _6842_/D fanout501/X VGND VGND VPWR VPWR _6842_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_62_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6773_ _6986_/CLK _6773_/D fanout491/X VGND VGND VPWR VPWR _6773_/Q sky130_fd_sc_hd__dfstp_1
X_3985_ _3985_/A0 _6394_/A0 _3991_/S VGND VGND VPWR VPWR _3985_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5724_ _6891_/Q _5655_/X _5667_/X _6875_/Q VGND VGND VPWR VPWR _5724_/X sky130_fd_sc_hd__a22o_1
X_5655_ _5938_/B _5700_/C _5699_/B VGND VGND VPWR VPWR _5655_/X sky130_fd_sc_hd__and3_4
XFILLER_148_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4606_ _4802_/C _4606_/B _4606_/C _4793_/B VGND VGND VPWR VPWR _4607_/D sky130_fd_sc_hd__and4b_1
X_5586_ _5586_/A0 hold999/X hold70/X VGND VGND VPWR VPWR _5586_/X sky130_fd_sc_hd__mux2_1
XFILLER_190_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold310 _5478_/X VGND VGND VPWR VPWR _7044_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 _6805_/Q VGND VGND VPWR VPWR hold321/X sky130_fd_sc_hd__dlygate4sd3_1
X_4537_ _4846_/A _4570_/B _4846_/B _4570_/D VGND VGND VPWR VPWR _4971_/B sky130_fd_sc_hd__and4_4
Xhold332 _5208_/X VGND VGND VPWR VPWR _6809_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold343 _6727_/Q VGND VGND VPWR VPWR hold343/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold354 _5270_/X VGND VGND VPWR VPWR _6859_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 _6659_/Q VGND VGND VPWR VPWR hold365/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold376 _5330_/X VGND VGND VPWR VPWR _6913_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4468_ _4489_/A _4484_/B _4352_/B VGND VGND VPWR VPWR _4940_/A sky130_fd_sc_hd__or3b_2
Xhold387 _6668_/Q VGND VGND VPWR VPWR hold387/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold398 _5294_/X VGND VGND VPWR VPWR _6881_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6207_ _7073_/Q _6272_/B _6202_/X _6204_/X _6206_/X VGND VGND VPWR VPWR _6207_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3419_ _6863_/Q _5268_/A _5340_/A _6927_/Q VGND VGND VPWR VPWR _3419_/X sky130_fd_sc_hd__a22o_1
X_7187_ _7187_/CLK _7187_/D fanout490/X VGND VGND VPWR VPWR _7187_/Q sky130_fd_sc_hd__dfrtp_1
X_4399_ _4420_/A _4596_/A VGND VGND VPWR VPWR _4400_/B sky130_fd_sc_hd__or2_2
XFILLER_98_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6138_ _6950_/Q _6024_/A _6212_/B1 _7046_/Q VGND VGND VPWR VPWR _6138_/X sky130_fd_sc_hd__a22o_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1010 _5337_/X VGND VGND VPWR VPWR _6919_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1021 _6983_/Q VGND VGND VPWR VPWR _5409_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1032 _5305_/X VGND VGND VPWR VPWR _6890_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1043 _6804_/Q VGND VGND VPWR VPWR _5201_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6069_ _6069_/A _6069_/B _6069_/C _6069_/D VGND VGND VPWR VPWR _6069_/X sky130_fd_sc_hd__or4_1
XFILLER_100_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1054 _5343_/X VGND VGND VPWR VPWR _6924_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1065 _7074_/Q VGND VGND VPWR VPWR _5512_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_133_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1076 _5404_/X VGND VGND VPWR VPWR _6978_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1087 _4048_/X VGND VGND VPWR VPWR _6537_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1098 hold1451/X VGND VGND VPWR VPWR _4207_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_205 _5988_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_216 _3958_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_227 _6329_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_238 hold9/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_249 _5705_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3770_ _6601_/Q _4135_/A _3547_/Y input98/X VGND VGND VPWR VPWR _3770_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5440_ hold565/X hold681/X _5447_/S VGND VGND VPWR VPWR _5440_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5371_ _5557_/A0 hold597/X _5375_/S VGND VGND VPWR VPWR _5371_/X sky130_fd_sc_hd__mux2_1
X_7110_ _7110_/CLK _7110_/D fanout507/X VGND VGND VPWR VPWR _7110_/Q sky130_fd_sc_hd__dfrtp_1
X_4322_ hold711/X _6396_/A0 _4323_/S VGND VGND VPWR VPWR _4322_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7041_ _7102_/CLK _7041_/D fanout503/X VGND VGND VPWR VPWR _7041_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_113_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4253_ _4253_/A0 _5476_/A0 _4257_/S VGND VGND VPWR VPWR _4253_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3204_ _7085_/Q VGND VGND VPWR VPWR _3204_/Y sky130_fd_sc_hd__inv_2
X_4184_ _4184_/A0 _3601_/X _4188_/S VGND VGND VPWR VPWR _6642_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_7_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A VGND VGND VPWR VPWR _7200_/CLK sky130_fd_sc_hd__clkbuf_8
X_6825_ _6825_/CLK _6825_/D fanout491/X VGND VGND VPWR VPWR _6825_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3968_ _3968_/A0 _5212_/C _3982_/S VGND VGND VPWR VPWR _3968_/X sky130_fd_sc_hd__mux2_1
X_6756_ _6759_/CLK _6756_/D fanout488/X VGND VGND VPWR VPWR _6756_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_149_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5707_ _6938_/Q _5705_/X _5706_/X _6498_/Q _5704_/X VGND VGND VPWR VPWR _5708_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6687_ _7094_/CLK _6687_/D fanout494/X VGND VGND VPWR VPWR _6687_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_109_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3899_ _5592_/B _3899_/B _7146_/Q _7147_/Q VGND VGND VPWR VPWR _3908_/B sky130_fd_sc_hd__and4b_1
XFILLER_149_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5638_ _7157_/Q _5643_/A VGND VGND VPWR VPWR _5638_/Y sky130_fd_sc_hd__nor2_1
XFILLER_164_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5569_ _5569_/A0 _5569_/A1 _5570_/S VGND VGND VPWR VPWR _5569_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold140 _6487_/Q VGND VGND VPWR VPWR hold140/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 _4292_/X VGND VGND VPWR VPWR _6739_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold162 _5272_/X VGND VGND VPWR VPWR _6861_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold173 hold173/A VGND VGND VPWR VPWR hold173/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 _5384_/X VGND VGND VPWR VPWR _6961_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 _6925_/Q VGND VGND VPWR VPWR hold195/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4940_ _4940_/A _5023_/B VGND VGND VPWR VPWR _4940_/Y sky130_fd_sc_hd__nor2_1
XFILLER_64_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4871_ _4871_/A _5094_/A VGND VGND VPWR VPWR _4871_/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3822_ _3821_/X _6467_/Q _3833_/S VGND VGND VPWR VPWR _6467_/D sky130_fd_sc_hd__mux2_1
X_6610_ _6963_/CLK _6610_/D fanout509/X VGND VGND VPWR VPWR _6610_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_177_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6541_ _3927_/A1 _6541_/D _6429_/X VGND VGND VPWR VPWR _6541_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_193_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3753_ _6736_/Q _4288_/A _5223_/A _6820_/Q _3732_/X VGND VGND VPWR VPWR _3755_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6472_ _3927_/A1 _6472_/D _6427_/X VGND VGND VPWR VPWR _6472_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_146_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3684_ _7075_/Q _5511_/A _3684_/B1 _7051_/Q VGND VGND VPWR VPWR _3684_/X sky130_fd_sc_hd__a22o_1
X_5423_ _5555_/A0 hold407/X _5429_/S VGND VGND VPWR VPWR _5423_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput201 _3201_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[33] sky130_fd_sc_hd__buf_12
Xoutput212 _3225_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[9] sky130_fd_sc_hd__buf_12
Xoutput223 _6549_/Q VGND VGND VPWR VPWR mgmt_gpio_out[19] sky130_fd_sc_hd__buf_12
X_5354_ hold85/X hold177/X _5357_/S VGND VGND VPWR VPWR _5354_/X sky130_fd_sc_hd__mux2_1
Xoutput234 _6831_/Q VGND VGND VPWR VPWR mgmt_gpio_out[29] sky130_fd_sc_hd__buf_12
Xoutput245 _6558_/Q VGND VGND VPWR VPWR mgmt_gpio_out[4] sky130_fd_sc_hd__buf_12
XFILLER_114_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput256 _3948_/A VGND VGND VPWR VPWR pad_flash_io0_ieb sky130_fd_sc_hd__buf_12
Xoutput267 _6794_/Q VGND VGND VPWR VPWR pll_div[1] sky130_fd_sc_hd__buf_12
X_4305_ _5549_/A0 hold579/X _4305_/S VGND VGND VPWR VPWR _4305_/X sky130_fd_sc_hd__mux2_1
Xoutput278 _6486_/Q VGND VGND VPWR VPWR pll_trim[12] sky130_fd_sc_hd__buf_12
Xoutput289 _6480_/Q VGND VGND VPWR VPWR pll_trim[22] sky130_fd_sc_hd__buf_12
X_5285_ _5579_/A0 hold518/X _5285_/S VGND VGND VPWR VPWR _5285_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7024_ _7080_/CLK _7024_/D fanout502/X VGND VGND VPWR VPWR _7024_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_101_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4236_ _5459_/A0 hold89/X hold59/X VGND VGND VPWR VPWR hold90/A sky130_fd_sc_hd__mux2_1
X_4167_ _4167_/A0 _3723_/X _4173_/S VGND VGND VPWR VPWR _6627_/D sky130_fd_sc_hd__mux2_1
X_4098_ hold441/X _5550_/A0 _4102_/S VGND VGND VPWR VPWR _4098_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_4_csclk clkbuf_leaf_4_csclk/A VGND VGND VPWR VPWR _6709_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6808_ _7033_/CLK _6808_/D fanout503/X VGND VGND VPWR VPWR _6808_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_168_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6739_ _6963_/CLK _6739_/D fanout510/X VGND VGND VPWR VPWR _6739_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_99_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout450 _5539_/A1 VGND VGND VPWR VPWR _5533_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout461 _5531_/A1 VGND VGND VPWR VPWR _6394_/A0 sky130_fd_sc_hd__buf_6
XFILLER_171_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout472 _5960_/B VGND VGND VPWR VPWR _5938_/B sky130_fd_sc_hd__buf_6
XFILLER_59_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout483 _3872_/Y VGND VGND VPWR VPWR _6407_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_120_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout494 fanout496/X VGND VGND VPWR VPWR fanout494/X sky130_fd_sc_hd__buf_8
XFILLER_19_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold909 _4242_/X VGND VGND VPWR VPWR _6687_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5070_ _6362_/A _5112_/C _5071_/C VGND VGND VPWR VPWR _5070_/Y sky130_fd_sc_hd__nor3_1
XFILLER_29_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1609 _7150_/Q VGND VGND VPWR VPWR _5620_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_4021_ _6397_/A0 hold560/X _4021_/S VGND VGND VPWR VPWR _4021_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5972_ _6000_/A _6039_/C VGND VGND VPWR VPWR _6006_/B sky130_fd_sc_hd__nand2_2
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4923_ _5153_/A _5109_/A _4963_/B _4923_/D VGND VGND VPWR VPWR _4924_/B sky130_fd_sc_hd__or4_1
XFILLER_178_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4854_ _4932_/A _5023_/B _4675_/A _4503_/C VGND VGND VPWR VPWR _4857_/B sky130_fd_sc_hd__o31a_1
X_3805_ _6543_/Q _3834_/B _3890_/B hold72/A VGND VGND VPWR VPWR _3806_/B sky130_fd_sc_hd__a31o_1
XFILLER_178_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4785_ _4759_/A _4485_/A _5015_/B VGND VGND VPWR VPWR _4785_/X sky130_fd_sc_hd__a21o_1
X_3736_ _7074_/Q _5511_/A _5448_/A _7018_/Q VGND VGND VPWR VPWR _3736_/X sky130_fd_sc_hd__a22o_1
X_6524_ _6708_/CLK _6524_/D _6432_/A VGND VGND VPWR VPWR _6524_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_174_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6455_ _3927_/A1 _6455_/D _6410_/X VGND VGND VPWR VPWR _6455_/Q sky130_fd_sc_hd__dfrtp_1
X_3667_ _6923_/Q _5340_/A _4010_/A _6507_/Q VGND VGND VPWR VPWR _3667_/X sky130_fd_sc_hd__a22o_1
XFILLER_109_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5406_ _5583_/A0 hold247/X _5411_/S VGND VGND VPWR VPWR _5406_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6386_ _6385_/X _6386_/A1 _6386_/S VGND VGND VPWR VPWR _7204_/D sky130_fd_sc_hd__mux2_1
X_3598_ _3872_/C _4085_/S _4264_/A _6719_/Q _3597_/X VGND VGND VPWR VPWR _3598_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_133_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5337_ _5586_/A0 _5337_/A1 _5339_/S VGND VGND VPWR VPWR _5337_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5268_ _5268_/A _5385_/B VGND VGND VPWR VPWR _5276_/S sky130_fd_sc_hd__nand2_8
X_4219_ hold44/X _4219_/A1 _4221_/S VGND VGND VPWR VPWR hold45/A sky130_fd_sc_hd__mux2_1
XFILLER_102_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7007_ _7071_/CLK _7007_/D fanout526/X VGND VGND VPWR VPWR _7007_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5199_ hold127/X hold175/X _5199_/S VGND VGND VPWR VPWR _5199_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4570_ _4846_/A _4570_/B _4846_/B _4570_/D VGND VGND VPWR VPWR _4814_/B sky130_fd_sc_hd__or4_4
X_3521_ _6918_/Q _5331_/A _5562_/A _7123_/Q VGND VGND VPWR VPWR _3524_/C sky130_fd_sc_hd__a22o_1
XFILLER_156_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap403 _6023_/A VGND VGND VPWR VPWR _6320_/A2 sky130_fd_sc_hd__buf_8
Xmax_cap414 _6027_/B VGND VGND VPWR VPWR _6340_/A2 sky130_fd_sc_hd__buf_12
Xhold706 _5399_/X VGND VGND VPWR VPWR _6974_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold717 _6615_/Q VGND VGND VPWR VPWR hold717/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold728 _4250_/X VGND VGND VPWR VPWR _6704_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6240_ _6601_/Q _5980_/Y _6036_/X _6516_/Q _6239_/X VGND VGND VPWR VPWR _6241_/D
+ sky130_fd_sc_hd__a221o_1
Xhold739 _7057_/Q VGND VGND VPWR VPWR hold739/X sky130_fd_sc_hd__dlygate4sd3_1
X_3452_ _7030_/Q _3326_/Y _4174_/A _6638_/Q VGND VGND VPWR VPWR _3452_/X sky130_fd_sc_hd__a22o_1
XFILLER_170_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6171_ _6195_/A2 _6170_/X _6171_/S VGND VGND VPWR VPWR _6171_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3383_ _6504_/Q _4001_/A _5439_/A _7016_/Q VGND VGND VPWR VPWR _3383_/X sky130_fd_sc_hd__a22o_1
X_5122_ _4582_/B _5016_/B _4504_/A _4504_/B VGND VGND VPWR VPWR _5123_/C sky130_fd_sc_hd__o211a_1
Xhold1406 _6641_/Q VGND VGND VPWR VPWR hold1406/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1417 _3994_/X VGND VGND VPWR VPWR _6491_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5053_ _5053_/A _5053_/B _5052_/X VGND VGND VPWR VPWR _5067_/A sky130_fd_sc_hd__or3b_1
Xhold1428 _6649_/Q VGND VGND VPWR VPWR _4192_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1439 _3528_/B VGND VGND VPWR VPWR _3471_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4004_ _5574_/A0 _4004_/A1 _4009_/S VGND VGND VPWR VPWR _4004_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5955_ _6674_/Q _5955_/A2 _5705_/X _6685_/Q VGND VGND VPWR VPWR _5955_/X sky130_fd_sc_hd__a22o_1
XFILLER_40_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4906_ _5021_/A _5023_/C _5021_/C VGND VGND VPWR VPWR _5079_/A sky130_fd_sc_hd__nor3_1
X_5886_ _6622_/Q _5661_/X _5697_/X _6732_/Q _5885_/X VGND VGND VPWR VPWR _5891_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_139_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4837_ _4652_/X _4836_/Y _4932_/A VGND VGND VPWR VPWR _4837_/X sky130_fd_sc_hd__a21o_1
XFILLER_178_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4768_ _4993_/A _4524_/B _4818_/B _4965_/B _4767_/X VGND VGND VPWR VPWR _4768_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_107_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6507_ _6707_/CLK _6507_/D _6433_/A VGND VGND VPWR VPWR _6507_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_134_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3719_ _7011_/Q _5439_/A _3471_/Y _6762_/Q VGND VGND VPWR VPWR _3719_/X sky130_fd_sc_hd__a22o_1
XFILLER_106_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4699_ _4699_/A _4699_/B _4860_/B _4699_/D VGND VGND VPWR VPWR _4699_/X sky130_fd_sc_hd__and4_1
XFILLER_134_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6438_ _6441_/A _6440_/B VGND VGND VPWR VPWR _6438_/X sky130_fd_sc_hd__and2_1
XFILLER_106_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6369_ _6698_/Q _6369_/A2 _6369_/B1 _6699_/Q VGND VGND VPWR VPWR _6369_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_22_csclk _6820_/CLK VGND VGND VPWR VPWR _7078_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold11 hold11/A VGND VGND VPWR VPWR hold11/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold22 hold22/A VGND VGND VPWR VPWR hold22/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold33 hold33/A VGND VGND VPWR VPWR hold33/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold44 hold44/A VGND VGND VPWR VPWR hold44/X sky130_fd_sc_hd__buf_4
Xhold55 hold55/A VGND VGND VPWR VPWR hold55/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 hold66/A VGND VGND VPWR VPWR hold66/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 hold77/A VGND VGND VPWR VPWR hold77/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 hold88/A VGND VGND VPWR VPWR hold88/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 hold99/A VGND VGND VPWR VPWR hold99/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_37_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7049_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_16_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_mgmt_gpio_in[4] mgmt_gpio_in[4] VGND VGND VPWR VPWR clkbuf_0_mgmt_gpio_in[4]/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_31_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_8 _5277_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_719 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5740_ _5740_/A _5740_/B _5740_/C _5740_/D VGND VGND VPWR VPWR _5740_/X sky130_fd_sc_hd__or4_1
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5671_ _7152_/Q _5706_/B _5699_/C VGND VGND VPWR VPWR _5671_/X sky130_fd_sc_hd__and3_4
XFILLER_188_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4622_ _4639_/B VGND VGND VPWR VPWR _4622_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4553_ _4935_/A _4553_/B VGND VGND VPWR VPWR _4792_/C sky130_fd_sc_hd__nor2_1
XFILLER_190_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold503 _4316_/X VGND VGND VPWR VPWR _6759_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold514 _6953_/Q VGND VGND VPWR VPWR hold514/X sky130_fd_sc_hd__dlygate4sd3_1
X_3504_ hold21/X _3538_/B VGND VGND VPWR VPWR _4147_/A sky130_fd_sc_hd__nor2_8
Xhold525 _5303_/X VGND VGND VPWR VPWR _6889_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold536 _6905_/Q VGND VGND VPWR VPWR hold536/X sky130_fd_sc_hd__dlygate4sd3_1
X_4484_ _4484_/A _4484_/B _4352_/B VGND VGND VPWR VPWR _4484_/X sky130_fd_sc_hd__or3b_1
Xhold547 _4139_/X VGND VGND VPWR VPWR _6604_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold558 _6620_/Q VGND VGND VPWR VPWR hold558/X sky130_fd_sc_hd__dlygate4sd3_1
X_6223_ _6511_/Q _5977_/X _6323_/B1 _6736_/Q VGND VGND VPWR VPWR _6223_/X sky130_fd_sc_hd__a22o_1
XFILLER_116_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold569 _6951_/Q VGND VGND VPWR VPWR hold569/X sky130_fd_sc_hd__dlygate4sd3_1
X_3435_ _6975_/Q _5394_/A _5277_/A _6871_/Q _3434_/X VGND VGND VPWR VPWR _3447_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_171_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6154_ _6959_/Q _6336_/A2 _6205_/B1 _7063_/Q VGND VGND VPWR VPWR _6154_/X sky130_fd_sc_hd__a22o_1
X_3366_ _6865_/Q _5268_/A _3983_/A _6489_/Q _3365_/X VGND VGND VPWR VPWR _3371_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1203 _6666_/Q VGND VGND VPWR VPWR _4212_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5105_ _4672_/A _5036_/A _5023_/C _5013_/A _4713_/A VGND VGND VPWR VPWR _5105_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1214 _4043_/X VGND VGND VPWR VPWR _6533_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6085_ _6085_/A _6085_/B VGND VGND VPWR VPWR _6085_/X sky130_fd_sc_hd__or2_2
XFILLER_58_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3297_ hold94/X _3301_/C hold18/X VGND VGND VPWR VPWR _3300_/A sky130_fd_sc_hd__or3b_4
Xhold1225 _5278_/X VGND VGND VPWR VPWR _6866_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1236 _6771_/Q VGND VGND VPWR VPWR _4331_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5036_ _5036_/A _5036_/B VGND VGND VPWR VPWR _5036_/Y sky130_fd_sc_hd__nand2_1
Xhold1247 _4271_/X VGND VGND VPWR VPWR _6721_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1258 hold1443/X VGND VGND VPWR VPWR _5503_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1269 _6706_/Q VGND VGND VPWR VPWR _4253_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6987_ _7139_/CLK _6987_/D fanout518/X VGND VGND VPWR VPWR _6987_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_179_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5938_ _6714_/Q _5938_/B VGND VGND VPWR VPWR _5938_/X sky130_fd_sc_hd__or2_1
XFILLER_179_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5869_ _5869_/A _5869_/B _5869_/C _5869_/D VGND VGND VPWR VPWR _5869_/X sky130_fd_sc_hd__or4_1
XFILLER_139_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput101 wb_adr_i[11] VGND VGND VPWR VPWR _4339_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_103_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput112 wb_adr_i[21] VGND VGND VPWR VPWR _4390_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_163_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput123 wb_adr_i[31] VGND VGND VPWR VPWR _3884_/A sky130_fd_sc_hd__clkbuf_1
Xinput134 wb_dat_i[11] VGND VGND VPWR VPWR _6372_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput145 wb_dat_i[21] VGND VGND VPWR VPWR _6378_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_102_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput156 wb_dat_i[31] VGND VGND VPWR VPWR _6384_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput167 wb_sel_i[2] VGND VGND VPWR VPWR _6358_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_76_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3220_ _6957_/Q VGND VGND VPWR VPWR _3220_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6910_ _7123_/CLK _6910_/D _6407_/A VGND VGND VPWR VPWR _6910_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6841_ _7140_/CLK hold82/X fanout522/X VGND VGND VPWR VPWR hold81/A sky130_fd_sc_hd__dfrtp_1
XFILLER_62_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6772_ _6986_/CLK _6772_/D fanout501/X VGND VGND VPWR VPWR _6772_/Q sky130_fd_sc_hd__dfrtp_1
X_3984_ _3984_/A0 _5212_/C _3991_/S VGND VGND VPWR VPWR _3984_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5723_ _7011_/Q _5686_/X _5703_/X _6851_/Q _5722_/X VGND VGND VPWR VPWR _5728_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_188_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5654_ _7148_/Q _7149_/Q VGND VGND VPWR VPWR _5699_/B sky130_fd_sc_hd__and2b_2
X_4605_ _4605_/A _4610_/A _5036_/A VGND VGND VPWR VPWR _4606_/C sky130_fd_sc_hd__or3_1
XFILLER_117_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5585_ hold85/X hold165/X hold70/X VGND VGND VPWR VPWR _5585_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold300 _4302_/X VGND VGND VPWR VPWR _6747_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold311 _6976_/Q VGND VGND VPWR VPWR hold311/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_191_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4536_ _4926_/A _4493_/X _4531_/X _4824_/A _4930_/A VGND VGND VPWR VPWR _4536_/Y
+ sky130_fd_sc_hd__a41oi_1
Xhold322 _5202_/X VGND VGND VPWR VPWR _6805_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold333 _6622_/Q VGND VGND VPWR VPWR hold333/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold344 _4278_/X VGND VGND VPWR VPWR _6727_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 _6818_/Q VGND VGND VPWR VPWR hold355/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 _4203_/X VGND VGND VPWR VPWR _6659_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4467_ _4467_/A _4654_/B _4467_/C VGND VGND VPWR VPWR _4484_/B sky130_fd_sc_hd__or3_2
Xhold377 _6685_/Q VGND VGND VPWR VPWR hold377/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold388 _4214_/X VGND VGND VPWR VPWR _6668_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6206_ _6977_/Q _6009_/X _6206_/B1 _6985_/Q _6205_/X VGND VGND VPWR VPWR _6206_/X
+ sky130_fd_sc_hd__a221o_1
Xhold399 _6833_/Q VGND VGND VPWR VPWR hold399/X sky130_fd_sc_hd__dlygate4sd3_1
X_3418_ _6951_/Q _5367_/A _5295_/A _6887_/Q VGND VGND VPWR VPWR _3418_/X sky130_fd_sc_hd__a22o_1
X_7186_ _7187_/CLK _7186_/D fanout490/X VGND VGND VPWR VPWR _7186_/Q sky130_fd_sc_hd__dfrtp_1
X_4398_ _4846_/A _4846_/B _4570_/D VGND VGND VPWR VPWR _4538_/B sky130_fd_sc_hd__and3_4
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3349_ _6505_/Q _3778_/A2 _3304_/Y input33/X VGND VGND VPWR VPWR _3349_/X sky130_fd_sc_hd__a22o_1
XFILLER_98_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6137_ _6926_/Q _6027_/B wire394/X _6894_/Q _6136_/X VGND VGND VPWR VPWR _6142_/B
+ sky130_fd_sc_hd__a221o_1
Xhold1000 _5586_/X VGND VGND VPWR VPWR _7140_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1011 _6975_/Q VGND VGND VPWR VPWR _5400_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1022 _5409_/X VGND VGND VPWR VPWR _6983_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1033 _7119_/Q VGND VGND VPWR VPWR _5563_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1044 _5201_/X VGND VGND VPWR VPWR _6804_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6068_ _6068_/A _6068_/B _6068_/C _6068_/D VGND VGND VPWR VPWR _6069_/D sky130_fd_sc_hd__or4_1
Xhold1055 _6884_/Q VGND VGND VPWR VPWR _5298_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1066 _5512_/X VGND VGND VPWR VPWR _7074_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1077 hold1515/X VGND VGND VPWR VPWR _5230_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1088 _6536_/Q VGND VGND VPWR VPWR _4047_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5019_ _5019_/A _5019_/B _5083_/C _5106_/B VGND VGND VPWR VPWR _5030_/A sky130_fd_sc_hd__or4_1
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1099 _6743_/Q VGND VGND VPWR VPWR _4297_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_206 _5994_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_217 input58/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_228 wire412/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_239 hold36/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5370_ _5574_/A0 _5370_/A1 _5375_/S VGND VGND VPWR VPWR _5370_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4321_ _4321_/A0 _6395_/A0 _4323_/S VGND VGND VPWR VPWR _4321_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7040_ _7102_/CLK _7040_/D fanout503/X VGND VGND VPWR VPWR _7040_/Q sky130_fd_sc_hd__dfrtp_2
X_4252_ _4252_/A _4330_/B VGND VGND VPWR VPWR _4257_/S sky130_fd_sc_hd__and2_2
XFILLER_113_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3203_ _6501_/Q VGND VGND VPWR VPWR _3203_/Y sky130_fd_sc_hd__inv_2
X_4183_ _4183_/A0 _3660_/X _4188_/S VGND VGND VPWR VPWR _6641_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6824_ _6825_/CLK _6824_/D fanout491/X VGND VGND VPWR VPWR _6824_/Q sky130_fd_sc_hd__dfrtp_1
X_6755_ _6755_/CLK _6755_/D fanout497/X VGND VGND VPWR VPWR _6755_/Q sky130_fd_sc_hd__dfrtp_1
X_3967_ input58/X hold564/X _3967_/S VGND VGND VPWR VPWR _3967_/X sky130_fd_sc_hd__mux2_8
X_5706_ _7152_/Q _5706_/B _5706_/C VGND VGND VPWR VPWR _5706_/X sky130_fd_sc_hd__and3_4
XFILLER_148_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6686_ _7094_/CLK _6686_/D fanout494/X VGND VGND VPWR VPWR _6686_/Q sky130_fd_sc_hd__dfrtp_2
X_3898_ _7144_/Q _7145_/Q VGND VGND VPWR VPWR _3899_/B sky130_fd_sc_hd__nor2_1
XFILLER_109_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5637_ _7157_/Q _5637_/B _6039_/A VGND VGND VPWR VPWR _5643_/B sky130_fd_sc_hd__and3_1
XFILLER_148_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5568_ _5586_/A0 hold987/X _5570_/S VGND VGND VPWR VPWR _5568_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold130 _4091_/X VGND VGND VPWR VPWR _6567_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_191_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold141 _3989_/X VGND VGND VPWR VPWR _6487_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_163_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4519_ _4871_/A _4994_/A _4515_/X _4850_/A _4518_/Y VGND VGND VPWR VPWR _4519_/X
+ sky130_fd_sc_hd__o2111a_1
Xhold152 _6838_/Q VGND VGND VPWR VPWR hold152/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold163 _6749_/Q VGND VGND VPWR VPWR hold163/X sky130_fd_sc_hd__dlygate4sd3_1
X_5499_ _5586_/A0 _5499_/A1 _5501_/S VGND VGND VPWR VPWR _5499_/X sky130_fd_sc_hd__mux2_1
Xhold174 _4110_/X VGND VGND VPWR VPWR _6579_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold185 _6729_/Q VGND VGND VPWR VPWR hold185/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 _5344_/X VGND VGND VPWR VPWR _6925_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7169_ _7182_/CLK _7169_/D fanout498/X VGND VGND VPWR VPWR _7169_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_58_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4870_ _4931_/B _4870_/B VGND VGND VPWR VPWR _4872_/B sky130_fd_sc_hd__nor2_1
XTAP_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3821_ hold17/A _3248_/Y _3821_/S VGND VGND VPWR VPWR _3821_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6540_ _7093_/CLK _6540_/D _6432_/A VGND VGND VPWR VPWR _6540_/Q sky130_fd_sc_hd__dfrtp_2
X_3752_ _6655_/Q _4198_/A _3733_/X VGND VGND VPWR VPWR _3755_/B sky130_fd_sc_hd__a21o_1
XFILLER_146_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6471_ _3945_/A1 _6471_/D _6426_/X VGND VGND VPWR VPWR _6471_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_185_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3683_ _6635_/Q _4174_/A _5187_/A _6794_/Q _3682_/X VGND VGND VPWR VPWR _3688_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5422_ _5536_/A1 _5422_/A1 _5429_/S VGND VGND VPWR VPWR _5422_/X sky130_fd_sc_hd__mux2_1
Xoutput202 _3200_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[34] sky130_fd_sc_hd__buf_12
Xoutput213 _3933_/X VGND VGND VPWR VPWR mgmt_gpio_out[0] sky130_fd_sc_hd__buf_12
Xoutput224 _3932_/X VGND VGND VPWR VPWR mgmt_gpio_out[1] sky130_fd_sc_hd__buf_12
Xoutput235 _6556_/Q VGND VGND VPWR VPWR mgmt_gpio_out[2] sky130_fd_sc_hd__buf_12
X_5353_ _5557_/A0 hold709/X _5357_/S VGND VGND VPWR VPWR _5353_/X sky130_fd_sc_hd__mux2_1
Xoutput246 _6559_/Q VGND VGND VPWR VPWR mgmt_gpio_out[5] sky130_fd_sc_hd__buf_12
Xoutput257 _3948_/Y VGND VGND VPWR VPWR pad_flash_io0_oeb sky130_fd_sc_hd__buf_12
XFILLER_160_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput268 _6795_/Q VGND VGND VPWR VPWR pll_div[2] sky130_fd_sc_hd__buf_12
X_4304_ hold36/X hold163/X _4305_/S VGND VGND VPWR VPWR _4304_/X sky130_fd_sc_hd__mux2_1
Xoutput279 _6487_/Q VGND VGND VPWR VPWR pll_trim[13] sky130_fd_sc_hd__buf_12
X_5284_ _5569_/A0 hold223/X _5285_/S VGND VGND VPWR VPWR _5284_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7023_ _7080_/CLK _7023_/D fanout502/X VGND VGND VPWR VPWR _7023_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_99_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4235_ _5521_/A0 hold964/X hold59/X VGND VGND VPWR VPWR _4235_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4166_ _4166_/A0 _3790_/X _4173_/S VGND VGND VPWR VPWR _6626_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4097_ hold379/X _4096_/X _4103_/S VGND VGND VPWR VPWR _4097_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6807_ _7102_/CLK _6807_/D fanout503/X VGND VGND VPWR VPWR _6807_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_168_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4999_ _4999_/A _4999_/B VGND VGND VPWR VPWR _4999_/Y sky130_fd_sc_hd__nand2_1
XFILLER_139_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6738_ _6740_/CLK _6738_/D fanout510/X VGND VGND VPWR VPWR _6738_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_23_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6669_ _6709_/CLK _6669_/D fanout494/X VGND VGND VPWR VPWR _6669_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_109_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout440 _5550_/A0 VGND VGND VPWR VPWR _5586_/A0 sky130_fd_sc_hd__buf_4
XFILLER_48_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout451 hold35/X VGND VGND VPWR VPWR _5539_/A1 sky130_fd_sc_hd__buf_8
XFILLER_120_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout462 _5555_/A0 VGND VGND VPWR VPWR _5531_/A1 sky130_fd_sc_hd__buf_6
XFILLER_171_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout473 _3195_/Y VGND VGND VPWR VPWR _6318_/S sky130_fd_sc_hd__buf_12
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout484 _3946_/B VGND VGND VPWR VPWR fanout484/X sky130_fd_sc_hd__buf_6
XFILLER_59_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout495 fanout496/X VGND VGND VPWR VPWR _6441_/A sky130_fd_sc_hd__buf_4
XFILLER_58_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4020_ _6396_/A0 hold617/X _4021_/S VGND VGND VPWR VPWR _4020_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5971_ _7154_/Q _7153_/Q VGND VGND VPWR VPWR _6039_/C sky130_fd_sc_hd__nor2_2
XFILLER_64_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4922_ _5177_/A _4922_/B _5177_/B _4920_/X VGND VGND VPWR VPWR _4923_/D sky130_fd_sc_hd__or4b_1
XFILLER_45_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4853_ _4683_/A _4707_/B _4447_/Y VGND VGND VPWR VPWR _4860_/C sky130_fd_sc_hd__o21a_1
XFILLER_193_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3804_ _6455_/Q _6454_/Q _6453_/Q VGND VGND VPWR VPWR _3890_/B sky130_fd_sc_hd__or3b_1
X_4784_ _4784_/A _4784_/B VGND VGND VPWR VPWR _5015_/B sky130_fd_sc_hd__nor2_1
XFILLER_119_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_opt_2_0_csclk _6820_/CLK VGND VGND VPWR VPWR clkbuf_opt_2_0_csclk/X sky130_fd_sc_hd__clkbuf_16
X_6523_ _6707_/CLK _6523_/D _6433_/A VGND VGND VPWR VPWR _6523_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_20_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3735_ _6482_/Q _3983_/A _3730_/X _5210_/A VGND VGND VPWR VPWR _3735_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6454_ _3945_/A1 _6454_/D _6409_/X VGND VGND VPWR VPWR _6454_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3666_ _6947_/Q _5367_/A _5358_/A _6939_/Q _3665_/X VGND VGND VPWR VPWR _3669_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_106_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5405_ _5459_/A0 hold335/X _5411_/S VGND VGND VPWR VPWR _5405_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6385_ _6698_/Q _6385_/A2 _6385_/B1 _6390_/A2 _6384_/X VGND VGND VPWR VPWR _6385_/X
+ sky130_fd_sc_hd__a221o_1
X_3597_ _7130_/Q _5571_/A _4204_/A _6663_/Q VGND VGND VPWR VPWR _3597_/X sky130_fd_sc_hd__a22o_1
XFILLER_133_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5336_ _5567_/A0 hold641/X _5339_/S VGND VGND VPWR VPWR _5336_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5267_ _5579_/A0 hold510/X _5267_/S VGND VGND VPWR VPWR _5267_/X sky130_fd_sc_hd__mux2_1
X_7006_ _7107_/CLK _7006_/D fanout514/X VGND VGND VPWR VPWR _7006_/Q sky130_fd_sc_hd__dfrtp_1
X_4218_ _5531_/A1 hold894/X _4221_/S VGND VGND VPWR VPWR _4218_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5198_ _6397_/A0 hold552/X _5199_/S VGND VGND VPWR VPWR _5198_/X sky130_fd_sc_hd__mux2_1
X_4149_ _6394_/A0 _4149_/A1 _4152_/S VGND VGND VPWR VPWR _4149_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3520_ _6730_/Q _4276_/A _4141_/A _6610_/Q VGND VGND VPWR VPWR _3524_/B sky130_fd_sc_hd__a22o_1
Xmax_cap404 _6040_/X VGND VGND VPWR VPWR _6212_/B1 sky130_fd_sc_hd__buf_8
XFILLER_6_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap415 _5992_/X VGND VGND VPWR VPWR _6024_/B sky130_fd_sc_hd__buf_12
Xhold707 _7014_/Q VGND VGND VPWR VPWR hold707/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold718 _4152_/X VGND VGND VPWR VPWR _6615_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold729 _7102_/Q VGND VGND VPWR VPWR hold729/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3451_ hold21/X _3729_/B VGND VGND VPWR VPWR _4174_/A sky130_fd_sc_hd__nor2_8
XFILLER_143_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3382_ _6480_/Q _3966_/A _5484_/A _7056_/Q VGND VGND VPWR VPWR _3382_/X sky130_fd_sc_hd__a22o_1
X_6170_ _6563_/Q _7179_/Q _6169_/X VGND VGND VPWR VPWR _6170_/X sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_3_csclk _7018_/CLK VGND VGND VPWR VPWR _6708_/CLK sky130_fd_sc_hd__clkbuf_16
X_5121_ _5140_/B _5121_/B VGND VGND VPWR VPWR _5139_/B sky130_fd_sc_hd__and2b_1
XFILLER_69_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1407 _6652_/Q VGND VGND VPWR VPWR hold1407/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1418 _6651_/Q VGND VGND VPWR VPWR _4194_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5052_ _4461_/B _5021_/B _4653_/C _4704_/B VGND VGND VPWR VPWR _5052_/X sky130_fd_sc_hd__o22a_1
Xhold1429 _7190_/Q VGND VGND VPWR VPWR _6350_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4003_ _5573_/A0 hold898/X _4009_/S VGND VGND VPWR VPWR _4003_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5954_ _6735_/Q _5697_/X _5953_/X VGND VGND VPWR VPWR _5957_/C sky130_fd_sc_hd__a21o_1
XFILLER_80_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4905_ _4905_/A _4905_/B VGND VGND VPWR VPWR _4925_/B sky130_fd_sc_hd__nand2_1
XFILLER_21_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5885_ _6532_/Q _5678_/X _5682_/X _6512_/Q VGND VGND VPWR VPWR _5885_/X sky130_fd_sc_hd__a22o_1
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4836_ _4836_/A _5001_/B VGND VGND VPWR VPWR _4836_/Y sky130_fd_sc_hd__nand2_1
XFILLER_178_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4767_ _4993_/A _4454_/Y _5049_/B _4983_/B _4766_/X VGND VGND VPWR VPWR _4767_/X
+ sky130_fd_sc_hd__a2111o_1
X_6506_ _6664_/CLK _6506_/D _6426_/A VGND VGND VPWR VPWR _6506_/Q sky130_fd_sc_hd__dfrtp_2
X_3718_ _7120_/Q _5562_/A _4104_/A input62/X _3717_/X VGND VGND VPWR VPWR _3721_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4698_ _4669_/X _4698_/B _4698_/C _4698_/D VGND VGND VPWR VPWR _4699_/D sky130_fd_sc_hd__and4b_1
XFILLER_106_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6437_ _6441_/A _6440_/B VGND VGND VPWR VPWR _6437_/X sky130_fd_sc_hd__and2_1
X_3649_ _6500_/Q _3778_/A2 _3547_/Y input97/X VGND VGND VPWR VPWR _3649_/X sky130_fd_sc_hd__a22o_1
XFILLER_136_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6368_ _6367_/X hold7/A _6386_/S VGND VGND VPWR VPWR _7198_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5319_ _5586_/A0 _5319_/A1 hold23/X VGND VGND VPWR VPWR _5319_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6299_ _6514_/Q _5977_/X _6323_/B1 _6739_/Q VGND VGND VPWR VPWR _6299_/X sky130_fd_sc_hd__a22o_1
Xhold12 hold12/A VGND VGND VPWR VPWR hold12/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold23 hold23/A VGND VGND VPWR VPWR hold23/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold34 hold34/A VGND VGND VPWR VPWR hold34/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 hold45/A VGND VGND VPWR VPWR hold45/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 hold56/A VGND VGND VPWR VPWR hold56/X sky130_fd_sc_hd__buf_6
Xhold67 hold67/A VGND VGND VPWR VPWR hold67/X sky130_fd_sc_hd__buf_6
Xhold78 hold78/A VGND VGND VPWR VPWR hold78/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold89 hold89/A VGND VGND VPWR VPWR hold89/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_9 _5466_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5670_ _5938_/B _5706_/B _5699_/C VGND VGND VPWR VPWR _5670_/X sky130_fd_sc_hd__and3_4
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4621_ _4793_/A _4621_/B _4621_/C VGND VGND VPWR VPWR _4639_/B sky130_fd_sc_hd__or3_4
XFILLER_175_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4552_ _4553_/B _4552_/B VGND VGND VPWR VPWR _4792_/B sky130_fd_sc_hd__nor2_1
XFILLER_116_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold504 _6937_/Q VGND VGND VPWR VPWR hold504/X sky130_fd_sc_hd__dlygate4sd3_1
X_3503_ _3528_/A _4111_/B VGND VGND VPWR VPWR _4198_/A sky130_fd_sc_hd__nor2_4
Xhold515 _5375_/X VGND VGND VPWR VPWR _6953_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold526 _6493_/Q VGND VGND VPWR VPWR hold526/X sky130_fd_sc_hd__dlygate4sd3_1
X_4483_ _4483_/A VGND VGND VPWR VPWR _5106_/A sky130_fd_sc_hd__inv_2
Xhold537 _5321_/X VGND VGND VPWR VPWR _6905_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 _6744_/Q VGND VGND VPWR VPWR hold548/X sky130_fd_sc_hd__dlygate4sd3_1
X_6222_ _6531_/Q _6272_/B VGND VGND VPWR VPWR _6222_/X sky130_fd_sc_hd__and2_1
XFILLER_131_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold559 _4158_/X VGND VGND VPWR VPWR _6620_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3434_ _7087_/Q _5520_/A _5349_/A _6935_/Q VGND VGND VPWR VPWR _3434_/X sky130_fd_sc_hd__a22o_1
XFILLER_171_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6153_ _6991_/Q _6203_/A2 _6024_/C _6911_/Q _6152_/X VGND VGND VPWR VPWR _6156_/C
+ sky130_fd_sc_hd__a221o_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3365_ _6953_/Q _5367_/A _5340_/A _6929_/Q VGND VGND VPWR VPWR _3365_/X sky130_fd_sc_hd__a22o_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5104_ _5104_/A _5104_/B _5104_/C _5104_/D VGND VGND VPWR VPWR _6779_/D sky130_fd_sc_hd__or4_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1204 _4212_/X VGND VGND VPWR VPWR _6666_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6084_ _6084_/A _6084_/B _6084_/C _6084_/D VGND VGND VPWR VPWR _6085_/B sky130_fd_sc_hd__or4_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3296_ _5212_/B _3495_/A VGND VGND VPWR VPWR _5520_/A sky130_fd_sc_hd__nor2_8
Xhold1215 hold1446/X VGND VGND VPWR VPWR _5359_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1226 _6566_/Q VGND VGND VPWR VPWR _4089_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1237 _4331_/X VGND VGND VPWR VPWR _6771_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1248 _6986_/Q VGND VGND VPWR VPWR _5413_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5035_ _5035_/A _5035_/B VGND VGND VPWR VPWR _5035_/Y sky130_fd_sc_hd__nand2_1
Xhold1259 _7018_/Q VGND VGND VPWR VPWR _5449_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6986_ _6986_/CLK _6986_/D fanout491/X VGND VGND VPWR VPWR _6986_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_25_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5937_ _6637_/Q _5655_/X _5693_/X _6658_/Q _5936_/X VGND VGND VPWR VPWR _5945_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_40_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5868_ _6675_/Q _5670_/X _5676_/X _6526_/Q _5867_/X VGND VGND VPWR VPWR _5869_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_179_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4819_ _4595_/B _4981_/C _4819_/C _4971_/B VGND VGND VPWR VPWR _4821_/C sky130_fd_sc_hd__and4bb_1
XFILLER_166_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5799_ _7007_/Q _5664_/X _5682_/X _7087_/Q _5798_/X VGND VGND VPWR VPWR _5799_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_119_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput102 wb_adr_i[12] VGND VGND VPWR VPWR _4338_/B sky130_fd_sc_hd__clkbuf_1
Xinput113 wb_adr_i[22] VGND VGND VPWR VPWR _4390_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_130_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput124 wb_adr_i[3] VGND VGND VPWR VPWR _4846_/B sky130_fd_sc_hd__clkbuf_16
Xinput135 wb_dat_i[12] VGND VGND VPWR VPWR _6376_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_193_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput146 wb_dat_i[22] VGND VGND VPWR VPWR _6382_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput157 wb_dat_i[3] VGND VGND VPWR VPWR _6373_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput168 wb_sel_i[3] VGND VGND VPWR VPWR _6357_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_76_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_560 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6840_ _7126_/CLK _6840_/D fanout524/X VGND VGND VPWR VPWR _6840_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_63_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6771_ _6825_/CLK _6771_/D fanout491/X VGND VGND VPWR VPWR _6771_/Q sky130_fd_sc_hd__dfrtp_2
X_3983_ _3983_/A _6392_/B VGND VGND VPWR VPWR _3991_/S sky130_fd_sc_hd__and2_2
XFILLER_22_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5722_ _7043_/Q _5848_/B1 _5691_/B _6971_/Q _5690_/X VGND VGND VPWR VPWR _5722_/X
+ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_21_csclk _6820_/CLK VGND VGND VPWR VPWR _7043_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_31_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5653_ _7151_/Q _7150_/Q VGND VGND VPWR VPWR _5700_/C sky130_fd_sc_hd__and2b_2
XFILLER_176_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4604_ _4621_/B _4971_/B _4793_/A VGND VGND VPWR VPWR _4606_/B sky130_fd_sc_hd__a21o_1
X_5584_ _5584_/A0 hold447/X hold70/X VGND VGND VPWR VPWR _5584_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_36_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7140_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_163_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold301 hold301/A VGND VGND VPWR VPWR hold301/X sky130_fd_sc_hd__dlygate4sd3_1
X_4535_ _4745_/A _4802_/A VGND VGND VPWR VPWR _4824_/A sky130_fd_sc_hd__or2_1
Xhold312 _5401_/X VGND VGND VPWR VPWR _6976_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 _7137_/Q VGND VGND VPWR VPWR hold323/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 _4161_/X VGND VGND VPWR VPWR _6622_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold345 _6891_/Q VGND VGND VPWR VPWR hold345/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold356 _5220_/X VGND VGND VPWR VPWR _6818_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4466_ _4846_/C _4466_/B VGND VGND VPWR VPWR _4832_/B sky130_fd_sc_hd__nand2_8
Xhold367 _6617_/Q VGND VGND VPWR VPWR hold367/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 _4239_/X VGND VGND VPWR VPWR _6685_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6205_ _6961_/Q _6336_/A2 _6205_/B1 _7065_/Q VGND VGND VPWR VPWR _6205_/X sky130_fd_sc_hd__a22o_1
XFILLER_171_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold389 _7017_/Q VGND VGND VPWR VPWR hold389/X sky130_fd_sc_hd__dlygate4sd3_1
X_3417_ _3714_/B _3525_/B VGND VGND VPWR VPWR _5193_/A sky130_fd_sc_hd__nor2_8
X_7185_ _7187_/CLK _7185_/D fanout490/X VGND VGND VPWR VPWR _7185_/Q sky130_fd_sc_hd__dfrtp_1
X_4397_ _4931_/A _4732_/A VGND VGND VPWR VPWR _4484_/A sky130_fd_sc_hd__nand2_1
XFILLER_131_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6136_ _6918_/Q wire412/X _6024_/D _6942_/Q VGND VGND VPWR VPWR _6136_/X sky130_fd_sc_hd__a22o_1
X_3348_ _6993_/Q _5412_/A _5484_/A _7057_/Q _3347_/X VGND VGND VPWR VPWR _3355_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1001 _6967_/Q VGND VGND VPWR VPWR _5391_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_133_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1012 _5400_/X VGND VGND VPWR VPWR _6975_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1023 _7055_/Q VGND VGND VPWR VPWR _5490_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_6067_ _6867_/Q _6199_/B1 _6025_/D _6963_/Q _6066_/X VGND VGND VPWR VPWR _6068_/D
+ sky130_fd_sc_hd__a221o_1
Xhold1034 _5563_/X VGND VGND VPWR VPWR _7119_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3279_ hold48/X hold19/X VGND VGND VPWR VPWR hold20/A sky130_fd_sc_hd__or2_2
Xhold1045 _6940_/Q VGND VGND VPWR VPWR _5361_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1056 _5298_/X VGND VGND VPWR VPWR _6884_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1067 _6791_/Q VGND VGND VPWR VPWR _5185_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5018_ _5018_/A _5023_/C _5018_/C VGND VGND VPWR VPWR _5106_/B sky130_fd_sc_hd__nor3_1
Xhold1078 _5230_/X VGND VGND VPWR VPWR _6824_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1089 _4047_/X VGND VGND VPWR VPWR _6536_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_207 _6027_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_218 _6803_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_229 _5569_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6969_ _6969_/CLK _6969_/D fanout506/X VGND VGND VPWR VPWR _6969_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_186_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold890 _7056_/Q VGND VGND VPWR VPWR hold890/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_95_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1590 _7169_/Q VGND VGND VPWR VPWR _5860_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4320_ _4320_/A0 _6394_/A0 _4323_/S VGND VGND VPWR VPWR _4320_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4251_ _5534_/A1 hold777/X _4251_/S VGND VGND VPWR VPWR _4251_/X sky130_fd_sc_hd__mux2_1
X_3202_ _7098_/Q VGND VGND VPWR VPWR _3202_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4182_ _4182_/A0 _3723_/X _4188_/S VGND VGND VPWR VPWR _6640_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6823_ _7138_/CLK _6823_/D fanout520/X VGND VGND VPWR VPWR _6823_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_168_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6754_ _6755_/CLK _6754_/D fanout497/X VGND VGND VPWR VPWR _6754_/Q sky130_fd_sc_hd__dfrtp_1
X_3966_ _3966_/A _5535_/B VGND VGND VPWR VPWR _3982_/S sky130_fd_sc_hd__and2_2
X_5705_ _5938_/B _5705_/B _5706_/C VGND VGND VPWR VPWR _5705_/X sky130_fd_sc_hd__and3_4
X_6685_ _6709_/CLK _6685_/D fanout511/X VGND VGND VPWR VPWR _6685_/Q sky130_fd_sc_hd__dfrtp_2
X_3897_ _5615_/A _6819_/Q _3896_/X VGND VGND VPWR VPWR _6562_/D sky130_fd_sc_hd__o21ai_1
XFILLER_176_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5636_ _5636_/A1 _5624_/B _5634_/Y _5635_/X VGND VGND VPWR VPWR _7156_/D sky130_fd_sc_hd__a31o_1
XFILLER_164_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_530 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5567_ _5567_/A0 hold655/X _5570_/S VGND VGND VPWR VPWR _5567_/X sky130_fd_sc_hd__mux2_1
Xhold120 _5456_/X VGND VGND VPWR VPWR _7025_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4518_ _5124_/A VGND VGND VPWR VPWR _4518_/Y sky130_fd_sc_hd__inv_2
Xhold131 _7202_/Q VGND VGND VPWR VPWR hold131/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold142 _7078_/Q VGND VGND VPWR VPWR hold142/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 _5246_/X VGND VGND VPWR VPWR _6838_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5498_ hold85/X hold121/X _5501_/S VGND VGND VPWR VPWR _5498_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold164 _4304_/X VGND VGND VPWR VPWR _6749_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 _6803_/Q VGND VGND VPWR VPWR hold175/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold186 _4280_/X VGND VGND VPWR VPWR _6729_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4449_ _4932_/A _4742_/A _4836_/A VGND VGND VPWR VPWR _4502_/A sky130_fd_sc_hd__and3b_1
XFILLER_104_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold197 _6837_/Q VGND VGND VPWR VPWR hold197/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7168_ _7182_/CLK _7168_/D fanout502/X VGND VGND VPWR VPWR _7168_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_58_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6119_ _6168_/A _6119_/B _6119_/C _6119_/D VGND VGND VPWR VPWR _6119_/X sky130_fd_sc_hd__or4_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7099_ _7115_/CLK _7099_/D fanout501/X VGND VGND VPWR VPWR _7099_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3820_ hold72/A _3823_/B VGND VGND VPWR VPWR _3820_/Y sky130_fd_sc_hd__nor2_1
XFILLER_177_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3751_ input71/X _3751_/A2 _4085_/S _3959_/A _3750_/X VGND VGND VPWR VPWR _3755_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_32_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6470_ _3945_/A1 _6470_/D _6425_/X VGND VGND VPWR VPWR hold91/A sky130_fd_sc_hd__dfrtp_1
XFILLER_146_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3682_ input12/X _3268_/Y _3340_/Y input21/X VGND VGND VPWR VPWR _3682_/X sky130_fd_sc_hd__a22o_2
XFILLER_145_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5421_ _5421_/A _5535_/B VGND VGND VPWR VPWR _5429_/S sky130_fd_sc_hd__nand2_8
XFILLER_173_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput203 _3922_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[35] sky130_fd_sc_hd__buf_12
XFILLER_126_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput214 _3926_/X VGND VGND VPWR VPWR mgmt_gpio_out[10] sky130_fd_sc_hd__buf_12
X_5352_ _5574_/A0 _5352_/A1 _5357_/S VGND VGND VPWR VPWR _5352_/X sky130_fd_sc_hd__mux2_1
Xoutput225 _6550_/Q VGND VGND VPWR VPWR mgmt_gpio_out[20] sky130_fd_sc_hd__buf_12
Xoutput236 _6832_/Q VGND VGND VPWR VPWR mgmt_gpio_out[30] sky130_fd_sc_hd__buf_12
Xoutput247 _3929_/X VGND VGND VPWR VPWR mgmt_gpio_out[6] sky130_fd_sc_hd__buf_12
XFILLER_114_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput258 _7213_/X VGND VGND VPWR VPWR pad_flash_io1_do sky130_fd_sc_hd__buf_12
X_4303_ hold44/X hold225/X _4305_/S VGND VGND VPWR VPWR _4303_/X sky130_fd_sc_hd__mux2_1
Xoutput269 _6796_/Q VGND VGND VPWR VPWR pll_div[3] sky130_fd_sc_hd__buf_12
X_5283_ _5586_/A0 _5283_/A1 _5285_/S VGND VGND VPWR VPWR _5283_/X sky130_fd_sc_hd__mux2_1
X_7022_ _7082_/CLK _7022_/D fanout518/X VGND VGND VPWR VPWR _7022_/Q sky130_fd_sc_hd__dfrtp_4
X_4234_ hold58/X _5580_/B VGND VGND VPWR VPWR hold59/A sky130_fd_sc_hd__nand2_2
XFILLER_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4165_ _6695_/Q _6348_/B VGND VGND VPWR VPWR _4173_/S sky130_fd_sc_hd__and2_4
XFILLER_114_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4096_ hold152/X hold85/X _4102_/S VGND VGND VPWR VPWR _4096_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6806_ _7074_/CLK _6806_/D fanout501/X VGND VGND VPWR VPWR _6806_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_168_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4998_ _4999_/A _4657_/C _4741_/C _4770_/C _4894_/C VGND VGND VPWR VPWR _5045_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_11_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3949_ _6459_/Q _3949_/B VGND VGND VPWR VPWR _3950_/A sky130_fd_sc_hd__or2_1
X_6737_ _6740_/CLK _6737_/D fanout510/X VGND VGND VPWR VPWR _6737_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6668_ _6709_/CLK _6668_/D fanout494/X VGND VGND VPWR VPWR _6668_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_139_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5619_ _5622_/B VGND VGND VPWR VPWR _5619_/Y sky130_fd_sc_hd__inv_2
X_6599_ _6759_/CLK _6599_/D fanout489/X VGND VGND VPWR VPWR _6599_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_192_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout441 hold127/X VGND VGND VPWR VPWR _5550_/A0 sky130_fd_sc_hd__buf_6
Xfanout452 hold36/X VGND VGND VPWR VPWR _5584_/A0 sky130_fd_sc_hd__buf_6
XFILLER_59_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout463 hold9/X VGND VGND VPWR VPWR _5555_/A0 sky130_fd_sc_hd__buf_6
XFILLER_120_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout474 _3981_/S VGND VGND VPWR VPWR _3971_/S sky130_fd_sc_hd__buf_12
XFILLER_171_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout485 _3946_/B VGND VGND VPWR VPWR fanout485/X sky130_fd_sc_hd__buf_4
Xfanout496 fanout497/X VGND VGND VPWR VPWR fanout496/X sky130_fd_sc_hd__buf_6
XFILLER_59_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5970_ _5970_/A0 _5969_/X _6171_/S VGND VGND VPWR VPWR _7174_/D sky130_fd_sc_hd__mux2_1
XFILLER_18_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4921_ _4674_/A _4684_/A _4622_/Y _4635_/Y VGND VGND VPWR VPWR _4922_/B sky130_fd_sc_hd__a31o_1
XFILLER_52_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4852_ _4674_/A _4684_/A _4595_/B _4506_/Y VGND VGND VPWR VPWR _4862_/B sky130_fd_sc_hd__a31o_1
XFILLER_178_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3803_ _6471_/Q _3838_/B VGND VGND VPWR VPWR _3890_/A sky130_fd_sc_hd__nand2_1
XFILLER_21_748 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4783_ _4783_/A _4802_/D VGND VGND VPWR VPWR _4783_/Y sky130_fd_sc_hd__nor2_1
X_6522_ _6707_/CLK _6522_/D _6433_/A VGND VGND VPWR VPWR _6522_/Q sky130_fd_sc_hd__dfrtp_2
X_3734_ _7026_/Q _5457_/A _5203_/A _6806_/Q VGND VGND VPWR VPWR _3734_/X sky130_fd_sc_hd__a22o_1
XFILLER_186_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6453_ _3945_/A1 _6453_/D _6408_/X VGND VGND VPWR VPWR _6453_/Q sky130_fd_sc_hd__dfrtp_1
X_3665_ _6767_/Q _4324_/A _4330_/A _6772_/Q VGND VGND VPWR VPWR _3665_/X sky130_fd_sc_hd__a22o_2
XFILLER_174_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5404_ _5581_/A0 _5404_/A1 _5411_/S VGND VGND VPWR VPWR _5404_/X sky130_fd_sc_hd__mux2_1
X_6384_ _6700_/Q _6384_/A2 _6384_/B1 _6699_/Q VGND VGND VPWR VPWR _6384_/X sky130_fd_sc_hd__a22o_1
X_3596_ _7013_/Q _5439_/A _4010_/A _6509_/Q _3557_/X VGND VGND VPWR VPWR _3600_/C
+ sky130_fd_sc_hd__a221o_1
X_5335_ _5557_/A0 hold605/X _5339_/S VGND VGND VPWR VPWR _5335_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5266_ _5578_/A0 hold823/X _5267_/S VGND VGND VPWR VPWR _5266_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7005_ _7075_/CLK _7005_/D fanout526/X VGND VGND VPWR VPWR _7005_/Q sky130_fd_sc_hd__dfrtp_4
X_4217_ _5521_/A0 hold954/X _4221_/S VGND VGND VPWR VPWR _4217_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5197_ _6396_/A0 hold593/X _5199_/S VGND VGND VPWR VPWR _5197_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4148_ _5212_/C _4148_/A1 _4152_/S VGND VGND VPWR VPWR _4148_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4079_ hold209/X _5558_/A0 _4085_/S VGND VGND VPWR VPWR _4079_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_82 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap405 _6036_/X VGND VGND VPWR VPWR _6329_/B1 sky130_fd_sc_hd__buf_12
XFILLER_128_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap416 _6029_/B VGND VGND VPWR VPWR _6338_/B1 sky130_fd_sc_hd__buf_8
XFILLER_116_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold708 _5444_/X VGND VGND VPWR VPWR _7014_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold719 _6754_/Q VGND VGND VPWR VPWR hold719/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_183_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3450_ _3495_/A _4111_/B VGND VGND VPWR VPWR _5529_/A sky130_fd_sc_hd__nor2_4
XFILLER_170_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3381_ _6976_/Q _5394_/A hold31/A _6880_/Q VGND VGND VPWR VPWR _3381_/X sky130_fd_sc_hd__a22o_1
XFILLER_97_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5120_ _5171_/A _5172_/A _5119_/Y VGND VGND VPWR VPWR _5121_/B sky130_fd_sc_hd__or3b_1
XFILLER_124_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5051_ _5044_/X _5048_/X _5050_/X VGND VGND VPWR VPWR _5104_/A sky130_fd_sc_hd__o21a_1
Xhold1408 _6653_/Q VGND VGND VPWR VPWR hold1408/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1419 _6648_/Q VGND VGND VPWR VPWR _4191_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4002_ _5536_/A1 _4002_/A1 _4009_/S VGND VGND VPWR VPWR _4002_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5953_ _6638_/Q _5655_/X _5659_/X _6705_/Q VGND VGND VPWR VPWR _5953_/X sky130_fd_sc_hd__a22o_1
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4904_ _4639_/A _4675_/A _4902_/X _4693_/A _4903_/X VGND VGND VPWR VPWR _4905_/B
+ sky130_fd_sc_hd__o221a_1
X_5884_ _6707_/Q _5675_/X _5683_/X _6612_/Q _5883_/X VGND VGND VPWR VPWR _5891_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_33_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4835_ _4932_/A _4835_/B VGND VGND VPWR VPWR _4857_/A sky130_fd_sc_hd__or2_1
XFILLER_178_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4766_ _4993_/A _4516_/B _4815_/A _4987_/B _4765_/X VGND VGND VPWR VPWR _4766_/X
+ sky130_fd_sc_hd__a2111o_1
X_6505_ _7102_/CLK _6505_/D fanout502/X VGND VGND VPWR VPWR _6505_/Q sky130_fd_sc_hd__dfrtp_4
X_3717_ _6475_/Q _3966_/A _3983_/A _6483_/Q VGND VGND VPWR VPWR _3717_/X sky130_fd_sc_hd__a22o_4
XFILLER_162_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4697_ _4784_/A _4683_/B _4696_/X _4653_/X VGND VGND VPWR VPWR _4698_/D sky130_fd_sc_hd__o211a_1
XFILLER_20_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3648_ _7092_/Q _5529_/A _4129_/A _6598_/Q _3647_/X VGND VGND VPWR VPWR _3651_/C
+ sky130_fd_sc_hd__a221o_1
X_6436_ _6441_/A _6440_/B VGND VGND VPWR VPWR _6436_/X sky130_fd_sc_hd__and2_1
XFILLER_161_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6367_ _6698_/Q _6367_/A2 _6367_/B1 _6390_/A2 _6366_/X VGND VGND VPWR VPWR _6367_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_88_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3579_ input55/X _5232_/A _4258_/A _6714_/Q _3578_/X VGND VGND VPWR VPWR _3582_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_161_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5318_ _5567_/A0 hold769/X hold23/X VGND VGND VPWR VPWR _5318_/X sky130_fd_sc_hd__mux2_1
X_6298_ _7093_/Q _5642_/X _5992_/X _6678_/Q VGND VGND VPWR VPWR _6298_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_718 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold13 hold13/A VGND VGND VPWR VPWR hold13/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 hold24/A VGND VGND VPWR VPWR hold24/X sky130_fd_sc_hd__dlygate4sd3_1
X_5249_ hold40/X hold81/X hold14/X VGND VGND VPWR VPWR hold82/A sky130_fd_sc_hd__mux2_1
XFILLER_29_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold35 hold35/A VGND VGND VPWR VPWR hold35/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 hold46/A VGND VGND VPWR VPWR hold46/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold57 hold57/A VGND VGND VPWR VPWR hold57/X sky130_fd_sc_hd__clkbuf_8
XFILLER_75_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold68 hold68/A VGND VGND VPWR VPWR hold68/X sky130_fd_sc_hd__clkbuf_16
XFILLER_29_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold79 hold79/A VGND VGND VPWR VPWR hold79/X sky130_fd_sc_hd__clkbuf_16
XFILLER_90_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4620_ _5108_/A _5021_/B VGND VGND VPWR VPWR _5115_/B sky130_fd_sc_hd__nor2_1
XFILLER_175_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_764 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4551_ _4341_/X _4971_/B _4588_/A VGND VGND VPWR VPWR _4552_/B sky130_fd_sc_hd__a21oi_1
XFILLER_144_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3502_ hold57/X hold21/X VGND VGND VPWR VPWR _4153_/A sky130_fd_sc_hd__nor2_2
XFILLER_156_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold505 _5357_/X VGND VGND VPWR VPWR _6937_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold516 _6494_/Q VGND VGND VPWR VPWR hold516/X sky130_fd_sc_hd__dlygate4sd3_1
X_4482_ _4596_/A _5013_/A VGND VGND VPWR VPWR _4483_/A sky130_fd_sc_hd__or2_2
Xhold527 _3996_/X VGND VGND VPWR VPWR _6493_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_183_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold538 _6977_/Q VGND VGND VPWR VPWR hold538/X sky130_fd_sc_hd__dlygate4sd3_1
X_6221_ _6726_/Q _6320_/A2 _6320_/B1 _6616_/Q VGND VGND VPWR VPWR _6221_/X sky130_fd_sc_hd__a22o_2
XFILLER_171_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold549 _4298_/X VGND VGND VPWR VPWR _6744_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3433_ _6503_/Q _3778_/A2 _5403_/A _6983_/Q _3432_/X VGND VGND VPWR VPWR _3447_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_131_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6152_ _7023_/Q _6204_/A2 _6025_/B _7108_/Q VGND VGND VPWR VPWR _6152_/X sky130_fd_sc_hd__a22o_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3364_ _7025_/Q _5448_/A _5544_/A _7110_/Q _3363_/X VGND VGND VPWR VPWR _3372_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_106_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5103_ _5103_/A _5103_/B VGND VGND VPWR VPWR _5104_/D sky130_fd_sc_hd__nor2_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6083_ _6948_/Q _6024_/A _6322_/B1 _7113_/Q _6082_/X VGND VGND VPWR VPWR _6084_/D
+ sky130_fd_sc_hd__a221o_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3295_ _5212_/A hold29/A VGND VGND VPWR VPWR _3295_/Y sky130_fd_sc_hd__nor2_8
XFILLER_57_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1205 _6962_/Q VGND VGND VPWR VPWR _5386_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1216 _6798_/Q VGND VGND VPWR VPWR _5194_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ _4962_/Y _4991_/Y _5033_/X _4232_/X _5034_/B2 VGND VGND VPWR VPWR _6778_/D
+ sky130_fd_sc_hd__o32a_1
Xhold1227 _4089_/X VGND VGND VPWR VPWR _6566_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1238 _6820_/Q VGND VGND VPWR VPWR _5224_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1249 _5413_/X VGND VGND VPWR VPWR _6986_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_65_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6985_ _6992_/CLK _6985_/D fanout517/X VGND VGND VPWR VPWR _6985_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5936_ _6624_/Q _5661_/X _5676_/X _6529_/Q VGND VGND VPWR VPWR _5936_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5867_ _6706_/Q _5675_/X _5697_/X _6731_/Q VGND VGND VPWR VPWR _5867_/X sky130_fd_sc_hd__a22o_1
XFILLER_139_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4818_ _4818_/A _4818_/B _4618_/C VGND VGND VPWR VPWR _4821_/B sky130_fd_sc_hd__or3b_1
X_5798_ _7071_/Q _5678_/X _5686_/X _7015_/Q _5797_/X VGND VGND VPWR VPWR _5798_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_135_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4749_ _4638_/B _4971_/B _4797_/A VGND VGND VPWR VPWR _4965_/B sky130_fd_sc_hd__and3b_2
XFILLER_147_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6419_ _6441_/A _6440_/B VGND VGND VPWR VPWR _6419_/X sky130_fd_sc_hd__and2_1
XFILLER_162_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput103 wb_adr_i[13] VGND VGND VPWR VPWR _4338_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_76_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput114 wb_adr_i[23] VGND VGND VPWR VPWR _4390_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput125 wb_adr_i[4] VGND VGND VPWR VPWR _4621_/B sky130_fd_sc_hd__buf_6
XFILLER_130_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput136 wb_dat_i[13] VGND VGND VPWR VPWR _6379_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_103_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput147 wb_dat_i[23] VGND VGND VPWR VPWR _6385_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_102_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput158 wb_dat_i[4] VGND VGND VPWR VPWR _6375_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput169 wb_stb_i VGND VGND VPWR VPWR input169/X sky130_fd_sc_hd__clkbuf_4
XFILLER_186_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_2_csclk _7018_/CLK VGND VGND VPWR VPWR _6707_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6770_ _6825_/CLK _6770_/D fanout490/X VGND VGND VPWR VPWR _6770_/Q sky130_fd_sc_hd__dfrtp_2
X_3982_ hold725/X _5552_/A0 _3982_/S VGND VGND VPWR VPWR _3982_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5721_ _6907_/Q _5685_/X _5966_/B1 _7035_/Q _5720_/X VGND VGND VPWR VPWR _5728_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_175_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5652_ _6319_/S VGND VGND VPWR VPWR _5652_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4603_ _4745_/A _5023_/B VGND VGND VPWR VPWR _5059_/A sky130_fd_sc_hd__nor2_2
X_5583_ _5583_/A0 hold323/X hold70/X VGND VGND VPWR VPWR _5583_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4534_ _4745_/A _4802_/A VGND VGND VPWR VPWR _4964_/A sky130_fd_sc_hd__nor2_1
Xhold302 _4326_/X VGND VGND VPWR VPWR _6767_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold313 _7036_/Q VGND VGND VPWR VPWR hold313/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold324 _5583_/X VGND VGND VPWR VPWR _7137_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 _6979_/Q VGND VGND VPWR VPWR hold335/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 _5306_/X VGND VGND VPWR VPWR _6891_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4465_ _4846_/C _4466_/B VGND VGND VPWR VPWR _4684_/A sky130_fd_sc_hd__and2_4
Xhold357 _7003_/Q VGND VGND VPWR VPWR hold357/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold368 _4155_/X VGND VGND VPWR VPWR _6617_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6204_ _7025_/Q _6204_/A2 _6025_/B _7110_/Q _6203_/X VGND VGND VPWR VPWR _6204_/X
+ sky130_fd_sc_hd__a221o_1
X_3416_ hold56/X hold75/X VGND VGND VPWR VPWR _3525_/B sky130_fd_sc_hd__nand2_8
XFILLER_131_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold379 _6570_/Q VGND VGND VPWR VPWR hold379/X sky130_fd_sc_hd__dlygate4sd3_1
X_7184_ _7187_/CLK _7184_/D fanout490/X VGND VGND VPWR VPWR _7184_/Q sky130_fd_sc_hd__dfrtp_1
X_4396_ _4846_/A _4596_/A _5021_/A VGND VGND VPWR VPWR _4396_/X sky130_fd_sc_hd__or3_2
X_6135_ _7115_/Q _6025_/C _6030_/X _6998_/Q _6134_/X VGND VGND VPWR VPWR _6143_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3347_ input19/X _3268_/Y _5250_/A _6849_/Q VGND VGND VPWR VPWR _3347_/X sky130_fd_sc_hd__a22o_1
XFILLER_100_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1002 _5391_/X VGND VGND VPWR VPWR _6967_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1013 _6943_/Q VGND VGND VPWR VPWR _5364_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6066_ _7051_/Q _5988_/X _6022_/B _6899_/Q VGND VGND VPWR VPWR _6066_/X sky130_fd_sc_hd__a22o_1
Xhold1024 _5490_/X VGND VGND VPWR VPWR _7055_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1035 _7002_/Q VGND VGND VPWR VPWR _5431_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_3278_ _3546_/A _3526_/A VGND VGND VPWR VPWR _3278_/Y sky130_fd_sc_hd__nor2_8
Xhold1046 _5361_/X VGND VGND VPWR VPWR _6940_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5017_ _5017_/A _5017_/B VGND VGND VPWR VPWR _5083_/C sky130_fd_sc_hd__nor2_1
Xhold1057 _6821_/Q VGND VGND VPWR VPWR _5226_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1068 _5185_/X VGND VGND VPWR VPWR _6791_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1079 hold1544/X VGND VGND VPWR VPWR _5231_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_208 _6021_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_219 _6488_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6968_ _6969_/CLK _6968_/D fanout506/X VGND VGND VPWR VPWR _6968_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_13_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5919_ _6753_/Q _5664_/X _5670_/X _6677_/Q VGND VGND VPWR VPWR _5919_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6899_ _7139_/CLK hold24/X fanout518/X VGND VGND VPWR VPWR _6899_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_179_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold880 _7104_/Q VGND VGND VPWR VPWR hold880/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold891 _5491_/X VGND VGND VPWR VPWR _7056_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_67_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1580 _6562_/Q VGND VGND VPWR VPWR _3193_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1591 _6577_/Q VGND VGND VPWR VPWR hold699/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_724 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4250_ _5533_/A1 hold727/X _4251_/S VGND VGND VPWR VPWR _4250_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3201_ _7106_/Q VGND VGND VPWR VPWR _3201_/Y sky130_fd_sc_hd__inv_2
X_4181_ _4181_/A0 _3790_/X _4188_/S VGND VGND VPWR VPWR _6639_/D sky130_fd_sc_hd__mux2_1
XFILLER_121_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6822_ _7138_/CLK hold10/X fanout520/X VGND VGND VPWR VPWR _6822_/Q sky130_fd_sc_hd__dfrtp_4
X_6753_ _6753_/CLK _6753_/D fanout491/X VGND VGND VPWR VPWR _6753_/Q sky130_fd_sc_hd__dfstp_1
X_3965_ hold12/X _3971_/S hold111/X VGND VGND VPWR VPWR hold13/A sky130_fd_sc_hd__o21ai_4
X_5704_ _6978_/Q _5702_/X _5703_/X _6850_/Q VGND VGND VPWR VPWR _5704_/X sky130_fd_sc_hd__a22o_2
X_3896_ _5648_/C _3896_/B VGND VGND VPWR VPWR _3896_/X sky130_fd_sc_hd__or2_1
X_6684_ _6709_/CLK hold60/X _6441_/A VGND VGND VPWR VPWR _6684_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_148_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5635_ _6564_/Q _6000_/A _6033_/A VGND VGND VPWR VPWR _5635_/X sky130_fd_sc_hd__and3_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5566_ _5584_/A0 hold443/X _5570_/S VGND VGND VPWR VPWR _5566_/X sky130_fd_sc_hd__mux2_1
Xhold110 _7206_/Q VGND VGND VPWR VPWR hold110/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 _7062_/Q VGND VGND VPWR VPWR hold121/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_163_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4517_ _4942_/A _5002_/A VGND VGND VPWR VPWR _5124_/A sky130_fd_sc_hd__nor2_2
Xhold132 _3977_/X VGND VGND VPWR VPWR hold132/X sky130_fd_sc_hd__dlygate4sd3_1
X_5497_ _5584_/A0 hold435/X _5501_/S VGND VGND VPWR VPWR _5497_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold143 _5516_/X VGND VGND VPWR VPWR _7078_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 _6999_/Q VGND VGND VPWR VPWR hold154/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 _7139_/Q VGND VGND VPWR VPWR hold165/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 _5199_/X VGND VGND VPWR VPWR _6803_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4448_ _4742_/A _4448_/B VGND VGND VPWR VPWR _4510_/A sky130_fd_sc_hd__nand2_1
XFILLER_171_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold187 _6998_/Q VGND VGND VPWR VPWR hold187/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 _5245_/X VGND VGND VPWR VPWR _6837_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7167_ _7181_/CLK _7167_/D fanout502/X VGND VGND VPWR VPWR _7167_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_113_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4379_ _4588_/A _4935_/A _4605_/A _4621_/B VGND VGND VPWR VPWR _4732_/A sky130_fd_sc_hd__nor4_4
XFILLER_86_621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6118_ _6965_/Q _6025_/D _6115_/X _6117_/X VGND VGND VPWR VPWR _6119_/D sky130_fd_sc_hd__a211o_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7098_ _7098_/CLK _7098_/D fanout506/X VGND VGND VPWR VPWR _7098_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6049_ _7027_/Q _6049_/B VGND VGND VPWR VPWR _6049_/X sky130_fd_sc_hd__and2_1
XFILLER_37_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_20_csclk _6820_/CLK VGND VGND VPWR VPWR _7107_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_64_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_35_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7142_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_91_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3750_ _6716_/Q _4264_/A _4204_/A _6660_/Q VGND VGND VPWR VPWR _3750_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3681_ _7083_/Q _5520_/A _4028_/A _6522_/Q _3680_/X VGND VGND VPWR VPWR _3688_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_158_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5420_ _5552_/A0 hold781/X _5420_/S VGND VGND VPWR VPWR _5420_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5351_ _5573_/A0 _5351_/A1 _5357_/S VGND VGND VPWR VPWR _5351_/X sky130_fd_sc_hd__mux2_1
Xoutput204 _3921_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[36] sky130_fd_sc_hd__buf_12
Xoutput215 _6569_/Q VGND VGND VPWR VPWR mgmt_gpio_out[11] sky130_fd_sc_hd__buf_12
XFILLER_160_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput226 _6551_/Q VGND VGND VPWR VPWR mgmt_gpio_out[21] sky130_fd_sc_hd__buf_12
XFILLER_99_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput237 _6833_/Q VGND VGND VPWR VPWR mgmt_gpio_out[31] sky130_fd_sc_hd__buf_12
Xoutput248 _6561_/Q VGND VGND VPWR VPWR mgmt_gpio_out[7] sky130_fd_sc_hd__buf_12
X_4302_ _5459_/A0 hold299/X _4305_/S VGND VGND VPWR VPWR _4302_/X sky130_fd_sc_hd__mux2_1
Xoutput259 _3950_/Y VGND VGND VPWR VPWR pad_flash_io1_ieb sky130_fd_sc_hd__buf_12
XFILLER_114_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5282_ _5567_/A0 hold773/X _5285_/S VGND VGND VPWR VPWR _5282_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4233_ _6346_/A _3971_/S _3191_/A _4230_/X _4232_/X VGND VGND VPWR VPWR _6680_/D
+ sky130_fd_sc_hd__a2111o_1
X_7021_ _7136_/CLK _7021_/D fanout521/X VGND VGND VPWR VPWR _7021_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_114_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4164_ hold669/X _5549_/A0 _4164_/S VGND VGND VPWR VPWR _4164_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4095_ hold413/X _4094_/X _4103_/S VGND VGND VPWR VPWR _4095_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6805_ _7002_/CLK _6805_/D fanout498/X VGND VGND VPWR VPWR _6805_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_169_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4997_ _4997_/A _5036_/B VGND VGND VPWR VPWR _5009_/A sky130_fd_sc_hd__nor2_1
XFILLER_23_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6736_ _7070_/CLK _6736_/D fanout510/X VGND VGND VPWR VPWR _6736_/Q sky130_fd_sc_hd__dfrtp_4
X_3948_ _3948_/A VGND VGND VPWR VPWR _3948_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6667_ _7093_/CLK _6667_/D _6432_/A VGND VGND VPWR VPWR _6667_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_109_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3879_ _4339_/A _4339_/B _3879_/C VGND VGND VPWR VPWR _3887_/A sky130_fd_sc_hd__or3_1
XFILLER_192_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5618_ _7150_/Q _5618_/B VGND VGND VPWR VPWR _5622_/B sky130_fd_sc_hd__or2_1
XFILLER_137_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6598_ _6759_/CLK _6598_/D fanout489/X VGND VGND VPWR VPWR _6598_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_124_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5549_ _5549_/A0 hold653/X _5552_/S VGND VGND VPWR VPWR _5549_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout442 hold133/X VGND VGND VPWR VPWR hold127/A sky130_fd_sc_hd__clkbuf_16
Xfanout453 hold36/X VGND VGND VPWR VPWR _5557_/A0 sky130_fd_sc_hd__clkbuf_4
Xfanout464 _5459_/A0 VGND VGND VPWR VPWR _5573_/A0 sky130_fd_sc_hd__buf_6
Xfanout475 _6563_/Q VGND VGND VPWR VPWR _5650_/A sky130_fd_sc_hd__buf_8
XFILLER_59_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout486 _3946_/B VGND VGND VPWR VPWR _6426_/A sky130_fd_sc_hd__buf_6
XFILLER_19_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout497 fanout527/X VGND VGND VPWR VPWR fanout497/X sky130_fd_sc_hd__buf_4
XFILLER_58_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_554 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_6_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A VGND VGND VPWR VPWR _3937_/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_97_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4920_ _4659_/B _5021_/B _4692_/B _4646_/A _4919_/X VGND VGND VPWR VPWR _4920_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_45_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4851_ _4639_/B _4692_/B _4510_/C VGND VGND VPWR VPWR _4862_/A sky130_fd_sc_hd__o21ai_1
XTAP_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3802_ _6473_/Q _6472_/Q _6471_/Q VGND VGND VPWR VPWR _3834_/B sky130_fd_sc_hd__and3_2
X_4782_ _4606_/B _4606_/C _4793_/B VGND VGND VPWR VPWR _4802_/D sky130_fd_sc_hd__a21bo_1
X_6521_ _6707_/CLK _6521_/D _6433_/A VGND VGND VPWR VPWR _6521_/Q sky130_fd_sc_hd__dfrtp_2
X_3733_ _6970_/Q _5394_/A _3334_/Y _6914_/Q VGND VGND VPWR VPWR _3733_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6452_ net499_2/A _6452_/D _6407_/X VGND VGND VPWR VPWR hold38/A sky130_fd_sc_hd__dfrtp_1
X_3664_ _6891_/Q _3280_/Y _4294_/A _6742_/Q VGND VGND VPWR VPWR _3669_/B sky130_fd_sc_hd__a22o_1
XFILLER_106_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5403_ _5403_/A _5571_/B VGND VGND VPWR VPWR _5411_/S sky130_fd_sc_hd__nand2_8
X_3595_ input14/X _3268_/Y _3300_/Y _6997_/Q _3556_/X VGND VGND VPWR VPWR _3600_/B
+ sky130_fd_sc_hd__a221o_2
X_6383_ _6382_/X _6383_/A1 _6386_/S VGND VGND VPWR VPWR _7203_/D sky130_fd_sc_hd__mux2_1
X_5334_ _5496_/A0 hold914/X _5339_/S VGND VGND VPWR VPWR _5334_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5265_ _5586_/A0 hold997/X _5267_/S VGND VGND VPWR VPWR _5265_/X sky130_fd_sc_hd__mux2_1
X_7004_ _7129_/CLK _7004_/D fanout526/X VGND VGND VPWR VPWR _7004_/Q sky130_fd_sc_hd__dfrtp_4
X_4216_ _4216_/A _5580_/B VGND VGND VPWR VPWR _4221_/S sky130_fd_sc_hd__nand2_2
X_5196_ _6395_/A0 _5196_/A1 _5199_/S VGND VGND VPWR VPWR _5196_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4147_ _4147_/A _6392_/B VGND VGND VPWR VPWR _4152_/S sky130_fd_sc_hd__nand2_4
XFILLER_95_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4078_ hold431/X _4077_/X _4086_/S VGND VGND VPWR VPWR _4078_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6719_ _7074_/CLK _6719_/D fanout501/X VGND VGND VPWR VPWR _6719_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_177_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap406 _6033_/X VGND VGND VPWR VPWR _6205_/B1 sky130_fd_sc_hd__buf_12
XFILLER_7_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap417 _5982_/X VGND VGND VPWR VPWR _6024_/A sky130_fd_sc_hd__buf_12
XFILLER_115_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold709 _6933_/Q VGND VGND VPWR VPWR hold709/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3380_ _7187_/Q _6817_/Q _6818_/Q VGND VGND VPWR VPWR _3380_/X sky130_fd_sc_hd__mux2_4
XFILLER_156_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5050_ _5050_/A _5050_/B _5050_/C VGND VGND VPWR VPWR _5050_/X sky130_fd_sc_hd__and3_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1409 _6644_/Q VGND VGND VPWR VPWR hold1409/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4001_ _4001_/A _5535_/B VGND VGND VPWR VPWR _4009_/S sky130_fd_sc_hd__nand2_8
XFILLER_77_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5952_ _6530_/Q _5676_/X _5703_/X _6605_/Q _5951_/X VGND VGND VPWR VPWR _5957_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_18_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4903_ _5013_/A _5016_/A _4781_/Y _4672_/A VGND VGND VPWR VPWR _4903_/X sky130_fd_sc_hd__o22a_1
X_5883_ _7208_/Q _5671_/X _5676_/X _6527_/Q VGND VGND VPWR VPWR _5883_/X sky130_fd_sc_hd__a22o_1
XFILLER_61_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4834_ _4947_/A _4933_/A _5035_/B _4832_/B _4784_/A VGND VGND VPWR VPWR _4835_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_60_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4765_ _4993_/A _4512_/B _4746_/Y _4985_/B _4764_/X VGND VGND VPWR VPWR _4765_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_193_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6504_ _7033_/CLK _6504_/D fanout502/X VGND VGND VPWR VPWR _6504_/Q sky130_fd_sc_hd__dfrtp_2
X_3716_ _7059_/Q _3329_/Y _5259_/A _6851_/Q _3715_/X VGND VGND VPWR VPWR _3721_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_147_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4696_ _5076_/A _4694_/B _4707_/B _4666_/B VGND VGND VPWR VPWR _4696_/X sky130_fd_sc_hd__o22a_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6435_ _6441_/A _6441_/B VGND VGND VPWR VPWR _6435_/X sky130_fd_sc_hd__and2_1
X_3647_ input13/X _3268_/Y _5225_/A _6821_/Q VGND VGND VPWR VPWR _3647_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6366_ _6700_/Q _6366_/A2 _6366_/B1 _6699_/Q VGND VGND VPWR VPWR _6366_/X sky130_fd_sc_hd__a22o_1
X_3578_ _7114_/Q _5553_/A _4276_/A _6729_/Q VGND VGND VPWR VPWR _3578_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5317_ _5557_/A0 hold645/X hold23/X VGND VGND VPWR VPWR _5317_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6297_ _6614_/Q _6023_/C _6020_/X _6709_/Q VGND VGND VPWR VPWR _6297_/X sky130_fd_sc_hd__a22o_1
XFILLER_142_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold14 hold14/A VGND VGND VPWR VPWR hold14/X sky130_fd_sc_hd__dlygate4sd3_1
X_5248_ _5569_/A0 hold123/X hold14/X VGND VGND VPWR VPWR _5248_/X sky130_fd_sc_hd__mux2_1
Xhold25 hold25/A VGND VGND VPWR VPWR hold25/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold36 hold36/A VGND VGND VPWR VPWR hold36/X sky130_fd_sc_hd__buf_8
XFILLER_29_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold47 hold47/A VGND VGND VPWR VPWR hold47/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 hold58/A VGND VGND VPWR VPWR hold58/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_48 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold69 hold69/A VGND VGND VPWR VPWR hold69/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5179_ _5023_/A _4679_/B _4679_/X _4510_/A _4510_/B VGND VGND VPWR VPWR _5180_/D
+ sky130_fd_sc_hd__o2111a_1
XFILLER_29_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4550_ _4621_/B _4971_/B VGND VGND VPWR VPWR _4793_/B sky130_fd_sc_hd__xnor2_1
XFILLER_128_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3501_ _7115_/Q _3278_/Y _5221_/B _6813_/Q _3500_/X VGND VGND VPWR VPWR _3515_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold506 _6921_/Q VGND VGND VPWR VPWR hold506/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4481_ _5018_/A _4638_/B VGND VGND VPWR VPWR _5013_/A sky130_fd_sc_hd__or2_4
XFILLER_156_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold517 _3997_/X VGND VGND VPWR VPWR _6494_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold528 _6477_/Q VGND VGND VPWR VPWR hold528/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6220_ _6220_/A0 _6219_/X _6319_/S VGND VGND VPWR VPWR _7182_/D sky130_fd_sc_hd__mux2_1
Xhold539 _5402_/X VGND VGND VPWR VPWR _6977_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3432_ _7063_/Q _5493_/A _5221_/B _3413_/X VGND VGND VPWR VPWR _3432_/X sky130_fd_sc_hd__a22o_1
XFILLER_103_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3363_ _7089_/Q _5520_/A hold22/A _6905_/Q _3362_/X VGND VGND VPWR VPWR _3363_/X
+ sky130_fd_sc_hd__a221o_1
X_6151_ _7031_/Q _6049_/B _6202_/B1 _7007_/Q _6148_/X VGND VGND VPWR VPWR _6156_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ _5102_/A _5102_/B VGND VGND VPWR VPWR _5103_/B sky130_fd_sc_hd__nor2_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3294_ _3536_/A _3546_/B VGND VGND VPWR VPWR _5535_/A sky130_fd_sc_hd__nor2_8
XFILLER_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6082_ _6940_/Q _6024_/D _6027_/D _6884_/Q VGND VGND VPWR VPWR _6082_/X sky130_fd_sc_hd__a22o_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1206 _5386_/X VGND VGND VPWR VPWR _6962_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1217 _5194_/X VGND VGND VPWR VPWR _6798_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1228 _6753_/Q VGND VGND VPWR VPWR _4309_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5033_ _6362_/A _5033_/B _5033_/C VGND VGND VPWR VPWR _5033_/X sky130_fd_sc_hd__or3_1
Xhold1239 _5224_/X VGND VGND VPWR VPWR _6820_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6984_ _7141_/CLK _6984_/D fanout504/X VGND VGND VPWR VPWR _6984_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_53_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5935_ _5935_/A _5935_/B _5935_/C _5935_/D VGND VGND VPWR VPWR _5935_/X sky130_fd_sc_hd__or4_1
XFILLER_80_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5866_ _6660_/Q _5685_/X _5865_/X VGND VGND VPWR VPWR _5869_/C sky130_fd_sc_hd__a21o_1
XFILLER_33_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4817_ _4983_/C _4817_/B _4817_/C _4816_/X VGND VGND VPWR VPWR _4818_/A sky130_fd_sc_hd__or4b_1
X_5797_ _6935_/Q _5670_/X _5671_/X _7063_/Q VGND VGND VPWR VPWR _5797_/X sky130_fd_sc_hd__a22o_1
XFILLER_178_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4748_ _4981_/B _4872_/A VGND VGND VPWR VPWR _4818_/B sky130_fd_sc_hd__nor2_1
XFILLER_135_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4679_ _5023_/B _4679_/B VGND VGND VPWR VPWR _4679_/X sky130_fd_sc_hd__or2_1
X_6418_ _6441_/A _6440_/B VGND VGND VPWR VPWR _6418_/X sky130_fd_sc_hd__and2_1
XFILLER_162_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6349_ _6349_/A0 _3790_/X _6356_/S VGND VGND VPWR VPWR _7189_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_759 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput104 wb_adr_i[14] VGND VGND VPWR VPWR _4338_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput115 wb_adr_i[24] VGND VGND VPWR VPWR _3880_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_48_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput126 wb_adr_i[5] VGND VGND VPWR VPWR _4605_/A sky130_fd_sc_hd__buf_6
Xinput137 wb_dat_i[14] VGND VGND VPWR VPWR _6381_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput148 wb_dat_i[24] VGND VGND VPWR VPWR _6364_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput159 wb_dat_i[5] VGND VGND VPWR VPWR _6378_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3981_ hold38/X hold469/X _3981_/S VGND VGND VPWR VPWR _3981_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5720_ _6923_/Q _5955_/A2 _5693_/X _6899_/Q VGND VGND VPWR VPWR _5720_/X sky130_fd_sc_hd__a22o_1
XFILLER_43_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5651_ _5651_/A _5651_/B VGND VGND VPWR VPWR _6171_/S sky130_fd_sc_hd__nor2_4
XFILLER_30_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4602_ _4846_/A _4570_/B _4570_/D _4778_/B _4601_/X VGND VGND VPWR VPWR _4647_/A
+ sky130_fd_sc_hd__a41o_1
XFILLER_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5582_ hold9/X _7136_/Q hold70/X VGND VGND VPWR VPWR _5582_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4533_ _4846_/C _4993_/A VGND VGND VPWR VPWR _4802_/A sky130_fd_sc_hd__nand2_8
XFILLER_116_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold303 _6728_/Q VGND VGND VPWR VPWR hold303/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold314 _5469_/X VGND VGND VPWR VPWR _7036_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold325 _6867_/Q VGND VGND VPWR VPWR hold325/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold336 _5405_/X VGND VGND VPWR VPWR _6979_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4464_ _4838_/B VGND VGND VPWR VPWR _4464_/Y sky130_fd_sc_hd__inv_2
Xhold347 _6843_/Q VGND VGND VPWR VPWR hold347/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold358 _5432_/X VGND VGND VPWR VPWR _7003_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6203_ _6993_/Q _6203_/A2 _6024_/C _6913_/Q VGND VGND VPWR VPWR _6203_/X sky130_fd_sc_hd__a22o_1
Xhold369 _6510_/Q VGND VGND VPWR VPWR hold369/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3415_ hold95/X _3729_/B VGND VGND VPWR VPWR _4104_/A sky130_fd_sc_hd__nor2_8
X_7183_ _7183_/CLK _7183_/D fanout490/X VGND VGND VPWR VPWR _7183_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4395_ _4461_/B VGND VGND VPWR VPWR _4395_/Y sky130_fd_sc_hd__inv_2
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6134_ _7139_/Q _6308_/A2 _6338_/B1 _7099_/Q _6123_/X VGND VGND VPWR VPWR _6134_/X
+ sky130_fd_sc_hd__a221o_4
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3346_ _6937_/Q _5349_/A _5331_/A _6921_/Q VGND VGND VPWR VPWR _3346_/X sky130_fd_sc_hd__a22o_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1003 _7063_/Q VGND VGND VPWR VPWR _5499_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6065_ _6851_/Q _6027_/A _6329_/B1 _7035_/Q _6048_/X VGND VGND VPWR VPWR _6068_/C
+ sky130_fd_sc_hd__a221o_1
Xhold1014 _5364_/X VGND VGND VPWR VPWR _6943_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3277_ hold28/X hold75/X VGND VGND VPWR VPWR _3526_/A sky130_fd_sc_hd__nand2_8
Xhold1025 _6503_/Q VGND VGND VPWR VPWR _4007_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1036 _5431_/X VGND VGND VPWR VPWR _7002_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1047 _7121_/Q VGND VGND VPWR VPWR _5565_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5016_ _5016_/A _5016_/B VGND VGND VPWR VPWR _5017_/B sky130_fd_sc_hd__and2_1
Xhold1058 _5226_/X VGND VGND VPWR VPWR _6821_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1069 _7103_/Q VGND VGND VPWR VPWR _5545_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_209 _6030_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6967_ _7108_/CLK _6967_/D fanout523/X VGND VGND VPWR VPWR _6967_/Q sky130_fd_sc_hd__dfrtp_2
X_5918_ _6708_/Q _5675_/X _5700_/X _6508_/Q _5917_/X VGND VGND VPWR VPWR _5923_/B
+ sky130_fd_sc_hd__a221o_1
X_6898_ _7139_/CLK _6898_/D fanout518/X VGND VGND VPWR VPWR _6898_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_179_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5849_ _6969_/Q _5675_/X _5700_/X _7033_/Q _5848_/X VGND VGND VPWR VPWR _5857_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_166_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold870 _6513_/Q VGND VGND VPWR VPWR hold870/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold881 _5546_/X VGND VGND VPWR VPWR _7104_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold892 _7000_/Q VGND VGND VPWR VPWR hold892/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1570 _6697_/Q VGND VGND VPWR VPWR _3191_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1581 _6817_/Q VGND VGND VPWR VPWR hold876/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_83_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1592 _7101_/Q VGND VGND VPWR VPWR hold902/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3200_ _7114_/Q VGND VGND VPWR VPWR _3200_/Y sky130_fd_sc_hd__inv_2
X_4180_ _6693_/Q _6348_/B VGND VGND VPWR VPWR _4188_/S sky130_fd_sc_hd__and2_4
XFILLER_79_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6821_ _7136_/CLK _6821_/D fanout520/X VGND VGND VPWR VPWR _6821_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6752_ _6755_/CLK _6752_/D fanout497/X VGND VGND VPWR VPWR _6752_/Q sky130_fd_sc_hd__dfrtp_2
X_3964_ hold12/X _3967_/S hold111/X VGND VGND VPWR VPWR _3964_/X sky130_fd_sc_hd__o21a_4
X_5703_ _5938_/B _5703_/B _5703_/C VGND VGND VPWR VPWR _5703_/X sky130_fd_sc_hd__and3_4
XFILLER_176_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6683_ _6683_/CLK hold63/X fanout511/X VGND VGND VPWR VPWR _6683_/Q sky130_fd_sc_hd__dfstp_1
X_3895_ _7144_/Q _7146_/Q _7147_/Q _7145_/Q VGND VGND VPWR VPWR _3896_/B sky130_fd_sc_hd__or4b_1
X_5634_ _5637_/B _6039_/A VGND VGND VPWR VPWR _5634_/Y sky130_fd_sc_hd__nand2_1
XFILLER_136_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5565_ _5574_/A0 _5565_/A1 _5570_/S VGND VGND VPWR VPWR _5565_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold100 hold100/A VGND VGND VPWR VPWR hold2/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold111 _3963_/Y VGND VGND VPWR VPWR hold111/X sky130_fd_sc_hd__dlygate4sd3_1
X_4516_ _4742_/A _4516_/B VGND VGND VPWR VPWR _4850_/A sky130_fd_sc_hd__nand2_1
Xhold122 _5498_/X VGND VGND VPWR VPWR _7062_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5496_ _5496_/A0 hold817/X _5501_/S VGND VGND VPWR VPWR _5496_/X sky130_fd_sc_hd__mux2_1
Xhold133 hold133/A VGND VGND VPWR VPWR hold133/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 _6479_/Q VGND VGND VPWR VPWR hold144/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold155 _5427_/X VGND VGND VPWR VPWR _6999_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 _5585_/X VGND VGND VPWR VPWR _7139_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4447_ _4742_/A _4759_/B VGND VGND VPWR VPWR _4447_/Y sky130_fd_sc_hd__nand2_1
Xhold177 _6934_/Q VGND VGND VPWR VPWR hold177/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 _5426_/X VGND VGND VPWR VPWR _6998_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold199 _6893_/Q VGND VGND VPWR VPWR hold199/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7166_ _7182_/CLK _7166_/D fanout500/X VGND VGND VPWR VPWR _7166_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4378_ _4546_/A _4547_/A VGND VGND VPWR VPWR _5018_/A sky130_fd_sc_hd__or2_4
XFILLER_86_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_1_csclk _7018_/CLK VGND VGND VPWR VPWR _7093_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6117_ _7138_/Q _6308_/A2 _6338_/B1 _7098_/Q _6116_/X VGND VGND VPWR VPWR _6117_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3329_ _3495_/A _3340_/B VGND VGND VPWR VPWR _3329_/Y sky130_fd_sc_hd__nor2_4
XFILLER_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7097_ _7098_/CLK _7097_/D fanout505/X VGND VGND VPWR VPWR _7097_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_85_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6048_ _6499_/Q _6323_/A2 _6024_/B _6931_/Q VGND VGND VPWR VPWR _6048_/X sky130_fd_sc_hd__a22o_1
XTAP_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3680_ _6707_/Q _4252_/A _4204_/A _6661_/Q VGND VGND VPWR VPWR _3680_/X sky130_fd_sc_hd__a22o_1
XFILLER_158_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5350_ _5581_/A0 _5350_/A1 _5357_/S VGND VGND VPWR VPWR _5350_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput205 _3920_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[37] sky130_fd_sc_hd__buf_12
Xoutput216 _6570_/Q VGND VGND VPWR VPWR mgmt_gpio_out[12] sky130_fd_sc_hd__buf_12
XFILLER_160_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput227 _6552_/Q VGND VGND VPWR VPWR mgmt_gpio_out[22] sky130_fd_sc_hd__buf_12
Xoutput238 _3923_/X VGND VGND VPWR VPWR mgmt_gpio_out[32] sky130_fd_sc_hd__buf_12
X_4301_ _5521_/A0 _4301_/A1 _4305_/S VGND VGND VPWR VPWR _4301_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput249 _3928_/X VGND VGND VPWR VPWR mgmt_gpio_out[8] sky130_fd_sc_hd__buf_12
X_5281_ _5557_/A0 hold667/X _5285_/S VGND VGND VPWR VPWR _5281_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7020_ _7050_/CLK _7020_/D fanout499/X VGND VGND VPWR VPWR _7020_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_114_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4232_ _6696_/Q _4232_/B VGND VGND VPWR VPWR _4232_/X sky130_fd_sc_hd__or2_2
XFILLER_141_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4163_ hold181/X hold36/X _4164_/S VGND VGND VPWR VPWR _4163_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4094_ hold197/X hold36/X _4102_/S VGND VGND VPWR VPWR _4094_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6804_ _7002_/CLK _6804_/D fanout498/X VGND VGND VPWR VPWR _6804_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4996_ _4996_/A _5036_/B VGND VGND VPWR VPWR _5008_/B sky130_fd_sc_hd__nor2_1
X_6735_ _6759_/CLK _6735_/D fanout489/X VGND VGND VPWR VPWR _6735_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3947_ _6460_/Q _3947_/B VGND VGND VPWR VPWR _3948_/A sky130_fd_sc_hd__nand2b_1
XFILLER_149_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6666_ _6764_/CLK _6666_/D _3946_/B VGND VGND VPWR VPWR _6666_/Q sky130_fd_sc_hd__dfrtp_1
X_3878_ _4339_/C _4339_/D _4338_/A _4338_/B VGND VGND VPWR VPWR _3879_/C sky130_fd_sc_hd__or4_1
XFILLER_109_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5617_ _5650_/B _5705_/B _5706_/B _5617_/B1 _5610_/X VGND VGND VPWR VPWR _7149_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_164_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6597_ _7211_/CLK _6597_/D fanout489/X VGND VGND VPWR VPWR _6597_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_136_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5548_ _5584_/A0 hold437/X _5552_/S VGND VGND VPWR VPWR _5548_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5479_ _5584_/A0 hold492/X hold79/X VGND VGND VPWR VPWR _5479_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout432 _4596_/X VGND VGND VPWR VPWR _5021_/B sky130_fd_sc_hd__buf_8
Xfanout443 _5558_/A0 VGND VGND VPWR VPWR _6397_/A0 sky130_fd_sc_hd__buf_8
X_7149_ _7183_/CLK _7149_/D fanout499/X VGND VGND VPWR VPWR _7149_/Q sky130_fd_sc_hd__dfstp_1
Xfanout454 hold35/X VGND VGND VPWR VPWR hold36/A sky130_fd_sc_hd__buf_8
XFILLER_101_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout465 hold9/X VGND VGND VPWR VPWR _5459_/A0 sky130_fd_sc_hd__buf_8
Xfanout487 fanout527/X VGND VGND VPWR VPWR _3946_/B sky130_fd_sc_hd__buf_6
Xfanout498 fanout500/X VGND VGND VPWR VPWR fanout498/X sky130_fd_sc_hd__buf_8
XFILLER_100_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4850_ _4850_/A _4850_/B VGND VGND VPWR VPWR _5124_/B sky130_fd_sc_hd__nand2_1
XTAP_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3801_ _3801_/A _3801_/B VGND VGND VPWR VPWR _6471_/D sky130_fd_sc_hd__xor2_1
XFILLER_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4781_ _4781_/A _4781_/B VGND VGND VPWR VPWR _4781_/Y sky130_fd_sc_hd__nand2_2
X_6520_ _6708_/CLK _6520_/D fanout494/X VGND VGND VPWR VPWR _6520_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_119_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3732_ input52/X _5232_/A hold69/A _7135_/Q VGND VGND VPWR VPWR _3732_/X sky130_fd_sc_hd__a22o_2
XFILLER_9_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6451_ net499_2/A _6451_/D _6406_/X VGND VGND VPWR VPWR hold1/A sky130_fd_sc_hd__dfrtp_1
X_3663_ _6987_/Q _3298_/Y _5394_/A _6971_/Q VGND VGND VPWR VPWR _3669_/A sky130_fd_sc_hd__a22o_1
X_5402_ hold538/X _5552_/A0 _5402_/S VGND VGND VPWR VPWR _5402_/X sky130_fd_sc_hd__mux2_1
X_6382_ _6698_/Q _6382_/A2 _6382_/B1 _6390_/A2 _6381_/X VGND VGND VPWR VPWR _6382_/X
+ sky130_fd_sc_hd__a221o_1
X_3594_ _7061_/Q _3329_/Y _5529_/A _7093_/Q _3555_/X VGND VGND VPWR VPWR _3600_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5333_ _5573_/A0 hold888/X _5339_/S VGND VGND VPWR VPWR _5333_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5264_ _5567_/A0 hold731/X _5267_/S VGND VGND VPWR VPWR _5264_/X sky130_fd_sc_hd__mux2_1
X_7003_ _7050_/CLK _7003_/D fanout499/X VGND VGND VPWR VPWR _7003_/Q sky130_fd_sc_hd__dfstp_4
X_4215_ hold363/X _5534_/A1 _4215_/S VGND VGND VPWR VPWR _4215_/X sky130_fd_sc_hd__mux2_1
X_5195_ _6394_/A0 _5195_/A1 _5199_/S VGND VGND VPWR VPWR _5195_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4146_ _5549_/A0 hold585/X _4146_/S VGND VGND VPWR VPWR _4146_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4077_ hold295/X _5539_/A1 _4085_/S VGND VGND VPWR VPWR _4077_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4979_ _5142_/A _5114_/B _4979_/C _4979_/D VGND VGND VPWR VPWR _4979_/X sky130_fd_sc_hd__or4_1
X_6718_ _7074_/CLK _6718_/D fanout501/X VGND VGND VPWR VPWR _6718_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6649_ _7187_/CLK _6649_/D VGND VGND VPWR VPWR _6649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_34_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7132_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_117_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_49_csclk _6970_/CLK VGND VGND VPWR VPWR _6883_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_87_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap407 _6020_/X VGND VGND VPWR VPWR _6025_/D sky130_fd_sc_hd__buf_12
Xmax_cap418 _5696_/X VGND VGND VPWR VPWR _5966_/B1 sky130_fd_sc_hd__buf_12
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4000_ hold583/X _5552_/A0 _4000_/S VGND VGND VPWR VPWR _4000_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5951_ _6775_/Q _5663_/X _5671_/X _7211_/Q VGND VGND VPWR VPWR _5951_/X sky130_fd_sc_hd__a22o_1
XFILLER_52_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4902_ _5023_/B _4675_/A _4900_/X _4666_/B _4668_/X VGND VGND VPWR VPWR _4902_/X
+ sky130_fd_sc_hd__o221a_1
X_5882_ _5882_/A0 _5881_/X _6319_/S VGND VGND VPWR VPWR _7170_/D sky130_fd_sc_hd__mux2_1
XFILLER_178_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4833_ _4461_/B _4832_/B _4484_/X VGND VGND VPWR VPWR _4833_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_33_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4764_ _4764_/A _4986_/B _4764_/C VGND VGND VPWR VPWR _4764_/X sky130_fd_sc_hd__or3_1
XFILLER_193_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6503_ _7055_/CLK _6503_/D fanout523/X VGND VGND VPWR VPWR _6503_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_159_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3715_ _6732_/Q _4282_/A _5229_/A _6825_/Q VGND VGND VPWR VPWR _3715_/X sky130_fd_sc_hd__a22o_2
XFILLER_174_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4695_ _5076_/A _4582_/B _4694_/B _5016_/B _4694_/X VGND VGND VPWR VPWR _4698_/C
+ sky130_fd_sc_hd__o221a_1
X_6434_ _6441_/A _6441_/B VGND VGND VPWR VPWR _6434_/X sky130_fd_sc_hd__and2_1
X_3646_ _6476_/Q _3966_/A _5466_/A _7036_/Q _3645_/X VGND VGND VPWR VPWR _3651_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_162_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6365_ _6364_/X _6365_/A1 _6386_/S VGND VGND VPWR VPWR _7197_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3577_ _6885_/Q _5295_/A _5322_/A _6909_/Q _3576_/X VGND VGND VPWR VPWR _3582_/B
+ sky130_fd_sc_hd__a221o_1
X_5316_ _5574_/A0 _5316_/A1 hold23/X VGND VGND VPWR VPWR _5316_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6296_ _6729_/Q _6320_/A2 _6320_/B1 _6619_/Q VGND VGND VPWR VPWR _6296_/X sky130_fd_sc_hd__a22o_2
XFILLER_130_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5247_ _5550_/A0 hold441/X hold14/X VGND VGND VPWR VPWR _5247_/X sky130_fd_sc_hd__mux2_1
Xhold15 hold15/A VGND VGND VPWR VPWR hold15/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 hold26/A VGND VGND VPWR VPWR hold26/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 hold37/A VGND VGND VPWR VPWR hold37/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold48 hold48/A VGND VGND VPWR VPWR hold48/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold59 hold59/A VGND VGND VPWR VPWR hold59/X sky130_fd_sc_hd__dlygate4sd3_1
X_5178_ _5178_/A _5178_/B _5178_/C _5178_/D VGND VGND VPWR VPWR _5178_/X sky130_fd_sc_hd__or4_1
XFILLER_56_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4129_ _4129_/A _6392_/B VGND VGND VPWR VPWR _4134_/S sky130_fd_sc_hd__and2_1
XFILLER_29_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_764 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3500_ input7/X _3295_/Y _3300_/Y _6998_/Q VGND VGND VPWR VPWR _3500_/X sky130_fd_sc_hd__a22o_1
XFILLER_190_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4480_ _4588_/A _4935_/A _4793_/A _4621_/B VGND VGND VPWR VPWR _4638_/B sky130_fd_sc_hd__or4_4
Xhold507 _5339_/X VGND VGND VPWR VPWR _6921_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 _6873_/Q VGND VGND VPWR VPWR hold518/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold529 _3974_/X VGND VGND VPWR VPWR _6477_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3431_ _3431_/A _3431_/B _3431_/C _3431_/D VGND VGND VPWR VPWR _3447_/A sky130_fd_sc_hd__or4_1
X_6150_ _7079_/Q _5994_/X _5998_/Y _7015_/Q _6149_/X VGND VGND VPWR VPWR _6156_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3362_ _6897_/Q _5304_/A _5322_/A _6913_/Q VGND VGND VPWR VPWR _3362_/X sky130_fd_sc_hd__a22o_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5101_ _5114_/C _5145_/B _5112_/D _5101_/D VGND VGND VPWR VPWR _5102_/B sky130_fd_sc_hd__or4_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6081_ _6852_/Q _6027_/A _6024_/B _6932_/Q _6080_/X VGND VGND VPWR VPWR _6084_/C
+ sky130_fd_sc_hd__a221o_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3293_ hold28/X _3313_/B VGND VGND VPWR VPWR _3546_/B sky130_fd_sc_hd__nand2_8
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1207 _6948_/Q VGND VGND VPWR VPWR _5370_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5032_ _5112_/C _5030_/X _5071_/C VGND VGND VPWR VPWR _5033_/C sky130_fd_sc_hd__o21ba_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1218 _6634_/Q VGND VGND VPWR VPWR _4175_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1229 _4309_/X VGND VGND VPWR VPWR _6753_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_731 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6983_ _7055_/CLK _6983_/D fanout523/X VGND VGND VPWR VPWR _6983_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_80_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5934_ _6663_/Q _5685_/X _5966_/B1 _6519_/Q _5933_/X VGND VGND VPWR VPWR _5935_/D
+ sky130_fd_sc_hd__a221o_1
X_5865_ _6665_/Q _5677_/X _5966_/B1 _6516_/Q VGND VGND VPWR VPWR _5865_/X sky130_fd_sc_hd__a22o_1
XFILLER_33_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4816_ _4997_/A _4802_/A _5076_/B _4677_/B VGND VGND VPWR VPWR _4816_/X sky130_fd_sc_hd__o22a_1
X_5796_ _6975_/Q _5960_/B _5691_/B VGND VGND VPWR VPWR _5796_/X sky130_fd_sc_hd__o21a_1
XFILLER_193_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4747_ _5003_/A _5036_/A VGND VGND VPWR VPWR _4985_/B sky130_fd_sc_hd__nor2_1
XFILLER_147_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4678_ _5018_/C _4692_/B VGND VGND VPWR VPWR _4916_/B sky130_fd_sc_hd__or2_2
XFILLER_162_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6417_ _6433_/A _6441_/B VGND VGND VPWR VPWR _6417_/X sky130_fd_sc_hd__and2_1
XFILLER_107_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3629_ input37/X _3751_/A2 _4204_/A _6662_/Q _3606_/X VGND VGND VPWR VPWR _3632_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_150_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6348_ _6692_/Q _6348_/B VGND VGND VPWR VPWR _6356_/S sky130_fd_sc_hd__and2_4
XFILLER_1_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_644 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6279_ _6713_/Q _6009_/X _6038_/Y _6723_/Q _6273_/X VGND VGND VPWR VPWR _6280_/D
+ sky130_fd_sc_hd__a221o_1
Xinput105 wb_adr_i[15] VGND VGND VPWR VPWR _4338_/C sky130_fd_sc_hd__clkbuf_1
Xinput116 wb_adr_i[25] VGND VGND VPWR VPWR input116/X sky130_fd_sc_hd__clkbuf_1
XFILLER_76_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput127 wb_adr_i[6] VGND VGND VPWR VPWR _4588_/A sky130_fd_sc_hd__buf_4
XFILLER_48_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput138 wb_dat_i[15] VGND VGND VPWR VPWR _6384_/B1 sky130_fd_sc_hd__clkbuf_1
Xinput149 wb_dat_i[25] VGND VGND VPWR VPWR _6366_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_57_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3980_ hold916/X _5587_/A0 _3982_/S VGND VGND VPWR VPWR _3980_/X sky130_fd_sc_hd__mux2_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5650_ _5650_/A _5650_/B VGND VGND VPWR VPWR _5650_/Y sky130_fd_sc_hd__nor2_4
XFILLER_188_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4601_ _4797_/A _4572_/Y _4600_/X _4952_/A _5112_/A VGND VGND VPWR VPWR _4601_/X
+ sky130_fd_sc_hd__a2111o_1
X_5581_ _5581_/A0 _5581_/A1 hold70/X VGND VGND VPWR VPWR _5581_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4532_ _4570_/D _4532_/B VGND VGND VPWR VPWR _4971_/A sky130_fd_sc_hd__nor2_2
XFILLER_191_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold304 _4279_/X VGND VGND VPWR VPWR _6728_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold315 _6963_/Q VGND VGND VPWR VPWR hold315/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold326 _5279_/X VGND VGND VPWR VPWR _6867_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4463_ _4474_/A _4944_/A _4462_/Y VGND VGND VPWR VPWR _4846_/D sky130_fd_sc_hd__nor3b_4
Xhold337 _6955_/Q VGND VGND VPWR VPWR hold337/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 _5252_/X VGND VGND VPWR VPWR _6843_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6202_ _7033_/Q _6049_/B _6202_/B1 _7009_/Q VGND VGND VPWR VPWR _6202_/X sky130_fd_sc_hd__a22o_1
XFILLER_171_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold359 _7035_/Q VGND VGND VPWR VPWR hold359/X sky130_fd_sc_hd__dlygate4sd3_1
X_3414_ hold56/X hold67/X VGND VGND VPWR VPWR _3729_/B sky130_fd_sc_hd__nand2_8
X_7182_ _7182_/CLK _7182_/D fanout499/X VGND VGND VPWR VPWR _7182_/Q sky130_fd_sc_hd__dfrtp_1
X_4394_ _4489_/A _4932_/A VGND VGND VPWR VPWR _4461_/B sky130_fd_sc_hd__or2_2
XFILLER_98_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6133_ _7070_/Q _6272_/B _6128_/X _6130_/X _6132_/X VGND VGND VPWR VPWR _6133_/X
+ sky130_fd_sc_hd__a2111o_2
X_3345_ _6497_/Q _3992_/A _5511_/A _7081_/Q VGND VGND VPWR VPWR _3345_/X sky130_fd_sc_hd__a22o_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6064_ _6859_/Q _6326_/A2 _6021_/Y _6883_/Q _6063_/X VGND VGND VPWR VPWR _6068_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_100_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1004 _5499_/X VGND VGND VPWR VPWR _7063_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3276_ hold74/X hold66/X VGND VGND VPWR VPWR hold75/A sky130_fd_sc_hd__nor2_8
Xhold1015 _6871_/Q VGND VGND VPWR VPWR _5283_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1026 _4007_/X VGND VGND VPWR VPWR _6503_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5015_ _5107_/C _5015_/B _5015_/C VGND VGND VPWR VPWR _5019_/B sky130_fd_sc_hd__or3_1
Xhold1037 _6860_/Q VGND VGND VPWR VPWR _5271_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1048 _5565_/X VGND VGND VPWR VPWR _7121_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1059 _6792_/Q VGND VGND VPWR VPWR _5186_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6966_ _7082_/CLK _6966_/D _3873_/A VGND VGND VPWR VPWR _6966_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_41_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5917_ _6773_/Q _5663_/X _5689_/X _5916_/X VGND VGND VPWR VPWR _5917_/X sky130_fd_sc_hd__a22o_1
X_6897_ _7065_/CLK _6897_/D fanout517/X VGND VGND VPWR VPWR _6897_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_167_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5848_ _7009_/Q _5664_/X _5848_/B1 _7049_/Q VGND VGND VPWR VPWR _5848_/X sky130_fd_sc_hd__a22o_1
X_5779_ _6950_/Q _5666_/X _5685_/X _6910_/Q VGND VGND VPWR VPWR _5779_/X sky130_fd_sc_hd__a22o_1
XFILLER_166_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold860 _7109_/Q VGND VGND VPWR VPWR hold860/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_174_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold871 _4019_/X VGND VGND VPWR VPWR _6513_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold882 _7032_/Q VGND VGND VPWR VPWR hold882/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold893 _5428_/X VGND VGND VPWR VPWR _7000_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1560 _3855_/X VGND VGND VPWR VPWR _6455_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1571 _6582_/Q VGND VGND VPWR VPWR hold783/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1582 _6594_/Q VGND VGND VPWR VPWR hold227/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1593 hold46/A VGND VGND VPWR VPWR _3815_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6820_ _6820_/CLK _6820_/D fanout511/X VGND VGND VPWR VPWR _6820_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_51_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6751_ _6759_/CLK _6751_/D fanout489/X VGND VGND VPWR VPWR _6751_/Q sky130_fd_sc_hd__dfrtp_2
X_3963_ hold110/X _3971_/S VGND VGND VPWR VPWR _3963_/Y sky130_fd_sc_hd__nand2b_1
X_5702_ _7152_/Q _5703_/B _5703_/C VGND VGND VPWR VPWR _5702_/X sky130_fd_sc_hd__and3_4
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_1_1_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
X_6682_ _6683_/CLK hold90/X fanout511/X VGND VGND VPWR VPWR hold89/A sky130_fd_sc_hd__dfrtp_4
XFILLER_31_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3894_ _6700_/Q _3876_/X _3894_/B1 VGND VGND VPWR VPWR _6700_/D sky130_fd_sc_hd__a21o_1
X_5633_ _7156_/Q _7155_/Q VGND VGND VPWR VPWR _6039_/A sky130_fd_sc_hd__and2_2
XFILLER_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5564_ _5573_/A0 hold878/X _5570_/S VGND VGND VPWR VPWR _5564_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4515_ _4515_/A _4515_/B _4515_/C _4863_/A VGND VGND VPWR VPWR _4515_/X sky130_fd_sc_hd__and4_1
Xhold101 hold2/X VGND VGND VPWR VPWR hold101/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 hold137/X VGND VGND VPWR VPWR _5203_/B sky130_fd_sc_hd__buf_6
X_5495_ _5573_/A0 hold850/X _5501_/S VGND VGND VPWR VPWR _5495_/X sky130_fd_sc_hd__mux2_1
Xhold123 hold123/A VGND VGND VPWR VPWR hold123/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 _3998_/X VGND VGND VPWR VPWR _6495_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 _3978_/X VGND VGND VPWR VPWR _6479_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 _6846_/Q VGND VGND VPWR VPWR hold156/X sky130_fd_sc_hd__dlygate4sd3_1
X_4446_ _4872_/A VGND VGND VPWR VPWR _4446_/Y sky130_fd_sc_hd__inv_2
Xhold167 _6502_/Q VGND VGND VPWR VPWR hold167/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold178 _5354_/X VGND VGND VPWR VPWR _6934_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 _6878_/Q VGND VGND VPWR VPWR hold189/X sky130_fd_sc_hd__dlygate4sd3_1
X_7165_ _7183_/CLK _7165_/D fanout500/X VGND VGND VPWR VPWR _7165_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4377_ _4546_/A _4547_/A VGND VGND VPWR VPWR _4657_/A sky130_fd_sc_hd__nor2_2
XFILLER_98_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6116_ _6973_/Q _6009_/X _6030_/X _6997_/Q VGND VGND VPWR VPWR _6116_/X sky130_fd_sc_hd__a22o_1
X_3328_ _3526_/A _3536_/A VGND VGND VPWR VPWR _5484_/A sky130_fd_sc_hd__nor2_4
X_7096_ _7137_/CLK _7096_/D fanout501/X VGND VGND VPWR VPWR _7096_/Q sky130_fd_sc_hd__dfstp_2
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6047_ _5650_/Y _6045_/X _6046_/X _5652_/Y _6071_/A2 VGND VGND VPWR VPWR _7175_/D
+ sky130_fd_sc_hd__a32o_1
X_3259_ hold64/X hold53/X hold72/X VGND VGND VPWR VPWR hold65/A sky130_fd_sc_hd__mux2_1
XTAP_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6949_ _7140_/CLK _6949_/D fanout522/X VGND VGND VPWR VPWR _6949_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_139_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold690 _4220_/X VGND VGND VPWR VPWR _6673_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1390 _7064_/Q VGND VGND VPWR VPWR _5500_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_691 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput206 _3189_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[3] sky130_fd_sc_hd__buf_12
Xoutput217 _3938_/X VGND VGND VPWR VPWR mgmt_gpio_out[13] sky130_fd_sc_hd__buf_12
X_4300_ _4300_/A _5580_/B VGND VGND VPWR VPWR _4305_/S sky130_fd_sc_hd__nand2_2
Xoutput228 _6553_/Q VGND VGND VPWR VPWR mgmt_gpio_out[23] sky130_fd_sc_hd__buf_12
XFILLER_99_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5280_ _5496_/A0 hold811/X _5285_/S VGND VGND VPWR VPWR _5280_/X sky130_fd_sc_hd__mux2_1
Xoutput239 _3924_/X VGND VGND VPWR VPWR mgmt_gpio_out[33] sky130_fd_sc_hd__buf_12
XFILLER_141_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4231_ _6696_/Q _4232_/B VGND VGND VPWR VPWR _6362_/A sky130_fd_sc_hd__nor2_8
XFILLER_141_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4162_ hold273/X hold44/X _4164_/S VGND VGND VPWR VPWR _4162_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4093_ _4093_/A0 _4092_/X _4103_/S VGND VGND VPWR VPWR _4093_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6803_ _7207_/CLK _6803_/D fanout488/X VGND VGND VPWR VPWR _6803_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_169_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4995_ _4995_/A _5036_/B VGND VGND VPWR VPWR _5007_/B sky130_fd_sc_hd__nor2_1
X_6734_ _7211_/CLK _6734_/D fanout489/X VGND VGND VPWR VPWR _6734_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_149_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3946_ _6459_/Q _3946_/B VGND VGND VPWR VPWR _3946_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_28 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6665_ _6764_/CLK _6665_/D _3946_/B VGND VGND VPWR VPWR _6665_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_137_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3877_ _6458_/Q hold12/A _6407_/B VGND VGND VPWR VPWR _3962_/B sky130_fd_sc_hd__o21ai_1
XFILLER_192_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5616_ _6562_/Q _5650_/B VGND VGND VPWR VPWR _5624_/B sky130_fd_sc_hd__nand2_1
XFILLER_176_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6596_ _6759_/CLK _6596_/D fanout489/X VGND VGND VPWR VPWR _6596_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_164_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5547_ _5574_/A0 _5547_/A1 _5552_/S VGND VGND VPWR VPWR _5547_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5478_ _5583_/A0 hold309/X hold79/X VGND VGND VPWR VPWR _5478_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4429_ _4933_/A _4944_/B VGND VGND VPWR VPWR _4836_/A sky130_fd_sc_hd__nor2_1
XFILLER_48_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7148_ _7181_/CLK _7148_/D fanout499/X VGND VGND VPWR VPWR _7148_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout444 _5558_/A0 VGND VGND VPWR VPWR _5534_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout455 _4327_/A1 VGND VGND VPWR VPWR _6395_/A0 sky130_fd_sc_hd__buf_6
Xfanout466 _5212_/C VGND VGND VPWR VPWR _6393_/A0 sky130_fd_sc_hd__buf_6
Xfanout477 _4693_/A VGND VGND VPWR VPWR _4814_/A sky130_fd_sc_hd__buf_6
Xfanout488 fanout491/X VGND VGND VPWR VPWR fanout488/X sky130_fd_sc_hd__buf_6
X_7079_ _7079_/CLK _7079_/D fanout517/X VGND VGND VPWR VPWR _7079_/Q sky130_fd_sc_hd__dfrtp_1
Xfanout499 fanout500/X VGND VGND VPWR VPWR fanout499/X sky130_fd_sc_hd__buf_8
XFILLER_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3800_ _3800_/A _3800_/B VGND VGND VPWR VPWR _6472_/D sky130_fd_sc_hd__nor2_1
XFILLER_178_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4780_ _4780_/A _4981_/C VGND VGND VPWR VPWR _5119_/A sky130_fd_sc_hd__nor2_1
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3731_ _3731_/A _4111_/B VGND VGND VPWR VPWR _5210_/A sky130_fd_sc_hd__nor2_1
XFILLER_159_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_0_csclk _7018_/CLK VGND VGND VPWR VPWR _6764_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_158_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3662_ _3661_/X _3662_/A1 _3917_/A VGND VGND VPWR VPWR _3662_/X sky130_fd_sc_hd__mux2_1
XFILLER_158_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6450_ net499_2/A _6450_/D _6405_/X VGND VGND VPWR VPWR _6450_/Q sky130_fd_sc_hd__dfrtp_1
X_5401_ hold311/X _5569_/A0 _5402_/S VGND VGND VPWR VPWR _5401_/X sky130_fd_sc_hd__mux2_1
X_6381_ _6700_/Q _6381_/A2 _6381_/B1 _6699_/Q VGND VGND VPWR VPWR _6381_/X sky130_fd_sc_hd__a22o_1
X_3593_ _3593_/A _3593_/B _3593_/C _3593_/D VGND VGND VPWR VPWR _3601_/C sky130_fd_sc_hd__or4_1
XFILLER_126_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5332_ _5521_/A0 _5332_/A1 _5339_/S VGND VGND VPWR VPWR _5332_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5263_ _5584_/A0 hold544/X _5267_/S VGND VGND VPWR VPWR _5263_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7002_ _7002_/CLK _7002_/D fanout500/X VGND VGND VPWR VPWR _7002_/Q sky130_fd_sc_hd__dfstp_1
X_4214_ hold387/X _5533_/A1 _4215_/S VGND VGND VPWR VPWR _4214_/X sky130_fd_sc_hd__mux2_1
X_5194_ _6393_/A0 _5194_/A1 _5199_/S VGND VGND VPWR VPWR _5194_/X sky130_fd_sc_hd__mux2_1
X_4145_ hold36/X _4145_/A1 _4146_/S VGND VGND VPWR VPWR _4145_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4076_ hold550/X _4075_/X _4086_/S VGND VGND VPWR VPWR _4076_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4978_ _4870_/B _4783_/Y _5095_/C _5145_/A VGND VGND VPWR VPWR _4979_/D sky130_fd_sc_hd__a211o_1
X_6717_ _7115_/CLK _6717_/D fanout501/X VGND VGND VPWR VPWR _6717_/Q sky130_fd_sc_hd__dfrtp_1
X_3929_ _6560_/Q input77/X _3957_/B VGND VGND VPWR VPWR _3929_/X sky130_fd_sc_hd__mux2_4
XFILLER_20_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6648_ _7187_/CLK _6648_/D VGND VGND VPWR VPWR _6648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6579_ _6579_/CLK _6579_/D _6407_/A VGND VGND VPWR VPWR _6579_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_117_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap408 _6022_/D VGND VGND VPWR VPWR _6323_/B1 sky130_fd_sc_hd__buf_12
XFILLER_171_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap419 _5689_/X VGND VGND VPWR VPWR _5691_/B sky130_fd_sc_hd__buf_12
XFILLER_143_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5950_ _6669_/Q _5677_/X _5688_/X _6610_/Q _5949_/X VGND VGND VPWR VPWR _5957_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_46_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4901_ _5027_/A _4677_/B _4679_/B _4689_/B _4900_/X VGND VGND VPWR VPWR _4905_/A
+ sky130_fd_sc_hd__a41o_1
X_5881_ _6563_/Q _7169_/Q _5880_/X VGND VGND VPWR VPWR _5881_/X sky130_fd_sc_hd__a21o_1
XFILLER_61_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4832_ _4932_/A _4832_/B _4839_/B VGND VGND VPWR VPWR _4843_/B sky130_fd_sc_hd__nor3_1
XANTENNA_190 _3308_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4763_ _4993_/A _4448_/B _4753_/Y _4762_/X VGND VGND VPWR VPWR _4764_/C sky130_fd_sc_hd__a211o_1
XFILLER_159_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6502_ _7139_/CLK _6502_/D fanout518/X VGND VGND VPWR VPWR _6502_/Q sky130_fd_sc_hd__dfrtp_1
X_3714_ _5241_/B _3714_/B VGND VGND VPWR VPWR _5229_/A sky130_fd_sc_hd__nor2_1
X_4694_ _4832_/B _4694_/B VGND VGND VPWR VPWR _4694_/X sky130_fd_sc_hd__or2_1
X_6433_ _6433_/A _6441_/B VGND VGND VPWR VPWR _6433_/X sky130_fd_sc_hd__and2_1
X_3645_ _7028_/Q _3326_/Y _4046_/A _6538_/Q VGND VGND VPWR VPWR _3645_/X sky130_fd_sc_hd__a22o_1
XFILLER_20_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3576_ _6893_/Q _5304_/A _4174_/A _6637_/Q VGND VGND VPWR VPWR _3576_/X sky130_fd_sc_hd__a22o_1
XFILLER_136_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6364_ _6700_/Q _6364_/A2 _6364_/B1 _6699_/Q _6363_/X VGND VGND VPWR VPWR _6364_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5315_ hold9/X _5315_/A1 hold23/X VGND VGND VPWR VPWR hold24/A sky130_fd_sc_hd__mux2_1
X_6295_ _6295_/A1 _6319_/S _6293_/X _6294_/X VGND VGND VPWR VPWR _7185_/D sky130_fd_sc_hd__o22a_1
XFILLER_0_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5246_ hold85/X hold152/X hold14/X VGND VGND VPWR VPWR _5246_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold16 hold16/A VGND VGND VPWR VPWR hold16/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 hold27/A VGND VGND VPWR VPWR hold27/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 hold38/A VGND VGND VPWR VPWR hold38/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 hold49/A VGND VGND VPWR VPWR hold49/X sky130_fd_sc_hd__dlygate4sd3_1
X_5177_ _5177_/A _5177_/B _5176_/X VGND VGND VPWR VPWR _5178_/D sky130_fd_sc_hd__or3b_1
XFILLER_68_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4128_ _5552_/A0 hold755/X _4128_/S VGND VGND VPWR VPWR _4128_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4059_ hold975/X _4058_/X _4069_/S VGND VGND VPWR VPWR _4059_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold508 _6945_/Q VGND VGND VPWR VPWR hold508/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold519 _5285_/X VGND VGND VPWR VPWR _6873_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3430_ input57/X _5232_/A hold69/A _7140_/Q _3418_/X VGND VGND VPWR VPWR _3431_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3361_ _6481_/Q _3966_/A hold30/A _6881_/Q _3360_/X VGND VGND VPWR VPWR _3373_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_112_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5100_ _5100_/A _5140_/A _5142_/B _5100_/D VGND VGND VPWR VPWR _5101_/D sky130_fd_sc_hd__or4_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6080_ _6500_/Q _6323_/A2 _5988_/X _7052_/Q VGND VGND VPWR VPWR _6080_/X sky130_fd_sc_hd__a22o_1
X_3292_ _3495_/A hold29/X VGND VGND VPWR VPWR _5502_/A sky130_fd_sc_hd__nor2_8
XFILLER_112_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5031_ _5031_/A _5031_/B _5031_/C VGND VGND VPWR VPWR _5071_/C sky130_fd_sc_hd__or3_2
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1208 _5370_/X VGND VGND VPWR VPWR _6948_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1219 _4175_/X VGND VGND VPWR VPWR _6634_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6982_ _7070_/CLK _6982_/D fanout510/X VGND VGND VPWR VPWR _6982_/Q sky130_fd_sc_hd__dfrtp_2
X_5933_ _6704_/Q _5659_/X _5699_/X _6539_/Q VGND VGND VPWR VPWR _5933_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_33_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7134_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_178_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5864_ _6721_/Q _5702_/X _5703_/X _6601_/Q _5863_/X VGND VGND VPWR VPWR _5869_/B
+ sky130_fd_sc_hd__a221o_1
X_4815_ _4815_/A _4987_/C _4815_/C _4814_/X VGND VGND VPWR VPWR _4817_/C sky130_fd_sc_hd__or4b_1
XFILLER_166_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5795_ _5795_/A0 _5794_/X _6319_/S VGND VGND VPWR VPWR _7166_/D sky130_fd_sc_hd__mux2_1
XFILLER_119_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_48_csclk _6931_/CLK VGND VGND VPWR VPWR _6923_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_119_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4746_ _4981_/B _4994_/A VGND VGND VPWR VPWR _4746_/Y sky130_fd_sc_hd__nor2_1
XFILLER_193_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4677_ _5023_/A _4677_/B VGND VGND VPWR VPWR _5054_/B sky130_fd_sc_hd__or2_1
XFILLER_134_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6416_ _6433_/A _6441_/B VGND VGND VPWR VPWR _6416_/X sky130_fd_sc_hd__and2_1
X_3628_ _6672_/Q _4216_/A _4159_/A _6623_/Q _3609_/X VGND VGND VPWR VPWR _3632_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6347_ _6347_/A1 _3888_/Y _6346_/Y _6345_/X VGND VGND VPWR VPWR _7188_/D sky130_fd_sc_hd__a31o_1
XFILLER_0_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3559_ _6501_/Q _3778_/A2 _4324_/A _6769_/Q VGND VGND VPWR VPWR _3559_/X sky130_fd_sc_hd__a22o_1
XFILLER_88_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6278_ _6773_/Q _6002_/Y _6007_/Y _6758_/Q _6277_/X VGND VGND VPWR VPWR _6280_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput106 wb_adr_i[16] VGND VGND VPWR VPWR _4337_/B sky130_fd_sc_hd__clkbuf_1
Xinput117 wb_adr_i[26] VGND VGND VPWR VPWR input117/X sky130_fd_sc_hd__clkbuf_1
Xinput128 wb_adr_i[7] VGND VGND VPWR VPWR _4935_/A sky130_fd_sc_hd__buf_6
X_5229_ _5229_/A _6392_/B VGND VGND VPWR VPWR _5231_/S sky130_fd_sc_hd__nand2_1
XFILLER_76_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput139 wb_dat_i[16] VGND VGND VPWR VPWR _6363_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_56_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_90 _6461_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_3_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_121_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4600_ _4367_/B _5106_/A _4574_/Y _4599_/X _5148_/A VGND VGND VPWR VPWR _4600_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_30_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5580_ hold69/X _5580_/B VGND VGND VPWR VPWR hold70/A sky130_fd_sc_hd__nand2_8
XFILLER_30_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4531_ _4846_/C _4369_/B _4464_/Y _5050_/A _4530_/X VGND VGND VPWR VPWR _4531_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_129_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold305 _7028_/Q VGND VGND VPWR VPWR hold305/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold316 _5387_/X VGND VGND VPWR VPWR _6963_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4462_ _4605_/A _4462_/B VGND VGND VPWR VPWR _4462_/Y sky130_fd_sc_hd__nor2_1
Xhold327 _6737_/Q VGND VGND VPWR VPWR hold327/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 _5378_/X VGND VGND VPWR VPWR _6955_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6201_ _7081_/Q _5994_/X _5998_/Y _7017_/Q _6198_/X VGND VGND VPWR VPWR _6201_/X
+ sky130_fd_sc_hd__a221o_1
Xhold349 hold349/A VGND VGND VPWR VPWR hold349/X sky130_fd_sc_hd__dlygate4sd3_1
X_3413_ _7174_/Q _6816_/Q _6818_/Q VGND VGND VPWR VPWR _3413_/X sky130_fd_sc_hd__mux2_8
XFILLER_144_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7181_ _7181_/CLK _7181_/D fanout505/X VGND VGND VPWR VPWR _7181_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_171_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4393_ _4351_/A _4351_/B _4391_/Y VGND VGND VPWR VPWR _4932_/A sky130_fd_sc_hd__a21o_4
XFILLER_98_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3344_ _3731_/A _3546_/B VGND VGND VPWR VPWR _3983_/A sky130_fd_sc_hd__nor2_8
X_6132_ _6974_/Q _6009_/X _6206_/B1 _6982_/Q _6131_/X VGND VGND VPWR VPWR _6132_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3275_ _3546_/A _5212_/B VGND VGND VPWR VPWR _5232_/A sky130_fd_sc_hd__nor2_8
X_6063_ _6947_/Q _6024_/A _6040_/X _7043_/Q VGND VGND VPWR VPWR _6063_/X sky130_fd_sc_hd__a22o_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1005 _6959_/Q VGND VGND VPWR VPWR _5382_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1016 _5283_/X VGND VGND VPWR VPWR _6871_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1027 _7132_/Q VGND VGND VPWR VPWR _5577_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5014_ _4400_/B _4718_/B _5013_/A VGND VGND VPWR VPWR _5015_/C sky130_fd_sc_hd__a21oi_1
Xhold1038 _5271_/X VGND VGND VPWR VPWR _6860_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 _6946_/Q VGND VGND VPWR VPWR _5368_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6965_ _7140_/CLK _6965_/D fanout522/X VGND VGND VPWR VPWR _6965_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_53_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5916_ _6713_/Q _5938_/B VGND VGND VPWR VPWR _5916_/X sky130_fd_sc_hd__or2_1
XFILLER_81_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6896_ _6969_/CLK _6896_/D fanout506/X VGND VGND VPWR VPWR _6896_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_22_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5847_ _5847_/A _5847_/B _5847_/C _5847_/D VGND VGND VPWR VPWR _5847_/X sky130_fd_sc_hd__or4_1
XFILLER_21_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5778_ _6926_/Q _5955_/A2 _5700_/X _7030_/Q _5777_/X VGND VGND VPWR VPWR _5785_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_154_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4729_ _4981_/B _5094_/A VGND VGND VPWR VPWR _4729_/Y sky130_fd_sc_hd__nand2_1
XFILLER_135_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold850 _7059_/Q VGND VGND VPWR VPWR hold850/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold861 _5551_/X VGND VGND VPWR VPWR _7109_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold872 _6772_/Q VGND VGND VPWR VPWR hold872/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold883 _5464_/X VGND VGND VPWR VPWR _7032_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold894 _6671_/Q VGND VGND VPWR VPWR hold894/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1550 _6542_/Q VGND VGND VPWR VPWR _3912_/B1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1561 _7185_/Q VGND VGND VPWR VPWR _6295_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1572 _6578_/Q VGND VGND VPWR VPWR hold799/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1583 hold64/A VGND VGND VPWR VPWR _3828_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1594 _6471_/Q VGND VGND VPWR VPWR _3801_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6750_ _6963_/CLK _6750_/D fanout509/X VGND VGND VPWR VPWR _6750_/Q sky130_fd_sc_hd__dfrtp_1
X_3962_ _6700_/Q _3962_/B VGND VGND VPWR VPWR _6692_/D sky130_fd_sc_hd__and2_1
XFILLER_189_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5701_ _7050_/Q _5699_/X _5700_/X _7026_/Q _5698_/X VGND VGND VPWR VPWR _5708_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_188_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6681_ _6683_/CLK _6681_/D fanout511/X VGND VGND VPWR VPWR _6681_/Q sky130_fd_sc_hd__dfrtp_4
X_3893_ _6699_/Q _3876_/X _3893_/B1 VGND VGND VPWR VPWR _6699_/D sky130_fd_sc_hd__a21o_1
XFILLER_31_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5632_ _5632_/A1 _5637_/B _5631_/Y VGND VGND VPWR VPWR _7155_/D sky130_fd_sc_hd__a21oi_1
XFILLER_129_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5563_ _5581_/A0 _5563_/A1 _5570_/S VGND VGND VPWR VPWR _5563_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4514_ _4516_/B _5001_/B VGND VGND VPWR VPWR _4863_/A sky130_fd_sc_hd__nand2_1
Xhold102 _5239_/X VGND VGND VPWR VPWR _6832_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold113 hold113/A VGND VGND VPWR VPWR _5385_/B sky130_fd_sc_hd__buf_8
X_5494_ _5581_/A0 _5494_/A1 _5501_/S VGND VGND VPWR VPWR _5494_/X sky130_fd_sc_hd__mux2_1
Xhold124 _5248_/X VGND VGND VPWR VPWR _6840_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 _6680_/Q VGND VGND VPWR VPWR _3981_/S sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold146 _6724_/Q VGND VGND VPWR VPWR hold146/X sky130_fd_sc_hd__dlygate4sd3_1
X_4445_ _4445_/A _4724_/B VGND VGND VPWR VPWR _4872_/A sky130_fd_sc_hd__or2_4
Xhold157 _5255_/X VGND VGND VPWR VPWR _6846_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 _4006_/X VGND VGND VPWR VPWR _6502_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold179 hold179/A VGND VGND VPWR VPWR hold179/X sky130_fd_sc_hd__dlygate4sd3_1
X_7164_ _7183_/CLK _7164_/D fanout500/X VGND VGND VPWR VPWR _7164_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_144_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4376_ _4570_/D _4376_/B VGND VGND VPWR VPWR _5023_/A sky130_fd_sc_hd__nand2_8
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6115_ _6501_/Q _6323_/A2 wire412/X _6917_/Q VGND VGND VPWR VPWR _6115_/X sky130_fd_sc_hd__a22o_1
X_3327_ _5212_/B _3534_/A VGND VGND VPWR VPWR _5448_/A sky130_fd_sc_hd__nor2_8
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7095_ _7137_/CLK _7095_/D fanout501/X VGND VGND VPWR VPWR _7095_/Q sky130_fd_sc_hd__dfstp_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6046_ _6842_/Q _6046_/B VGND VGND VPWR VPWR _6046_/X sky130_fd_sc_hd__or2_1
X_3258_ hold73/X _3258_/A1 _3971_/S VGND VGND VPWR VPWR hold74/A sky130_fd_sc_hd__mux2_2
XFILLER_39_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3189_ _6869_/Q VGND VGND VPWR VPWR _3189_/Y sky130_fd_sc_hd__inv_2
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6948_ _7135_/CLK _6948_/D fanout526/X VGND VGND VPWR VPWR _6948_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_169_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6879_ _7126_/CLK _6879_/D fanout523/X VGND VGND VPWR VPWR _6879_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_139_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold680 _5508_/X VGND VGND VPWR VPWR _7071_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold691 _7130_/Q VGND VGND VPWR VPWR hold691/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1380 _5582_/X VGND VGND VPWR VPWR hold6/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1391 _7077_/Q VGND VGND VPWR VPWR _5515_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput207 _3230_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[4] sky130_fd_sc_hd__buf_12
XFILLER_99_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput218 _3937_/X VGND VGND VPWR VPWR mgmt_gpio_out[14] sky130_fd_sc_hd__clkbuf_1
XFILLER_153_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput229 _6826_/Q VGND VGND VPWR VPWR mgmt_gpio_out[24] sky130_fd_sc_hd__buf_12
XFILLER_99_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4230_ _6692_/Q _6693_/Q _6695_/Q _6694_/Q VGND VGND VPWR VPWR _4230_/X sky130_fd_sc_hd__or4_1
XFILLER_141_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4161_ hold333/X _5459_/A0 _4164_/S VGND VGND VPWR VPWR _4161_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4092_ hold868/X _5496_/A0 _4102_/S VGND VGND VPWR VPWR _4092_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6802_ _7207_/CLK _6802_/D fanout488/X VGND VGND VPWR VPWR _6802_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_51_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4994_ _4994_/A _5036_/B VGND VGND VPWR VPWR _5008_/A sky130_fd_sc_hd__nor2_1
XFILLER_90_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6733_ _7211_/CLK _6733_/D fanout489/X VGND VGND VPWR VPWR _6733_/Q sky130_fd_sc_hd__dfstp_2
X_3945_ input83/X _3945_/A1 _6459_/Q VGND VGND VPWR VPWR _3945_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6664_ _6664_/CLK _6664_/D _3946_/B VGND VGND VPWR VPWR _6664_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_31_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3876_ _6458_/Q hold12/A _6407_/B VGND VGND VPWR VPWR _3876_/X sky130_fd_sc_hd__o21a_1
XFILLER_177_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5615_ _5615_/A _6564_/Q VGND VGND VPWR VPWR _5643_/A sky130_fd_sc_hd__nor2_1
XFILLER_136_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6595_ _7033_/CLK _6595_/D fanout504/X VGND VGND VPWR VPWR _6595_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5546_ _5573_/A0 hold880/X _5552_/S VGND VGND VPWR VPWR _5546_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5477_ _5573_/A0 hold844/X hold79/X VGND VGND VPWR VPWR _5477_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4428_ _4605_/A _4428_/B VGND VGND VPWR VPWR _4944_/B sky130_fd_sc_hd__nand2_1
Xclkbuf_2_3__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR net499_2/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_48_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7147_ _7181_/CLK _7147_/D fanout502/X VGND VGND VPWR VPWR _7147_/Q sky130_fd_sc_hd__dfrtp_1
Xfanout434 hold40/X VGND VGND VPWR VPWR _5552_/A0 sky130_fd_sc_hd__buf_8
Xfanout445 hold84/X VGND VGND VPWR VPWR _5558_/A0 sky130_fd_sc_hd__buf_6
XFILLER_101_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4359_ _4610_/A _4781_/A VGND VGND VPWR VPWR _4428_/B sky130_fd_sc_hd__xnor2_2
XFILLER_86_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout456 _5583_/A0 VGND VGND VPWR VPWR _4327_/A1 sky130_fd_sc_hd__buf_4
Xfanout467 _5476_/A0 VGND VGND VPWR VPWR _5212_/C sky130_fd_sc_hd__clkbuf_8
Xfanout489 fanout491/X VGND VGND VPWR VPWR fanout489/X sky130_fd_sc_hd__buf_4
X_7078_ _7078_/CLK _7078_/D fanout515/X VGND VGND VPWR VPWR _7078_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_100_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6029_ _6040_/B _6029_/B _6029_/C _6029_/D VGND VGND VPWR VPWR _6046_/B sky130_fd_sc_hd__or4_4
XFILLER_100_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3730_ _6460_/Q _6445_/Q _6811_/Q VGND VGND VPWR VPWR _3730_/X sky130_fd_sc_hd__or3_4
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3661_ _3660_/X _6784_/Q _3791_/A VGND VGND VPWR VPWR _3661_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5400_ _5400_/A0 _5586_/A0 _5402_/S VGND VGND VPWR VPWR _5400_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6380_ _6379_/X _6380_/A1 _6386_/S VGND VGND VPWR VPWR _7202_/D sky130_fd_sc_hd__mux2_1
X_3592_ input6/X _3295_/Y _3304_/Y input29/X _3554_/X VGND VGND VPWR VPWR _3593_/D
+ sky130_fd_sc_hd__a221o_2
XFILLER_127_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5331_ _5331_/A _5571_/B VGND VGND VPWR VPWR _5339_/S sky130_fd_sc_hd__nand2_8
XFILLER_161_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5262_ _5574_/A0 _5262_/A1 _5267_/S VGND VGND VPWR VPWR _5262_/X sky130_fd_sc_hd__mux2_1
X_7001_ _7102_/CLK _7001_/D fanout503/X VGND VGND VPWR VPWR _7001_/Q sky130_fd_sc_hd__dfrtp_4
X_4213_ hold856/X _4327_/A1 _4215_/S VGND VGND VPWR VPWR _4213_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5193_ _5193_/A _6392_/B VGND VGND VPWR VPWR _5199_/S sky130_fd_sc_hd__nand2_2
XFILLER_68_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4144_ hold44/X hold241/X _4146_/S VGND VGND VPWR VPWR _4144_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4075_ hold329/X _5583_/A0 _4085_/S VGND VGND VPWR VPWR _4075_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_4_0_csclk clkbuf_3_5_0_csclk/A VGND VGND VPWR VPWR _6820_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_64_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4977_ _5094_/B _4971_/Y _4976_/X VGND VGND VPWR VPWR _5145_/A sky130_fd_sc_hd__o21ai_1
X_6716_ _7074_/CLK _6716_/D fanout501/X VGND VGND VPWR VPWR _6716_/Q sky130_fd_sc_hd__dfrtp_1
X_3928_ _6566_/Q _3872_/C _6462_/Q VGND VGND VPWR VPWR _3928_/X sky130_fd_sc_hd__mux2_1
XFILLER_165_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6647_ _7187_/CLK _6647_/D VGND VGND VPWR VPWR _6647_/Q sky130_fd_sc_hd__dfxtp_1
X_3859_ input58/X _3856_/B _3853_/B _3859_/B2 _3858_/X VGND VGND VPWR VPWR _6453_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_165_746 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6578_ _6579_/CLK _6578_/D _6407_/A VGND VGND VPWR VPWR _6578_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_124_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5529_ _5529_/A _6392_/B VGND VGND VPWR VPWR _5534_/S sky130_fd_sc_hd__and2_2
XFILLER_3_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_74 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap409 _6016_/X VGND VGND VPWR VPWR _6024_/D sky130_fd_sc_hd__buf_12
XFILLER_40_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4900_ _5023_/B _5016_/A VGND VGND VPWR VPWR _4900_/X sky130_fd_sc_hd__and2_1
XFILLER_46_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5880_ _6596_/Q _5691_/Y _5869_/X _5879_/X _6318_/S VGND VGND VPWR VPWR _5880_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_73_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4831_ _5023_/B _4689_/B _4524_/Y VGND VGND VPWR VPWR _5162_/A sky130_fd_sc_hd__o21ai_1
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_180 _3927_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_191 _4083_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4762_ _4993_/A _4759_/B _4984_/B _4761_/X VGND VGND VPWR VPWR _4762_/X sky130_fd_sc_hd__a211o_1
XFILLER_159_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6501_ _7108_/CLK _6501_/D fanout523/X VGND VGND VPWR VPWR _6501_/Q sky130_fd_sc_hd__dfrtp_4
X_3713_ _6859_/Q _5268_/A _3318_/Y _6883_/Q _3712_/X VGND VGND VPWR VPWR _3721_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4693_ _4693_/A _4832_/B _4784_/A VGND VGND VPWR VPWR _4698_/B sky130_fd_sc_hd__or3_1
X_6432_ _6432_/A _6441_/B VGND VGND VPWR VPWR _6432_/X sky130_fd_sc_hd__and2_1
X_3644_ _6800_/Q _5193_/A _4016_/A _6513_/Q _3643_/X VGND VGND VPWR VPWR _3651_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_134_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6363_ _6698_/Q _6363_/A2 _6363_/B1 _6390_/A2 VGND VGND VPWR VPWR _6363_/X sky130_fd_sc_hd__a22o_1
X_3575_ _6853_/Q _5259_/A _4141_/A _6609_/Q _3574_/X VGND VGND VPWR VPWR _3582_/A
+ sky130_fd_sc_hd__a221o_1
X_5314_ _5581_/A0 _5314_/A1 hold23/X VGND VGND VPWR VPWR _5314_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6294_ _7184_/Q _5592_/Y _5650_/Y VGND VGND VPWR VPWR _6294_/X sky130_fd_sc_hd__o21ba_1
XFILLER_114_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5245_ hold36/X hold197/X hold14/X VGND VGND VPWR VPWR _5245_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold17 hold17/A VGND VGND VPWR VPWR hold17/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold28 hold28/A VGND VGND VPWR VPWR hold28/X sky130_fd_sc_hd__buf_6
XFILLER_102_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5176_ _4659_/B _5027_/B _5108_/B _4679_/B VGND VGND VPWR VPWR _5176_/X sky130_fd_sc_hd__o22a_1
XFILLER_152_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold39 hold39/A VGND VGND VPWR VPWR hold39/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4127_ _5569_/A0 hold227/X _4128_/S VGND VGND VPWR VPWR _4127_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4058_ hold783/X _5496_/A0 _4068_/S VGND VGND VPWR VPWR _4058_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_5_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A VGND VGND VPWR VPWR _7196_/CLK sky130_fd_sc_hd__clkbuf_8
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_726 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold509 _5366_/X VGND VGND VPWR VPWR _6945_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_524 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3360_ _7102_/Q _5535_/A _3357_/X _3359_/X VGND VGND VPWR VPWR _3360_/X sky130_fd_sc_hd__a211o_1
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3291_ _3303_/A hold28/X VGND VGND VPWR VPWR hold29/A sky130_fd_sc_hd__nand2_8
XFILLER_151_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5030_ _5030_/A _5073_/B _5079_/B _5029_/X VGND VGND VPWR VPWR _5030_/X sky130_fd_sc_hd__or4b_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1209 hold1610/X VGND VGND VPWR VPWR _4105_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6981_ _7140_/CLK _6981_/D fanout522/X VGND VGND VPWR VPWR _6981_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_19_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5932_ _6734_/Q _5697_/X _5931_/X VGND VGND VPWR VPWR _5935_/C sky130_fd_sc_hd__a21o_1
XFILLER_80_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5863_ _6670_/Q _5955_/A2 _5688_/X _6606_/Q VGND VGND VPWR VPWR _5863_/X sky130_fd_sc_hd__a22o_1
XFILLER_178_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4814_ _4814_/A _4814_/B _4814_/C VGND VGND VPWR VPWR _4814_/X sky130_fd_sc_hd__or3_1
XFILLER_21_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5794_ _5650_/A _5794_/A2 _5793_/X VGND VGND VPWR VPWR _5794_/X sky130_fd_sc_hd__a21o_1
XFILLER_119_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4745_ _4745_/A _4871_/A VGND VGND VPWR VPWR _4875_/B sky130_fd_sc_hd__nor2_1
XFILLER_193_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4676_ _4646_/A _4683_/B _4692_/B _4675_/A VGND VGND VPWR VPWR _4676_/X sky130_fd_sc_hd__o22a_1
XFILLER_107_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6415_ _6426_/A _6441_/B VGND VGND VPWR VPWR _6415_/X sky130_fd_sc_hd__and2_1
X_3627_ _3627_/A _3627_/B _3627_/C _3627_/D VGND VGND VPWR VPWR _3633_/C sky130_fd_sc_hd__or4_1
XFILLER_134_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6346_ _6346_/A _6697_/Q VGND VGND VPWR VPWR _6346_/Y sky130_fd_sc_hd__nand2_1
X_3558_ _6925_/Q _5340_/A _4252_/A _6709_/Q VGND VGND VPWR VPWR _3583_/A sky130_fd_sc_hd__a22o_1
XFILLER_1_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6277_ _6733_/Q _5997_/Y _6015_/X _6662_/Q VGND VGND VPWR VPWR _6277_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3489_ _3530_/B _4120_/B VGND VGND VPWR VPWR _4258_/A sky130_fd_sc_hd__nor2_4
Xinput107 wb_adr_i[17] VGND VGND VPWR VPWR _4337_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_76_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput118 wb_adr_i[27] VGND VGND VPWR VPWR _3885_/A sky130_fd_sc_hd__clkbuf_1
X_5228_ hold979/X _5581_/A0 _5228_/S VGND VGND VPWR VPWR _5228_/X sky130_fd_sc_hd__mux2_1
Xinput129 wb_adr_i[8] VGND VGND VPWR VPWR _4339_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_56_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5159_ _5159_/A _5159_/B _5159_/C VGND VGND VPWR VPWR _5160_/C sky130_fd_sc_hd__nand3_1
XFILLER_84_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_2_1_0_csclk clkbuf_2_1_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_3_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_80 _6169_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_91 _6461_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4530_ _4530_/A _4530_/B _4530_/C _4530_/D VGND VGND VPWR VPWR _4530_/X sky130_fd_sc_hd__and4_1
XFILLER_7_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold306 _5460_/X VGND VGND VPWR VPWR _7028_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4461_ _5076_/A _4461_/B VGND VGND VPWR VPWR _5126_/A sky130_fd_sc_hd__nor2_1
Xhold317 _6988_/Q VGND VGND VPWR VPWR hold317/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold328 _4290_/X VGND VGND VPWR VPWR _6737_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6200_ _6905_/Q _6022_/B _6025_/D _6969_/Q VGND VGND VPWR VPWR _6216_/B sky130_fd_sc_hd__a22o_1
Xhold339 _6907_/Q VGND VGND VPWR VPWR hold339/X sky130_fd_sc_hd__dlygate4sd3_1
X_3412_ _3411_/X _3412_/A1 _3917_/A VGND VGND VPWR VPWR _6789_/D sky130_fd_sc_hd__mux2_1
X_7180_ _7181_/CLK _7180_/D fanout506/X VGND VGND VPWR VPWR _7180_/Q sky130_fd_sc_hd__dfrtp_1
X_4392_ _4390_/C _4390_/D _4467_/A _4674_/A VGND VGND VPWR VPWR _4560_/A sky130_fd_sc_hd__a31o_2
XFILLER_171_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6131_ _6958_/Q _6336_/A2 _6205_/B1 _7062_/Q VGND VGND VPWR VPWR _6131_/X sky130_fd_sc_hd__a22o_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3343_ _3528_/A _3546_/B VGND VGND VPWR VPWR _5322_/A sky130_fd_sc_hd__nor2_8
XFILLER_97_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6062_ _6923_/Q _6340_/A2 wire394/X _6891_/Q _6061_/X VGND VGND VPWR VPWR _6068_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3274_ hold28/X hold67/X VGND VGND VPWR VPWR _5212_/B sky130_fd_sc_hd__nand2_8
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1006 _5382_/X VGND VGND VPWR VPWR _6959_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1017 _6932_/Q VGND VGND VPWR VPWR _5352_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ _5013_/A _5076_/B VGND VGND VPWR VPWR _5013_/X sky130_fd_sc_hd__or2_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1028 _5577_/X VGND VGND VPWR VPWR _7132_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1039 hold1562/X VGND VGND VPWR VPWR _4074_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6964_ _7075_/CLK _6964_/D fanout514/X VGND VGND VPWR VPWR _6964_/Q sky130_fd_sc_hd__dfrtp_2
X_5915_ _6688_/Q _5666_/X _5697_/X _6733_/Q _5914_/X VGND VGND VPWR VPWR _5923_/A
+ sky130_fd_sc_hd__a221o_1
X_6895_ _7079_/CLK _6895_/D fanout516/X VGND VGND VPWR VPWR _6895_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5846_ _6889_/Q _5846_/A2 _5666_/X _6953_/Q _5845_/X VGND VGND VPWR VPWR _5847_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_42_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5777_ _7038_/Q _5696_/X _5697_/X _6990_/Q VGND VGND VPWR VPWR _5777_/X sky130_fd_sc_hd__a22o_1
X_4728_ _4759_/A _4870_/B VGND VGND VPWR VPWR _4728_/Y sky130_fd_sc_hd__nor2_1
XFILLER_147_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4659_ _5023_/A _4659_/B VGND VGND VPWR VPWR _5065_/B sky130_fd_sc_hd__nor2_1
XFILLER_162_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold840 _6571_/Q VGND VGND VPWR VPWR hold840/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold851 _5495_/X VGND VGND VPWR VPWR _7059_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_107_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold862 _7083_/Q VGND VGND VPWR VPWR hold862/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold873 _4332_/X VGND VGND VPWR VPWR _6772_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold884 _6960_/Q VGND VGND VPWR VPWR hold884/X sky130_fd_sc_hd__dlygate4sd3_1
X_6329_ _6664_/Q _6024_/C _6329_/B1 _6520_/Q VGND VGND VPWR VPWR _6329_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold895 _4218_/X VGND VGND VPWR VPWR _6671_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_107_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1540 _7172_/Q VGND VGND VPWR VPWR _5926_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1551 _7155_/Q VGND VGND VPWR VPWR _5632_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1562 _6555_/Q VGND VGND VPWR VPWR hold1562/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1573 _6579_/Q VGND VGND VPWR VPWR hold173/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1584 _7187_/Q VGND VGND VPWR VPWR _6344_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_177_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1595 _6593_/Q VGND VGND VPWR VPWR hold193/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_32_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7126_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_79_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_47_csclk _6931_/CLK VGND VGND VPWR VPWR _7128_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_36_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3961_ _6825_/Q _3961_/B VGND VGND VPWR VPWR _3961_/X sky130_fd_sc_hd__and2_2
XFILLER_189_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5700_ _7152_/Q _5706_/B _5700_/C VGND VGND VPWR VPWR _5700_/X sky130_fd_sc_hd__and3_4
XFILLER_50_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6680_ _7200_/CLK _6680_/D _6348_/B VGND VGND VPWR VPWR _6680_/Q sky130_fd_sc_hd__dfrtp_4
X_3892_ _6698_/Q _3876_/X _3892_/B1 VGND VGND VPWR VPWR _6698_/D sky130_fd_sc_hd__a21o_1
XFILLER_176_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5631_ _7155_/Q _5624_/B _5637_/B VGND VGND VPWR VPWR _5631_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_148_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5562_ _5562_/A _5571_/B VGND VGND VPWR VPWR _5562_/Y sky130_fd_sc_hd__nand2_4
XFILLER_129_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4513_ _4516_/B _4657_/C VGND VGND VPWR VPWR _4515_/C sky130_fd_sc_hd__nand2_1
XFILLER_191_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold103 _6467_/Q VGND VGND VPWR VPWR _3248_/A sky130_fd_sc_hd__dlygate4sd3_1
X_5493_ _5493_/A _5571_/B VGND VGND VPWR VPWR _5493_/Y sky130_fd_sc_hd__nand2_8
Xhold114 _5313_/B VGND VGND VPWR VPWR _5571_/B sky130_fd_sc_hd__buf_12
Xhold125 _6450_/Q VGND VGND VPWR VPWR hold125/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4444_ _4434_/B _4444_/B VGND VGND VPWR VPWR _4724_/B sky130_fd_sc_hd__nand2b_2
Xhold136 _3971_/S VGND VGND VPWR VPWR _3967_/S sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 _4274_/X VGND VGND VPWR VPWR _6724_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 _7200_/Q VGND VGND VPWR VPWR hold158/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold169 _6619_/Q VGND VGND VPWR VPWR hold169/X sky130_fd_sc_hd__dlygate4sd3_1
X_7163_ _7183_/CLK _7163_/D fanout508/X VGND VGND VPWR VPWR _7163_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_113_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4375_ _4846_/A _4846_/B _4570_/B VGND VGND VPWR VPWR _4951_/B sky130_fd_sc_hd__nor3b_2
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6114_ _6925_/Q _6027_/B wire394/X _6893_/Q _6113_/X VGND VGND VPWR VPWR _6119_/C
+ sky130_fd_sc_hd__a221o_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3326_ _5241_/B _3534_/A VGND VGND VPWR VPWR _3326_/Y sky130_fd_sc_hd__nor2_8
XFILLER_112_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7094_ _7094_/CLK _7094_/D fanout494/X VGND VGND VPWR VPWR _7094_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6045_ _6045_/A _6045_/B _6045_/C VGND VGND VPWR VPWR _6045_/X sky130_fd_sc_hd__or3_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3257_ hold16/X hold64/X hold72/X VGND VGND VPWR VPWR hold73/A sky130_fd_sc_hd__mux2_1
XTAP_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3188_ _3188_/A VGND VGND VPWR VPWR _6346_/A sky130_fd_sc_hd__inv_2
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6947_ _7043_/CLK _6947_/D fanout514/X VGND VGND VPWR VPWR _6947_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_41_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6878_ _7135_/CLK _6878_/D fanout519/X VGND VGND VPWR VPWR _6878_/Q sky130_fd_sc_hd__dfrtp_2
X_5829_ _6920_/Q _5677_/X _5691_/B _5828_/X VGND VGND VPWR VPWR _5829_/X sky130_fd_sc_hd__a22o_1
XFILLER_139_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold670 _4164_/X VGND VGND VPWR VPWR _6625_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold681 _7010_/Q VGND VGND VPWR VPWR hold681/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 _5575_/X VGND VGND VPWR VPWR _7130_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1370 _6585_/Q VGND VGND VPWR VPWR _4117_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1381 _6822_/Q VGND VGND VPWR VPWR _5227_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1392 _7201_/Q VGND VGND VPWR VPWR _3975_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput208 _3229_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[5] sky130_fd_sc_hd__buf_12
XFILLER_154_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput219 _3936_/X VGND VGND VPWR VPWR mgmt_gpio_out[15] sky130_fd_sc_hd__clkbuf_1
XFILLER_5_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4160_ _4160_/A0 _5521_/A0 _4164_/S VGND VGND VPWR VPWR _4160_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4091_ hold129/X _4090_/X _4103_/S VGND VGND VPWR VPWR _4091_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6801_ _7207_/CLK _6801_/D fanout488/X VGND VGND VPWR VPWR _6801_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_90_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4993_ _4993_/A _4993_/B VGND VGND VPWR VPWR _5036_/B sky130_fd_sc_hd__nor2_4
XFILLER_23_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6732_ _7211_/CLK _6732_/D fanout489/X VGND VGND VPWR VPWR _6732_/Q sky130_fd_sc_hd__dfrtp_2
X_3944_ _6460_/Q _3946_/B VGND VGND VPWR VPWR _3944_/Y sky130_fd_sc_hd__nor2_1
X_6663_ _6664_/CLK _6663_/D fanout485/X VGND VGND VPWR VPWR _6663_/Q sky130_fd_sc_hd__dfrtp_4
X_3875_ _7160_/Q _6813_/Q _6818_/Q VGND VGND VPWR VPWR _5592_/B sky130_fd_sc_hd__mux2_4
XFILLER_139_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5614_ _7149_/Q _7148_/Q VGND VGND VPWR VPWR _5706_/B sky130_fd_sc_hd__and2_2
X_6594_ _6664_/CLK _6594_/D _6426_/A VGND VGND VPWR VPWR _6594_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_164_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5545_ _5581_/A0 _5545_/A1 _5552_/S VGND VGND VPWR VPWR _5545_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_0_0_csclk clkbuf_3_1_0_csclk/A VGND VGND VPWR VPWR _6753_/CLK sky130_fd_sc_hd__clkbuf_8
X_5476_ _5476_/A0 _5476_/A1 hold79/X VGND VGND VPWR VPWR _5476_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7215_ _7215_/A VGND VGND VPWR VPWR _7215_/X sky130_fd_sc_hd__buf_2
X_4427_ _4354_/A _4354_/B _4355_/Y _4350_/B VGND VGND VPWR VPWR _4933_/A sky130_fd_sc_hd__a211o_2
XFILLER_160_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7146_ _7181_/CLK _7146_/D fanout502/X VGND VGND VPWR VPWR _7146_/Q sky130_fd_sc_hd__dfrtp_1
Xfanout424 _4718_/B VGND VGND VPWR VPWR _5076_/B sky130_fd_sc_hd__buf_6
X_4358_ _4621_/B _4781_/A VGND VGND VPWR VPWR _4360_/B sky130_fd_sc_hd__and2_1
Xfanout435 hold40/X VGND VGND VPWR VPWR _5579_/A0 sky130_fd_sc_hd__buf_6
Xfanout446 hold85/X VGND VGND VPWR VPWR _5549_/A0 sky130_fd_sc_hd__buf_6
XFILLER_58_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout457 hold43/X VGND VGND VPWR VPWR _5583_/A0 sky130_fd_sc_hd__buf_8
X_3309_ hold48/X hold18/X _3301_/C VGND VGND VPWR VPWR hold49/A sky130_fd_sc_hd__or3b_4
Xfanout468 _5536_/A1 VGND VGND VPWR VPWR _5476_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_100_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7077_ _7110_/CLK _7077_/D fanout506/X VGND VGND VPWR VPWR _7077_/Q sky130_fd_sc_hd__dfrtp_4
X_4289_ _5521_/A0 _4289_/A1 _4293_/S VGND VGND VPWR VPWR _4289_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6028_ _6040_/B _6029_/B _6029_/C _6029_/D VGND VGND VPWR VPWR _6028_/Y sky130_fd_sc_hd__nor4_1
XFILLER_39_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3660_ _3660_/A _3660_/B _3660_/C VGND VGND VPWR VPWR _3660_/X sky130_fd_sc_hd__or3_4
X_3591_ _6477_/Q _3966_/A _3992_/A _6493_/Q _3560_/X VGND VGND VPWR VPWR _3593_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5330_ hold375/X _5579_/A0 _5330_/S VGND VGND VPWR VPWR _5330_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5261_ _5573_/A0 hold928/X _5267_/S VGND VGND VPWR VPWR _5261_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7000_ _7102_/CLK _7000_/D fanout503/X VGND VGND VPWR VPWR _7000_/Q sky130_fd_sc_hd__dfrtp_2
X_4212_ _4212_/A0 _6394_/A0 _4215_/S VGND VGND VPWR VPWR _4212_/X sky130_fd_sc_hd__mux2_1
X_5192_ _6397_/A0 hold478/X _5192_/S VGND VGND VPWR VPWR _5192_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4143_ _5459_/A0 hold289/X _4146_/S VGND VGND VPWR VPWR _4143_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4074_ _4074_/A0 _4073_/X _4086_/S VGND VGND VPWR VPWR _4074_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4976_ _5076_/B _5016_/A _5024_/A VGND VGND VPWR VPWR _4976_/X sky130_fd_sc_hd__a21o_1
X_6715_ _6963_/CLK _6715_/D fanout509/X VGND VGND VPWR VPWR _6715_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_189_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3927_ _6567_/Q _3927_/A1 _6461_/Q VGND VGND VPWR VPWR _3927_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3858_ _6541_/Q _3858_/B VGND VGND VPWR VPWR _3858_/X sky130_fd_sc_hd__and2b_1
X_6646_ _7196_/CLK _6646_/D VGND VGND VPWR VPWR _6646_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3789_ _3789_/A _3789_/B _3789_/C _3789_/D VGND VGND VPWR VPWR _3790_/D sky130_fd_sc_hd__or4_1
X_6577_ _6764_/CLK _6577_/D _6426_/A VGND VGND VPWR VPWR _6577_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_164_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5528_ _5579_/A0 hold415/X _5528_/S VGND VGND VPWR VPWR _5528_/X sky130_fd_sc_hd__mux2_1
X_5459_ _5459_/A0 hold341/X _5465_/S VGND VGND VPWR VPWR _5459_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7129_ _7129_/CLK _7129_/D fanout518/X VGND VGND VPWR VPWR _7129_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_47_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_170 _5574_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4830_ _5076_/A _4832_/B _4940_/A VGND VGND VPWR VPWR _5126_/B sky130_fd_sc_hd__a21oi_1
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_181 _3927_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_192 _3658_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4761_ _4761_/A _4761_/B _4761_/C _4760_/X VGND VGND VPWR VPWR _4761_/X sky130_fd_sc_hd__or4b_1
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3712_ input96/X _3547_/Y _5200_/A _6805_/Q VGND VGND VPWR VPWR _3712_/X sky130_fd_sc_hd__a22o_1
X_6500_ _7139_/CLK _6500_/D fanout518/X VGND VGND VPWR VPWR _6500_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_119_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4692_ _4814_/C _4692_/B VGND VGND VPWR VPWR _4863_/B sky130_fd_sc_hd__or2_1
XFILLER_174_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3643_ _7209_/Q _6392_/A _5187_/A _6795_/Q VGND VGND VPWR VPWR _3643_/X sky130_fd_sc_hd__a22o_1
X_6431_ _6432_/A _6441_/B VGND VGND VPWR VPWR _6431_/X sky130_fd_sc_hd__and2_1
XFILLER_147_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6362_ _6362_/A _6362_/B _6362_/C _6360_/X VGND VGND VPWR VPWR _6386_/S sky130_fd_sc_hd__or4b_4
X_3574_ _6684_/Q hold58/A _4246_/A _6704_/Q VGND VGND VPWR VPWR _3574_/X sky130_fd_sc_hd__a22o_1
X_5313_ hold22/X _5313_/B VGND VGND VPWR VPWR hold23/A sky130_fd_sc_hd__nand2_4
XFILLER_114_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6293_ _6598_/Q _6046_/B _6280_/X _6292_/X _6318_/S VGND VGND VPWR VPWR _6293_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_115_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5244_ _5496_/A0 hold868/X hold14/X VGND VGND VPWR VPWR _5244_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold18 hold18/A VGND VGND VPWR VPWR hold18/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 hold29/A VGND VGND VPWR VPWR hold29/X sky130_fd_sc_hd__buf_6
XFILLER_130_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5175_ _5137_/D _5174_/X _5148_/Y VGND VGND VPWR VPWR _5183_/B sky130_fd_sc_hd__o21a_1
XFILLER_69_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4126_ hold127/X hold193/X _4128_/S VGND VGND VPWR VPWR _4126_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4057_ hold425/X _4056_/X _4069_/S VGND VGND VPWR VPWR _4057_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4959_ _5123_/A _5163_/A _5163_/B VGND VGND VPWR VPWR _4959_/X sky130_fd_sc_hd__and3_1
XFILLER_177_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6629_ _7196_/CLK _6629_/D VGND VGND VPWR VPWR _6629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3290_ _3731_/A _3726_/B VGND VGND VPWR VPWR _3966_/A sky130_fd_sc_hd__nor2_8
XFILLER_111_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6980_ _7012_/CLK _6980_/D fanout505/X VGND VGND VPWR VPWR _6980_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_80_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5931_ _6614_/Q _5683_/X _5700_/X _6509_/Q VGND VGND VPWR VPWR _5931_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5862_ _7207_/Q _5671_/X _5682_/X _6511_/Q _5861_/X VGND VGND VPWR VPWR _5869_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_61_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4813_ _4985_/C _4813_/B _4813_/C _4813_/D VGND VGND VPWR VPWR _4815_/C sky130_fd_sc_hd__or4_1
X_5793_ _6846_/Q _5691_/Y _5785_/X _5792_/X _3195_/Y VGND VGND VPWR VPWR _5793_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_21_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4744_ _4758_/A _4758_/B _4744_/C VGND VGND VPWR VPWR _4744_/X sky130_fd_sc_hd__and3_1
XFILLER_159_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4675_ _4675_/A _4692_/B VGND VGND VPWR VPWR _4675_/Y sky130_fd_sc_hd__nor2_1
XFILLER_147_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6414_ _6426_/A _6441_/B VGND VGND VPWR VPWR _6414_/X sky130_fd_sc_hd__and2_1
X_3626_ input54/X _5232_/A _4300_/A _6748_/Q _3614_/X VGND VGND VPWR VPWR _3627_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_147_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3557_ _7029_/Q _3326_/Y _5403_/A _6981_/Q VGND VGND VPWR VPWR _3557_/X sky130_fd_sc_hd__a22o_1
X_6345_ _6346_/A _3888_/B _6692_/Q VGND VGND VPWR VPWR _6345_/X sky130_fd_sc_hd__o21a_1
X_6276_ _6508_/Q _6049_/B _6006_/Y _6753_/Q _6272_/X VGND VGND VPWR VPWR _6280_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3488_ _6878_/Q hold31/A _4104_/A _7214_/A VGND VGND VPWR VPWR _3488_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5227_ _5227_/A0 hold9/X _5228_/S VGND VGND VPWR VPWR hold10/A sky130_fd_sc_hd__mux2_1
Xinput108 wb_adr_i[18] VGND VGND VPWR VPWR _4337_/D sky130_fd_sc_hd__clkbuf_1
Xinput119 wb_adr_i[28] VGND VGND VPWR VPWR _3885_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_69_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5158_ _5158_/A _5158_/B _5158_/C VGND VGND VPWR VPWR _5159_/C sky130_fd_sc_hd__nor3_1
XFILLER_84_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4109_ _5567_/A0 hold799/X _4110_/S VGND VGND VPWR VPWR _4109_/X sky130_fd_sc_hd__mux2_1
X_5089_ _4996_/A _5094_/A _4659_/B _5021_/B VGND VGND VPWR VPWR _5089_/X sky130_fd_sc_hd__o22a_1
XFILLER_71_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_70 _5702_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_81 _6296_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_92 mask_rev_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4460_ _4759_/B _5001_/B VGND VGND VPWR VPWR _4860_/A sky130_fd_sc_hd__nand2_1
Xhold307 _7076_/Q VGND VGND VPWR VPWR hold307/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold318 _5415_/X VGND VGND VPWR VPWR _6988_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold329 _6590_/Q VGND VGND VPWR VPWR hold329/X sky130_fd_sc_hd__dlygate4sd3_1
X_3411_ _3410_/X _3449_/A1 _3791_/A VGND VGND VPWR VPWR _3411_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4391_ _4390_/C _4390_/D _4467_/A _4674_/A VGND VGND VPWR VPWR _4391_/Y sky130_fd_sc_hd__a31oi_2
XFILLER_98_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6130_ _7022_/Q _6204_/A2 _6007_/Y _7107_/Q _6129_/X VGND VGND VPWR VPWR _6130_/X
+ sky130_fd_sc_hd__a221o_1
X_3342_ _3546_/A hold76/X VGND VGND VPWR VPWR _5544_/A sky130_fd_sc_hd__nor2_8
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ _6915_/Q wire412/X _6024_/D _6939_/Q VGND VGND VPWR VPWR _6061_/X sky130_fd_sc_hd__a22o_1
X_3273_ hold66/X hold74/X VGND VGND VPWR VPWR hold67/A sky130_fd_sc_hd__and2b_4
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1007 hold1598/X VGND VGND VPWR VPWR _4093_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5012_ _4657_/A _4999_/A _4999_/B _5130_/B VGND VGND VPWR VPWR _5112_/C sky130_fd_sc_hd__a31o_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1018 _5352_/X VGND VGND VPWR VPWR _6932_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1029 _7111_/Q VGND VGND VPWR VPWR _5554_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6963_ _6963_/CLK _6963_/D fanout509/X VGND VGND VPWR VPWR _6963_/Q sky130_fd_sc_hd__dfstp_1
X_5914_ _7209_/Q _5671_/X _5706_/X _7092_/Q VGND VGND VPWR VPWR _5914_/X sky130_fd_sc_hd__a22o_1
XFILLER_62_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6894_ _7123_/CLK _6894_/D _6407_/A VGND VGND VPWR VPWR _6894_/Q sky130_fd_sc_hd__dfrtp_4
X_5845_ _6873_/Q _5683_/X _5703_/X _6857_/Q VGND VGND VPWR VPWR _5845_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5776_ _6918_/Q _5677_/X _5694_/X _7078_/Q VGND VGND VPWR VPWR _5776_/X sky130_fd_sc_hd__a22o_1
XFILLER_158_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4727_ _4739_/A _4724_/A _4726_/Y _6698_/Q VGND VGND VPWR VPWR _4992_/C sky130_fd_sc_hd__o31a_1
XFILLER_175_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4658_ _5021_/A _4784_/B VGND VGND VPWR VPWR _4713_/A sky130_fd_sc_hd__or2_1
XFILLER_135_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput90 spimemio_flash_io2_oeb VGND VGND VPWR VPWR input90/X sky130_fd_sc_hd__clkbuf_2
Xhold830 _6523_/Q VGND VGND VPWR VPWR hold830/X sky130_fd_sc_hd__dlygate4sd3_1
X_3609_ _6916_/Q _3334_/Y hold50/A _6677_/Q VGND VGND VPWR VPWR _3609_/X sky130_fd_sc_hd__a22o_1
Xhold841 _4099_/X VGND VGND VPWR VPWR _6571_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold852 _7088_/Q VGND VGND VPWR VPWR hold852/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4589_ _4814_/A _4675_/A VGND VGND VPWR VPWR _4694_/B sky130_fd_sc_hd__or2_4
XFILLER_150_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold863 _5522_/X VGND VGND VPWR VPWR _7083_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold874 _6703_/Q VGND VGND VPWR VPWR hold874/X sky130_fd_sc_hd__dlygate4sd3_1
X_6328_ _6605_/Q _5980_/Y _6038_/Y _6725_/Q _6327_/X VGND VGND VPWR VPWR _6331_/C
+ sky130_fd_sc_hd__a221o_1
Xhold885 _5383_/X VGND VGND VPWR VPWR _6960_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 _7128_/Q VGND VGND VPWR VPWR hold896/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6259_ _6747_/Q _6322_/B1 _6030_/X _6742_/Q _6258_/X VGND VGND VPWR VPWR _6267_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_29_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1530 _7170_/Q VGND VGND VPWR VPWR _5882_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1541 _7161_/Q VGND VGND VPWR VPWR _5649_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1552 hold16/A VGND VGND VPWR VPWR _3825_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1563 _6453_/Q VGND VGND VPWR VPWR _3859_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1574 _7154_/Q VGND VGND VPWR VPWR _5630_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1585 _7097_/Q VGND VGND VPWR VPWR hold265/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1596 _7117_/Q VGND VGND VPWR VPWR hold866/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3960_ _6824_/Q _3960_/B VGND VGND VPWR VPWR _3960_/X sky130_fd_sc_hd__and2_2
XFILLER_51_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3891_ _6541_/Q _3890_/A _3890_/Y _6543_/Q VGND VGND VPWR VPWR _6541_/D sky130_fd_sc_hd__a22o_1
XFILLER_189_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5630_ _5650_/B _6014_/A _6040_/A _5610_/X _5630_/B2 VGND VGND VPWR VPWR _7154_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5561_ _5579_/A0 hold433/X _5561_/S VGND VGND VPWR VPWR _5561_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4512_ _4742_/A _4512_/B VGND VGND VPWR VPWR _4515_/B sky130_fd_sc_hd__nand2_1
X_5492_ _5552_/A0 hold739/X _5492_/S VGND VGND VPWR VPWR _5492_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold104 _3253_/X VGND VGND VPWR VPWR hold104/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_156_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold115 _5562_/Y VGND VGND VPWR VPWR _5570_/S sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold126 hold132/X VGND VGND VPWR VPWR hold133/A sky130_fd_sc_hd__dlygate4sd3_1
X_4443_ _4445_/A _4453_/C VGND VGND VPWR VPWR _5003_/A sky130_fd_sc_hd__or2_4
XFILLER_171_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold137 _3964_/X VGND VGND VPWR VPWR hold137/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 _6714_/Q VGND VGND VPWR VPWR hold148/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold159 _3973_/X VGND VGND VPWR VPWR hold35/A sky130_fd_sc_hd__dlygate4sd3_1
X_7162_ _7183_/CLK _7162_/D fanout508/X VGND VGND VPWR VPWR _7162_/Q sky130_fd_sc_hd__dfrtp_1
X_4374_ _4745_/A _4532_/B VGND VGND VPWR VPWR _5112_/A sky130_fd_sc_hd__nor2_1
XFILLER_171_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3325_ hold29/X _3334_/A VGND VGND VPWR VPWR _5358_/A sky130_fd_sc_hd__nor2_8
X_6113_ _6941_/Q _6024_/D _6329_/B1 _7037_/Q VGND VGND VPWR VPWR _6113_/X sky130_fd_sc_hd__a22o_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7093_ _7093_/CLK _7093_/D fanout496/X VGND VGND VPWR VPWR _7093_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3256_ _3731_/A VGND VGND VPWR VPWR _3256_/Y sky130_fd_sc_hd__inv_2
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6044_ _6044_/A _6044_/B _6044_/C _6044_/D VGND VGND VPWR VPWR _6045_/C sky130_fd_sc_hd__or4_4
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3187_ _4654_/A VGND VGND VPWR VPWR _4546_/A sky130_fd_sc_hd__clkinv_2
XFILLER_94_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6946_ _7139_/CLK _6946_/D fanout518/X VGND VGND VPWR VPWR _6946_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_41_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6877_ _7138_/CLK _6877_/D fanout520/X VGND VGND VPWR VPWR _6877_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5828_ _6976_/Q _5960_/B VGND VGND VPWR VPWR _5828_/X sky130_fd_sc_hd__or2_1
XFILLER_167_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5759_ _7005_/Q _5664_/X _5688_/X _6861_/Q VGND VGND VPWR VPWR _5759_/X sky130_fd_sc_hd__a22o_1
XFILLER_135_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold660 _5398_/X VGND VGND VPWR VPWR _6973_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold671 _6535_/Q VGND VGND VPWR VPWR hold671/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold682 _5440_/X VGND VGND VPWR VPWR _7010_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold693 _6637_/Q VGND VGND VPWR VPWR hold693/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_618 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1360 hold1360/A VGND VGND VPWR VPWR wb_dat_o[20] sky130_fd_sc_hd__buf_12
XFILLER_45_523 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1371 _6587_/Q VGND VGND VPWR VPWR _4119_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1382 _6684_/Q VGND VGND VPWR VPWR _4238_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1393 _6672_/Q VGND VGND VPWR VPWR _4219_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput209 _3228_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[6] sky130_fd_sc_hd__buf_12
XFILLER_5_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4090_ _5243_/A1 hold9/X _4102_/S VGND VGND VPWR VPWR _4090_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6800_ _7207_/CLK _6800_/D fanout484/X VGND VGND VPWR VPWR _6800_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_91_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4992_ _4875_/X _4992_/B _4992_/C VGND VGND VPWR VPWR _5050_/C sky130_fd_sc_hd__and3b_1
X_6731_ _7211_/CLK _6731_/D fanout489/X VGND VGND VPWR VPWR _6731_/Q sky130_fd_sc_hd__dfrtp_2
X_3943_ input84/X _3872_/C _6460_/Q VGND VGND VPWR VPWR _3943_/X sky130_fd_sc_hd__mux2_2
XFILLER_16_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6662_ _6664_/CLK _6662_/D _3946_/B VGND VGND VPWR VPWR _6662_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_31_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3874_ _6457_/Q _3874_/A2 _6543_/Q _3834_/B VGND VGND VPWR VPWR _6442_/D sky130_fd_sc_hd__o211a_1
XFILLER_149_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5613_ _6564_/Q _5705_/B VGND VGND VPWR VPWR _5618_/B sky130_fd_sc_hd__nand2_1
X_6593_ _6969_/CLK _6593_/D fanout506/X VGND VGND VPWR VPWR _6593_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_191_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5544_ _5544_/A _5571_/B VGND VGND VPWR VPWR _5552_/S sky130_fd_sc_hd__nand2_8
XFILLER_145_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5475_ hold78/X _5571_/B VGND VGND VPWR VPWR hold79/A sky130_fd_sc_hd__nand2_8
XFILLER_117_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7214_ _7214_/A VGND VGND VPWR VPWR _7214_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_160_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4426_ _4462_/B _4426_/B VGND VGND VPWR VPWR _4947_/A sky130_fd_sc_hd__nand2_1
X_7145_ _7182_/CLK _7145_/D fanout502/X VGND VGND VPWR VPWR _7145_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_99_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout425 _4330_/B VGND VGND VPWR VPWR _6392_/B sky130_fd_sc_hd__buf_12
XFILLER_59_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4357_ _4621_/B _4781_/A VGND VGND VPWR VPWR _4360_/A sky130_fd_sc_hd__nor2_1
Xfanout436 hold39/X VGND VGND VPWR VPWR hold40/A sky130_fd_sc_hd__buf_6
XFILLER_86_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout447 hold85/X VGND VGND VPWR VPWR _5567_/A0 sky130_fd_sc_hd__buf_4
X_3308_ hold96/X _4111_/B VGND VGND VPWR VPWR _3308_/Y sky130_fd_sc_hd__nor2_8
Xfanout458 _5496_/A0 VGND VGND VPWR VPWR _5574_/A0 sky130_fd_sc_hd__clkbuf_8
X_7076_ _7137_/CLK _7076_/D fanout501/X VGND VGND VPWR VPWR _7076_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout469 hold565/X VGND VGND VPWR VPWR _5536_/A1 sky130_fd_sc_hd__buf_8
XFILLER_86_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4288_ _4288_/A _5580_/B VGND VGND VPWR VPWR _4293_/S sky130_fd_sc_hd__nand2_2
XFILLER_100_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6027_ _6027_/A _6027_/B _6027_/C _6027_/D VGND VGND VPWR VPWR _6029_/D sky130_fd_sc_hd__or4_1
X_3239_ _4605_/A VGND VGND VPWR VPWR _4793_/A sky130_fd_sc_hd__inv_2
XFILLER_86_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6929_ _6992_/CLK _6929_/D fanout517/X VGND VGND VPWR VPWR _6929_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_31_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7108_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_168_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_46_csclk _6931_/CLK VGND VGND VPWR VPWR _7037_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold490 _6501_/Q VGND VGND VPWR VPWR hold490/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_1_0_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_150_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1190 _4055_/X VGND VGND VPWR VPWR _6546_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3590_ _7077_/Q _5511_/A _4129_/A _6599_/Q _3561_/X VGND VGND VPWR VPWR _3593_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_139_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5260_ _5521_/A0 _5260_/A1 _5267_/S VGND VGND VPWR VPWR _5260_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4211_ _4211_/A0 _6393_/A0 _4215_/S VGND VGND VPWR VPWR _4211_/X sky130_fd_sc_hd__mux2_1
X_5191_ _6396_/A0 hold534/X _5192_/S VGND VGND VPWR VPWR _5191_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4142_ _5521_/A0 _4142_/A1 _4146_/S VGND VGND VPWR VPWR _4142_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4073_ hold922/X _5531_/A1 _4083_/S VGND VGND VPWR VPWR _4073_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4975_ _4971_/A _4797_/A _4607_/D _4974_/Y _4574_/Y VGND VGND VPWR VPWR _5095_/C
+ sky130_fd_sc_hd__a311o_1
X_6714_ _6725_/CLK _6714_/D fanout509/X VGND VGND VPWR VPWR _6714_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_51_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3926_ _6568_/Q input58/X _6462_/Q VGND VGND VPWR VPWR _3926_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6645_ _7196_/CLK _6645_/D VGND VGND VPWR VPWR _6645_/Q sky130_fd_sc_hd__dfxtp_1
X_3857_ _3858_/B _3857_/B VGND VGND VPWR VPWR _6454_/D sky130_fd_sc_hd__xnor2_1
XFILLER_165_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6576_ _7130_/CLK _6576_/D fanout519/X VGND VGND VPWR VPWR _6576_/Q sky130_fd_sc_hd__dfrtp_2
X_3788_ _3788_/A _3788_/B _3788_/C _3788_/D VGND VGND VPWR VPWR _3789_/D sky130_fd_sc_hd__or4_1
XFILLER_152_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5527_ _5578_/A0 hold852/X _5528_/S VGND VGND VPWR VPWR _5527_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_634 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5458_ _5536_/A1 _5458_/A1 _5465_/S VGND VGND VPWR VPWR _5458_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4409_ _4341_/X _4538_/B _4408_/Y VGND VGND VPWR VPWR _4433_/C sky130_fd_sc_hd__a21o_1
X_5389_ _5557_/A0 hold607/X _5393_/S VGND VGND VPWR VPWR _5389_/X sky130_fd_sc_hd__mux2_1
X_7128_ _7128_/CLK _7128_/D fanout514/X VGND VGND VPWR VPWR _7128_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_101_531 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7059_ _7078_/CLK _7059_/D fanout515/X VGND VGND VPWR VPWR _7059_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_131_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_160 _6206_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_171 _5531_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_182 _3927_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_193 _4022_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4760_ _4981_/B _4995_/A _4802_/A _4424_/Y _4758_/Y VGND VGND VPWR VPWR _4760_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3711_ _3714_/B hold76/X VGND VGND VPWR VPWR _5200_/A sky130_fd_sc_hd__nor2_2
XFILLER_147_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4691_ _4707_/A _4704_/B VGND VGND VPWR VPWR _4708_/B sky130_fd_sc_hd__or2_1
XFILLER_119_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6430_ _6433_/A _6441_/B VGND VGND VPWR VPWR _6430_/X sky130_fd_sc_hd__and2_1
XFILLER_146_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3642_ _3642_/A _3642_/B _3642_/C _3642_/D VGND VGND VPWR VPWR _3660_/B sky130_fd_sc_hd__or4_1
XFILLER_174_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6361_ _6358_/A _6389_/A2 _6699_/Q VGND VGND VPWR VPWR _6362_/B sky130_fd_sc_hd__a21boi_1
X_3573_ _3573_/A _3573_/B _3573_/C _3573_/D VGND VGND VPWR VPWR _3583_/C sky130_fd_sc_hd__or4_1
XFILLER_161_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5312_ _5579_/A0 hold554/X _5312_/S VGND VGND VPWR VPWR _5312_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6292_ _6292_/A _6292_/B _6292_/C VGND VGND VPWR VPWR _6292_/X sky130_fd_sc_hd__or3_1
XFILLER_114_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5243_ hold9/X _5243_/A1 hold14/X VGND VGND VPWR VPWR _5243_/X sky130_fd_sc_hd__mux2_1
Xhold19 hold19/A VGND VGND VPWR VPWR hold19/X sky130_fd_sc_hd__dlygate4sd3_1
X_5174_ _5174_/A _5174_/B _5174_/C _5173_/X VGND VGND VPWR VPWR _5174_/X sky130_fd_sc_hd__or4b_1
XFILLER_68_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4125_ _5558_/A0 hold209/X _4128_/S VGND VGND VPWR VPWR _4125_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_448 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4056_ hold237/X _5459_/A0 _4068_/S VGND VGND VPWR VPWR _4056_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4958_ _5002_/A _5035_/B _4832_/B _5108_/A _4957_/Y VGND VGND VPWR VPWR _5163_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_184_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3909_ _5650_/A _3908_/B _3906_/X _6819_/Q _6562_/Q VGND VGND VPWR VPWR _6564_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_177_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4889_ _4996_/A _5003_/A _4872_/B VGND VGND VPWR VPWR _4890_/D sky130_fd_sc_hd__a21oi_1
XFILLER_137_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6628_ _7193_/CLK _6628_/D VGND VGND VPWR VPWR _6628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6559_ _6969_/CLK _6559_/D fanout506/X VGND VGND VPWR VPWR _6559_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire431 _3887_/Y VGND VGND VPWR VPWR _3888_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_156_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5930_ _6754_/Q _5664_/X _5702_/X _6724_/Q _5929_/X VGND VGND VPWR VPWR _5935_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_80_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5861_ _6701_/Q _5659_/X _5693_/X _6655_/Q VGND VGND VPWR VPWR _5861_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4812_ _4984_/C _5090_/A _4805_/X _4811_/X VGND VGND VPWR VPWR _4813_/D sky130_fd_sc_hd__or4bb_1
XFILLER_61_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5792_ _5792_/A _5792_/B _5792_/C VGND VGND VPWR VPWR _5792_/X sky130_fd_sc_hd__or3_1
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4743_ _4981_/B _5003_/A VGND VGND VPWR VPWR _4764_/A sky130_fd_sc_hd__nor2_1
XFILLER_119_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4674_ _4674_/A _4684_/A VGND VGND VPWR VPWR _4692_/B sky130_fd_sc_hd__nand2_8
X_6413_ _6433_/A _6440_/B VGND VGND VPWR VPWR _6413_/X sky130_fd_sc_hd__and2_1
X_3625_ _6972_/Q _5394_/A _4252_/A _6708_/Q _3613_/X VGND VGND VPWR VPWR _3627_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_135_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6344_ _6344_/A1 _6319_/S _6342_/X _6343_/X VGND VGND VPWR VPWR _7187_/D sky130_fd_sc_hd__o22a_1
X_3556_ _6604_/Q _4135_/A _4312_/A _6759_/Q VGND VGND VPWR VPWR _3556_/X sky130_fd_sc_hd__a22o_1
XFILLER_103_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6275_ _6523_/Q _5994_/X _5998_/Y _6763_/Q _6274_/X VGND VGND VPWR VPWR _6280_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_163_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3487_ _7054_/Q _3684_/B1 _4083_/S _3487_/B2 _3486_/X VGND VGND VPWR VPWR _3499_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_115_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5226_ _5226_/A0 _5574_/A0 _5228_/S VGND VGND VPWR VPWR _5226_/X sky130_fd_sc_hd__mux2_1
Xinput109 wb_adr_i[19] VGND VGND VPWR VPWR _4337_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_130_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5157_ _5110_/C _5153_/X _5178_/C _5156_/Y VGND VGND VPWR VPWR _5157_/X sky130_fd_sc_hd__o31a_1
XFILLER_56_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4108_ _6396_/A0 hold699/X _4110_/S VGND VGND VPWR VPWR _4108_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5088_ _6779_/Q _6362_/A _5070_/Y _5087_/X VGND VGND VPWR VPWR _5104_/C sky130_fd_sc_hd__a22o_1
X_4039_ hold467/X _6397_/A0 _4039_/S VGND VGND VPWR VPWR _4039_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_60 _5663_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_71 _5703_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_82 _6332_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_93 mask_rev_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold308 _5514_/X VGND VGND VPWR VPWR _7076_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold319 _6952_/Q VGND VGND VPWR VPWR hold319/X sky130_fd_sc_hd__dlygate4sd3_1
X_3410_ _3410_/A _3410_/B VGND VGND VPWR VPWR _3410_/X sky130_fd_sc_hd__or2_4
XFILLER_109_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4390_ _4390_/A _4654_/A _4390_/C _4390_/D VGND VGND VPWR VPWR _4693_/A sky130_fd_sc_hd__or4_4
XFILLER_98_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3341_ _3534_/A hold76/X VGND VGND VPWR VPWR _3341_/Y sky130_fd_sc_hd__nor2_2
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6060_ _7112_/Q _6322_/B1 _6030_/X _6995_/Q _6059_/X VGND VGND VPWR VPWR _6069_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_140_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3272_ hold27/X hold55/X VGND VGND VPWR VPWR hold28/A sky130_fd_sc_hd__and2b_4
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1008 _4093_/X VGND VGND VPWR VPWR _6568_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5011_ _4873_/Y _5130_/B _5010_/X _5050_/C VGND VGND VPWR VPWR _5033_/B sky130_fd_sc_hd__o31a_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1019 _6903_/Q VGND VGND VPWR VPWR _5319_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6962_ _6990_/CLK _6962_/D _3873_/A VGND VGND VPWR VPWR _6962_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_53_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5913_ _5913_/A _5913_/B _5913_/C _5913_/D VGND VGND VPWR VPWR _5913_/X sky130_fd_sc_hd__or4_1
X_6893_ _6925_/CLK _6893_/D fanout516/X VGND VGND VPWR VPWR _6893_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_21_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5844_ _6881_/Q _5667_/X _5843_/X VGND VGND VPWR VPWR _5847_/C sky130_fd_sc_hd__a21o_1
XFILLER_34_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5775_ _6886_/Q _5846_/A2 _5848_/B1 _7046_/Q VGND VGND VPWR VPWR _5775_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4726_ _5001_/C VGND VGND VPWR VPWR _4726_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4657_ _4657_/A _4999_/A _4657_/C VGND VGND VPWR VPWR _5130_/A sky130_fd_sc_hd__and3_1
XFILLER_175_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput80 spi_sck VGND VGND VPWR VPWR input80/X sky130_fd_sc_hd__clkbuf_1
Xhold820 _5397_/X VGND VGND VPWR VPWR _6972_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3608_ _7113_/Q _5553_/A _5562_/A _7121_/Q VGND VGND VPWR VPWR _3608_/X sky130_fd_sc_hd__a22o_1
XFILLER_174_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput91 spimemio_flash_io3_do VGND VGND VPWR VPWR input91/X sky130_fd_sc_hd__clkbuf_1
Xhold831 _4031_/X VGND VGND VPWR VPWR _6523_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4588_ _4588_/A _4605_/A _4621_/B _4935_/A VGND VGND VPWR VPWR _4675_/A sky130_fd_sc_hd__or4bb_4
Xhold842 _6864_/Q VGND VGND VPWR VPWR hold842/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold853 _5527_/X VGND VGND VPWR VPWR _7088_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6327_ _6679_/Q _5992_/X _6020_/X _6710_/Q VGND VGND VPWR VPWR _6327_/X sky130_fd_sc_hd__a22o_1
Xhold864 _6987_/Q VGND VGND VPWR VPWR hold864/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold875 _4249_/X VGND VGND VPWR VPWR _6703_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3539_ _6854_/Q _5259_/A hold50/A _6679_/Q VGND VGND VPWR VPWR _3539_/X sky130_fd_sc_hd__a22o_2
XFILLER_107_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold886 _7048_/Q VGND VGND VPWR VPWR hold886/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold897 _5573_/X VGND VGND VPWR VPWR _7128_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6258_ _6717_/Q _6023_/B _6338_/B1 _6767_/Q _6246_/X VGND VGND VPWR VPWR _6258_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5209_ hold285/X _5539_/A1 _5209_/S VGND VGND VPWR VPWR _5209_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6189_ _7088_/Q _5977_/X _6025_/C _7117_/Q _6188_/X VGND VGND VPWR VPWR _6192_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1520 hold42/A VGND VGND VPWR VPWR _3865_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1531 _6780_/Q VGND VGND VPWR VPWR hold1531/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1542 _6653_/Q VGND VGND VPWR VPWR _4196_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1553 _6691_/Q VGND VGND VPWR VPWR _3188_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1564 _6545_/Q VGND VGND VPWR VPWR _3913_/B1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1575 _7184_/Q VGND VGND VPWR VPWR _6270_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1586 _6456_/Q VGND VGND VPWR VPWR _3847_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1597 _6564_/Q VGND VGND VPWR VPWR _3901_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_189_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3890_ _3890_/A _3890_/B VGND VGND VPWR VPWR _3890_/Y sky130_fd_sc_hd__nor2_1
XFILLER_188_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5560_ _5578_/A0 hold866/X _5561_/S VGND VGND VPWR VPWR _5560_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4511_ _4871_/A _5003_/A _4508_/X _4510_/X VGND VGND VPWR VPWR _4515_/A sky130_fd_sc_hd__o211a_1
XFILLER_144_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5491_ _5587_/A0 hold890/X _5492_/S VGND VGND VPWR VPWR _5491_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold105 _3254_/X VGND VGND VPWR VPWR _3301_/C sky130_fd_sc_hd__dlygate4sd3_1
X_4442_ _4445_/A _4453_/C VGND VGND VPWR VPWR _4512_/B sky130_fd_sc_hd__nor2_2
Xhold116 _5569_/X VGND VGND VPWR VPWR _7125_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 hold127/A VGND VGND VPWR VPWR hold127/X sky130_fd_sc_hd__clkbuf_16
Xhold138 _4141_/Y VGND VGND VPWR VPWR _4146_/S sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 _4262_/X VGND VGND VPWR VPWR _6714_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7161_ _7181_/CLK _7161_/D fanout499/X VGND VGND VPWR VPWR _7161_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_144_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4373_ _4846_/B _4781_/B VGND VGND VPWR VPWR _4532_/B sky130_fd_sc_hd__or2_2
XFILLER_98_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6112_ _7085_/Q _5977_/X _6025_/A _6861_/Q _6111_/X VGND VGND VPWR VPWR _6119_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3324_ _3526_/A _3334_/A VGND VGND VPWR VPWR _5340_/A sky130_fd_sc_hd__nor2_8
X_7092_ _7209_/CLK _7092_/D fanout485/X VGND VGND VPWR VPWR _7092_/Q sky130_fd_sc_hd__dfstp_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6043_ _6954_/Q _6336_/A2 _6037_/X _6042_/X VGND VGND VPWR VPWR _6044_/D sky130_fd_sc_hd__a211o_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3255_ _3301_/C hold48/X hold18/X VGND VGND VPWR VPWR _3255_/X sky130_fd_sc_hd__or3b_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3186_ _6445_/Q VGND VGND VPWR VPWR _3868_/A sky130_fd_sc_hd__inv_2
XFILLER_27_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6945_ _6992_/CLK _6945_/D fanout517/X VGND VGND VPWR VPWR _6945_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_53_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6876_ _7129_/CLK _6876_/D fanout518/X VGND VGND VPWR VPWR _6876_/Q sky130_fd_sc_hd__dfrtp_2
X_5827_ _7000_/Q _5656_/X _5696_/X _7040_/Q _5826_/X VGND VGND VPWR VPWR _5835_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_22_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5758_ _6893_/Q _5655_/X _5756_/X _5757_/X VGND VGND VPWR VPWR _5771_/A sky130_fd_sc_hd__a211o_1
XFILLER_182_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4709_ _4471_/B _4677_/B _5054_/B _4708_/X VGND VGND VPWR VPWR _4709_/X sky130_fd_sc_hd__o211a_1
X_5689_ _5705_/B _5703_/B VGND VGND VPWR VPWR _5689_/X sky130_fd_sc_hd__and2_4
XFILLER_108_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold650 _5435_/X VGND VGND VPWR VPWR _7006_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold661 _6862_/Q VGND VGND VPWR VPWR hold661/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold672 _4045_/X VGND VGND VPWR VPWR _6535_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap391 _6038_/Y VGND VGND VPWR VPWR _6206_/B1 sky130_fd_sc_hd__buf_12
Xhold683 _6768_/Q VGND VGND VPWR VPWR hold683/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 _4178_/X VGND VGND VPWR VPWR _6637_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1350 hold1350/A VGND VGND VPWR VPWR wb_dat_o[28] sky130_fd_sc_hd__buf_12
XFILLER_85_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1361 _6354_/A0 VGND VGND VPWR VPWR hold1361/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1372 _6586_/Q VGND VGND VPWR VPWR _4118_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1383 _7125_/Q VGND VGND VPWR VPWR _5569_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1394 _6806_/Q VGND VGND VPWR VPWR _5204_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4991_ _5103_/A _4991_/B VGND VGND VPWR VPWR _4991_/Y sky130_fd_sc_hd__nor2_1
XFILLER_91_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6730_ _6740_/CLK _6730_/D _3873_/A VGND VGND VPWR VPWR _6730_/Q sky130_fd_sc_hd__dfstp_1
X_3942_ _3971_/S _3942_/A2 _6407_/B _3941_/Y VGND VGND VPWR VPWR _3942_/X sky130_fd_sc_hd__a22o_2
XFILLER_189_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6661_ _6664_/CLK _6661_/D fanout485/X VGND VGND VPWR VPWR _6661_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_32_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3873_ _3873_/A _6407_/B VGND VGND VPWR VPWR _3873_/X sky130_fd_sc_hd__and2_1
XFILLER_176_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5612_ _7149_/Q _7148_/Q VGND VGND VPWR VPWR _5705_/B sky130_fd_sc_hd__nor2_4
X_6592_ _7141_/CLK _6592_/D fanout504/X VGND VGND VPWR VPWR _6592_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_191_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5543_ hold729/X _5552_/A0 _5543_/S VGND VGND VPWR VPWR _5543_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5474_ hold733/X _5552_/A0 _5474_/S VGND VGND VPWR VPWR _5474_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7213_ _7213_/A VGND VGND VPWR VPWR _7213_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_105_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4425_ _4742_/A _4485_/A VGND VGND VPWR VPWR _4504_/A sky130_fd_sc_hd__nand2_1
XFILLER_144_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7144_ _7181_/CLK _7144_/D fanout502/X VGND VGND VPWR VPWR _7144_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_113_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4356_ _4354_/A _4354_/B _4355_/Y _4350_/B VGND VGND VPWR VPWR _4944_/A sky130_fd_sc_hd__o2bb2ai_2
XFILLER_98_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout426 _5535_/B VGND VGND VPWR VPWR _4330_/B sky130_fd_sc_hd__buf_8
XFILLER_86_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout437 _5569_/A0 VGND VGND VPWR VPWR _5587_/A0 sky130_fd_sc_hd__buf_6
XFILLER_113_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3307_ hold67/X _3378_/B VGND VGND VPWR VPWR _4111_/B sky130_fd_sc_hd__nand2_8
Xfanout448 hold84/X VGND VGND VPWR VPWR hold85/A sky130_fd_sc_hd__buf_6
X_7075_ _7075_/CLK _7075_/D fanout515/X VGND VGND VPWR VPWR _7075_/Q sky130_fd_sc_hd__dfstp_1
Xfanout459 hold44/X VGND VGND VPWR VPWR _5496_/A0 sky130_fd_sc_hd__buf_4
X_4287_ _6397_/A0 hold455/X _4287_/S VGND VGND VPWR VPWR _4287_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6026_ _6026_/A _6026_/B _6026_/C _6026_/D VGND VGND VPWR VPWR _6029_/C sky130_fd_sc_hd__or4_1
XFILLER_100_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3238_ _4570_/D VGND VGND VPWR VPWR _4846_/C sky130_fd_sc_hd__clkinv_8
XFILLER_67_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6928_ _6977_/CLK _6928_/D fanout507/X VGND VGND VPWR VPWR _6928_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6859_ _6883_/CLK _6859_/D fanout505/X VGND VGND VPWR VPWR _6859_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_168_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold480 _6745_/Q VGND VGND VPWR VPWR hold480/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold491 _4005_/X VGND VGND VPWR VPWR _6501_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1180 _7095_/Q VGND VGND VPWR VPWR _5536_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1191 _6994_/Q VGND VGND VPWR VPWR _5422_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4210_ _4210_/A _4330_/B VGND VGND VPWR VPWR _4215_/S sky130_fd_sc_hd__and2_2
X_5190_ _6395_/A0 _5190_/A1 _5192_/S VGND VGND VPWR VPWR _5190_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4141_ _4141_/A _5580_/B VGND VGND VPWR VPWR _4141_/Y sky130_fd_sc_hd__nand2_2
X_4072_ _4072_/A0 _4071_/X _4086_/S VGND VGND VPWR VPWR _4072_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4974_ _4981_/B _5021_/B _4794_/A _5021_/A VGND VGND VPWR VPWR _4974_/Y sky130_fd_sc_hd__a211oi_1
X_3925_ _6577_/Q input81/X _3958_/B VGND VGND VPWR VPWR _3925_/X sky130_fd_sc_hd__mux2_8
XFILLER_51_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6713_ _6963_/CLK _6713_/D fanout509/X VGND VGND VPWR VPWR _6713_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_149_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6644_ _7193_/CLK _6644_/D VGND VGND VPWR VPWR _6644_/Q sky130_fd_sc_hd__dfxtp_1
X_3856_ _6454_/Q _3856_/B VGND VGND VPWR VPWR _3857_/B sky130_fd_sc_hd__nor2_1
XFILLER_137_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6575_ _6764_/CLK _6575_/D _6426_/A VGND VGND VPWR VPWR _6575_/Q sky130_fd_sc_hd__dfrtp_1
X_3787_ _7010_/Q _5439_/A _3727_/Y _6812_/Q _3734_/X VGND VGND VPWR VPWR _3788_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_164_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5526_ _5550_/A0 hold419/X _5528_/S VGND VGND VPWR VPWR _5526_/X sky130_fd_sc_hd__mux2_1
X_5457_ _5457_/A _5535_/B VGND VGND VPWR VPWR _5465_/S sky130_fd_sc_hd__nand2_8
XFILLER_160_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4408_ _4621_/B _4538_/B _4605_/A VGND VGND VPWR VPWR _4408_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_182_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5388_ _5496_/A0 hold815/X _5393_/S VGND VGND VPWR VPWR _5388_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7127_ _7130_/CLK _7127_/D fanout521/X VGND VGND VPWR VPWR _7127_/Q sky130_fd_sc_hd__dfstp_1
X_4339_ _4339_/A _4339_/B _4339_/C _4339_/D VGND VGND VPWR VPWR _4348_/C sky130_fd_sc_hd__and4_1
XFILLER_101_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7058_ _7135_/CLK _7058_/D fanout521/X VGND VGND VPWR VPWR _7058_/Q sky130_fd_sc_hd__dfstp_4
X_6009_ _6040_/B _6039_/C _6030_/C VGND VGND VPWR VPWR _6009_/X sky130_fd_sc_hd__and3_4
XFILLER_39_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_150 _6496_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_161 _6027_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_172 _5555_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_183 _3927_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_194 _3499_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3710_ _3710_/A _3710_/B _3710_/C _3710_/D VGND VGND VPWR VPWR _3722_/C sky130_fd_sc_hd__or4_1
XFILLER_147_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4690_ _4707_/A _4692_/B VGND VGND VPWR VPWR _4708_/A sky130_fd_sc_hd__or2_1
XFILLER_186_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3641_ input26/X _3304_/Y _4040_/A _6533_/Q _3640_/X VGND VGND VPWR VPWR _3642_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6360_ _6358_/A _6360_/A2 _6696_/Q VGND VGND VPWR VPWR _6360_/X sky130_fd_sc_hd__a21bo_1
X_3572_ _6861_/Q _5268_/A _4147_/A _6614_/Q _3571_/X VGND VGND VPWR VPWR _3573_/D
+ sky130_fd_sc_hd__a221o_1
X_5311_ _5578_/A0 hold846/X _5312_/S VGND VGND VPWR VPWR _5311_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6291_ _6291_/A _6291_/B _6291_/C _6291_/D VGND VGND VPWR VPWR _6292_/C sky130_fd_sc_hd__or4_2
XFILLER_142_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5242_ _5581_/A0 hold918/X hold14/X VGND VGND VPWR VPWR _5242_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_30_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7053_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_68_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5173_ _4981_/B _5003_/A _5036_/B _4996_/A _4510_/C VGND VGND VPWR VPWR _5173_/X
+ sky130_fd_sc_hd__o221a_1
X_4124_ _5539_/A1 hold295/X _4128_/S VGND VGND VPWR VPWR _4124_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput1 debug_mode VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__clkbuf_2
X_4055_ _4055_/A0 _4054_/X _4069_/S VGND VGND VPWR VPWR _4055_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_45_csclk _6931_/CLK VGND VGND VPWR VPWR _7071_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4957_ _4957_/A _4957_/B VGND VGND VPWR VPWR _4957_/Y sky130_fd_sc_hd__nand2_1
XFILLER_52_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3908_ _5650_/A _3908_/B VGND VGND VPWR VPWR _3908_/Y sky130_fd_sc_hd__nand2_1
X_4888_ _4759_/B _4871_/Y _4984_/B _5065_/A VGND VGND VPWR VPWR _4890_/C sky130_fd_sc_hd__a211o_1
XFILLER_138_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3839_ _6471_/Q _3839_/B VGND VGND VPWR VPWR _3840_/S sky130_fd_sc_hd__nor2_1
X_6627_ _7196_/CLK _6627_/D VGND VGND VPWR VPWR _6627_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6558_ _7141_/CLK _6558_/D fanout504/X VGND VGND VPWR VPWR _6558_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5509_ _5587_/A0 hold834/X _5510_/S VGND VGND VPWR VPWR _5509_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6489_ _6825_/CLK _6489_/D fanout498/X VGND VGND VPWR VPWR _6489_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_106_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire476 hold11/X VGND VGND VPWR VPWR hold12/A sky130_fd_sc_hd__buf_4
XFILLER_171_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5860_ _5860_/A0 _5859_/X _6319_/S VGND VGND VPWR VPWR _7169_/D sky130_fd_sc_hd__mux2_1
XFILLER_61_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4811_ _4814_/B _4694_/B _4759_/Y _4786_/Y _4810_/X VGND VGND VPWR VPWR _4811_/X
+ sky130_fd_sc_hd__o2111a_1
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5791_ _6934_/Q _5670_/X _5686_/X _7014_/Q _5790_/X VGND VGND VPWR VPWR _5792_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_61_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4742_ _4742_/A _4758_/A _4742_/C VGND VGND VPWR VPWR _5134_/A sky130_fd_sc_hd__and3_1
X_4673_ _4694_/B _5016_/B VGND VGND VPWR VPWR _5107_/C sky130_fd_sc_hd__nor2_1
X_6412_ _6433_/A _6441_/B VGND VGND VPWR VPWR _6412_/X sky130_fd_sc_hd__and2_1
X_3624_ _6908_/Q _5322_/A _4147_/A _6613_/Q _3611_/X VGND VGND VPWR VPWR _3627_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_174_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6343_ _7186_/Q _5592_/Y _5650_/Y VGND VGND VPWR VPWR _6343_/X sky130_fd_sc_hd__o21ba_1
XFILLER_127_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3555_ _6845_/Q _5250_/A _4046_/A _6539_/Q VGND VGND VPWR VPWR _3555_/X sky130_fd_sc_hd__a22o_1
XFILLER_127_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6274_ _6513_/Q _5977_/X _6323_/B1 _6738_/Q VGND VGND VPWR VPWR _6274_/X sky130_fd_sc_hd__a22o_1
X_3486_ _6982_/Q _5403_/A _6392_/A _7211_/Q VGND VGND VPWR VPWR _3486_/X sky130_fd_sc_hd__a22o_1
X_5225_ _5225_/A _5535_/B VGND VGND VPWR VPWR _5228_/S sky130_fd_sc_hd__and2_4
XFILLER_69_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5156_ _5156_/A _5156_/B _5156_/C VGND VGND VPWR VPWR _5156_/Y sky130_fd_sc_hd__nor3_1
XFILLER_29_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4107_ hold44/X hold281/X _4110_/S VGND VGND VPWR VPWR _4107_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5087_ _5155_/B _5087_/B VGND VGND VPWR VPWR _5087_/X sky130_fd_sc_hd__or2_1
XFILLER_84_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4038_ hold496/X _6396_/A0 _4039_/S VGND VGND VPWR VPWR _4038_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5989_ _6000_/A _6033_/A _6020_/C VGND VGND VPWR VPWR _6022_/B sky130_fd_sc_hd__and3_4
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_50 _4128_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_61 _5664_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_72 _5705_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_83 _6930_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_94 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput190 _3211_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[23] sky130_fd_sc_hd__buf_12
XFILLER_94_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold309 _7044_/Q VGND VGND VPWR VPWR hold309/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3340_ _5212_/A _3340_/B VGND VGND VPWR VPWR _3340_/Y sky130_fd_sc_hd__nor2_8
Xclkbuf_3_4_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A VGND VGND VPWR VPWR _7193_/CLK sky130_fd_sc_hd__clkbuf_8
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3271_ hold94/X hold19/X VGND VGND VPWR VPWR hold95/A sky130_fd_sc_hd__or2_4
XFILLER_97_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _5042_/C _5148_/B _5134_/B _5010_/D VGND VGND VPWR VPWR _5010_/X sky130_fd_sc_hd__or4_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1009 _6919_/Q VGND VGND VPWR VPWR _5337_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6961_ _7141_/CLK _6961_/D fanout506/X VGND VGND VPWR VPWR _6961_/Q sky130_fd_sc_hd__dfrtp_4
X_5912_ _6528_/Q _5676_/X _5703_/X _6603_/Q _5911_/X VGND VGND VPWR VPWR _5913_/D
+ sky130_fd_sc_hd__a221o_1
X_6892_ _6925_/CLK _6892_/D fanout516/X VGND VGND VPWR VPWR _6892_/Q sky130_fd_sc_hd__dfrtp_4
X_5843_ _7025_/Q _5663_/X _5682_/X _7089_/Q VGND VGND VPWR VPWR _5843_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5774_ _5794_/A2 _5773_/X _6319_/S VGND VGND VPWR VPWR _5774_/X sky130_fd_sc_hd__mux2_1
XFILLER_166_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4725_ _4731_/C _4731_/B _4724_/B _4547_/A VGND VGND VPWR VPWR _5001_/C sky130_fd_sc_hd__a211oi_4
XFILLER_135_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4656_ _5021_/A _4942_/A VGND VGND VPWR VPWR _4656_/Y sky130_fd_sc_hd__nor2_1
XFILLER_190_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3607_ _3714_/B _4111_/B VGND VGND VPWR VPWR _5225_/A sky130_fd_sc_hd__nor2_2
Xinput70 mgmt_gpio_in[7] VGND VGND VPWR VPWR _3960_/B sky130_fd_sc_hd__buf_2
Xinput81 spi_sdo VGND VGND VPWR VPWR input81/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold810 _5338_/X VGND VGND VPWR VPWR _6920_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_174_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold821 _7016_/Q VGND VGND VPWR VPWR hold821/X sky130_fd_sc_hd__dlygate4sd3_1
X_4587_ _5016_/A _4677_/B VGND VGND VPWR VPWR _4965_/A sky130_fd_sc_hd__nor2_1
XFILLER_116_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold832 _6936_/Q VGND VGND VPWR VPWR hold832/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput92 spimemio_flash_io3_oeb VGND VGND VPWR VPWR input92/X sky130_fd_sc_hd__clkbuf_2
Xhold843 _5275_/X VGND VGND VPWR VPWR _6864_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6326_ _6610_/Q _6326_/A2 _6033_/X _7211_/Q _6325_/X VGND VGND VPWR VPWR _6331_/B
+ sky130_fd_sc_hd__a221o_1
X_3538_ hold49/X _3538_/B VGND VGND VPWR VPWR hold50/A sky130_fd_sc_hd__nor2_4
Xhold854 _6892_/Q VGND VGND VPWR VPWR hold854/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold865 _5414_/X VGND VGND VPWR VPWR _6987_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 hold876/A VGND VGND VPWR VPWR hold876/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold887 _5482_/X VGND VGND VPWR VPWR _7048_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_107_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold898 _6499_/Q VGND VGND VPWR VPWR hold898/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_107_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6257_ _6257_/A _6257_/B _6257_/C _6257_/D VGND VGND VPWR VPWR _6257_/X sky130_fd_sc_hd__or4_1
XFILLER_88_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3469_ _6846_/Q _5250_/A _5511_/A _7078_/Q VGND VGND VPWR VPWR _3469_/X sky130_fd_sc_hd__a22o_1
XFILLER_103_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5208_ hold331/X _5583_/A0 _5209_/S VGND VGND VPWR VPWR _5208_/X sky130_fd_sc_hd__mux2_1
XFILLER_190_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6188_ _6960_/Q _6336_/A2 _6205_/B1 _7064_/Q VGND VGND VPWR VPWR _6188_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1510 _6171_/X VGND VGND VPWR VPWR _7180_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1521 _6450_/Q VGND VGND VPWR VPWR _3862_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5139_ _5139_/A _5139_/B _5139_/C _5139_/D VGND VGND VPWR VPWR _6780_/D sky130_fd_sc_hd__or4_1
Xhold1532 _7200_/Q VGND VGND VPWR VPWR _6374_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1543 _6445_/Q VGND VGND VPWR VPWR _3914_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1554 _3911_/Y VGND VGND VPWR VPWR _6691_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1565 _3841_/X VGND VGND VPWR VPWR _6459_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1576 _6591_/Q VGND VGND VPWR VPWR hold295/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1587 _6595_/Q VGND VGND VPWR VPWR hold755/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1598 _6568_/Q VGND VGND VPWR VPWR hold1598/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4510_ _4510_/A _4510_/B _4510_/C VGND VGND VPWR VPWR _4510_/X sky130_fd_sc_hd__and3_1
XFILLER_117_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5490_ _5586_/A0 _5490_/A1 _5492_/S VGND VGND VPWR VPWR _5490_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold106 _3281_/X VGND VGND VPWR VPWR _3525_/A sky130_fd_sc_hd__dlygate4sd3_1
X_4441_ _4441_/A _4453_/C VGND VGND VPWR VPWR _4994_/A sky130_fd_sc_hd__or2_2
XFILLER_172_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold117 _6880_/Q VGND VGND VPWR VPWR hold117/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold128 _4117_/X VGND VGND VPWR VPWR _6585_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 _4145_/X VGND VGND VPWR VPWR _6609_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7160_ _7182_/CLK _7160_/D fanout499/X VGND VGND VPWR VPWR _7160_/Q sky130_fd_sc_hd__dfrtp_1
X_4372_ _4846_/B _4781_/B VGND VGND VPWR VPWR _4993_/A sky130_fd_sc_hd__nor2_8
XFILLER_171_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6111_ _7005_/Q _6202_/B1 _6024_/C _6909_/Q VGND VGND VPWR VPWR _6111_/X sky130_fd_sc_hd__a22o_1
XFILLER_125_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3323_ _3546_/B _3476_/A VGND VGND VPWR VPWR _5466_/A sky130_fd_sc_hd__nor2_8
XFILLER_98_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7091_ _7094_/CLK _7091_/D fanout494/X VGND VGND VPWR VPWR _7091_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6042_ _6978_/Q _6206_/B1 _6272_/B _7066_/Q _6041_/X VGND VGND VPWR VPWR _6042_/X
+ sky130_fd_sc_hd__a221o_1
X_3254_ hold104/X _5168_/A1 _3971_/S VGND VGND VPWR VPWR _3254_/X sky130_fd_sc_hd__mux2_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3185_ hold25/A VGND VGND VPWR VPWR _3830_/A sky130_fd_sc_hd__inv_2
XFILLER_54_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6944_ _6977_/CLK _6944_/D fanout517/X VGND VGND VPWR VPWR _6944_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_179_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6875_ _7135_/CLK hold33/X fanout519/X VGND VGND VPWR VPWR _6875_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_22_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5826_ _6936_/Q _5670_/X _5672_/X _6928_/Q VGND VGND VPWR VPWR _5826_/X sky130_fd_sc_hd__a22o_1
XFILLER_139_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5757_ _6917_/Q _5677_/X _5694_/X _7077_/Q _5754_/X VGND VGND VPWR VPWR _5757_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4708_ _4708_/A _4708_/B _4708_/C _4850_/B VGND VGND VPWR VPWR _4708_/X sky130_fd_sc_hd__and4_1
XFILLER_175_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5688_ _5938_/B _5703_/B _5699_/B VGND VGND VPWR VPWR _5688_/X sky130_fd_sc_hd__and3_4
XFILLER_108_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4639_ _4639_/A _4639_/B VGND VGND VPWR VPWR _4985_/A sky130_fd_sc_hd__nor2_1
XFILLER_150_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold640 _5480_/X VGND VGND VPWR VPWR _7046_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold651 _7067_/Q VGND VGND VPWR VPWR hold651/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap370 hold107/X VGND VGND VPWR VPWR _5493_/A sky130_fd_sc_hd__buf_8
Xhold662 _5273_/X VGND VGND VPWR VPWR _6862_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap381 _3530_/B VGND VGND VPWR VPWR _3334_/A sky130_fd_sc_hd__buf_12
Xhold673 _7031_/Q VGND VGND VPWR VPWR hold673/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap392 _6021_/Y VGND VGND VPWR VPWR _6027_/D sky130_fd_sc_hd__buf_12
Xhold684 _4327_/X VGND VGND VPWR VPWR _6768_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6309_ _6749_/Q _6322_/B1 _6030_/X _6744_/Q _6308_/X VGND VGND VPWR VPWR _6316_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold695 _7094_/Q VGND VGND VPWR VPWR hold695/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1340 hold1340/A VGND VGND VPWR VPWR wb_dat_o[31] sky130_fd_sc_hd__buf_12
Xhold1351 _4194_/A0 VGND VGND VPWR VPWR hold1351/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1362 hold1362/A VGND VGND VPWR VPWR wb_dat_o[29] sky130_fd_sc_hd__buf_12
Xhold1373 _6835_/Q VGND VGND VPWR VPWR _5243_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1384 _6678_/Q VGND VGND VPWR VPWR _4226_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1395 _6495_/Q VGND VGND VPWR VPWR _3998_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xnet499_2 net499_2/A VGND VGND VPWR VPWR _3941_/B sky130_fd_sc_hd__inv_2
X_4990_ _4979_/X _4990_/B VGND VGND VPWR VPWR _4991_/B sky130_fd_sc_hd__and2b_1
XFILLER_90_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3941_ _3971_/S _3941_/B VGND VGND VPWR VPWR _3941_/Y sky130_fd_sc_hd__nor2_2
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6660_ _6664_/CLK _6660_/D fanout485/X VGND VGND VPWR VPWR _6660_/Q sky130_fd_sc_hd__dfrtp_4
X_3872_ _6820_/Q _6869_/Q _3872_/C VGND VGND VPWR VPWR _3872_/Y sky130_fd_sc_hd__nor3_2
XFILLER_189_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5611_ _6564_/Q _5609_/Y _5611_/S VGND VGND VPWR VPWR _7148_/D sky130_fd_sc_hd__mux2_1
XFILLER_149_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6591_ _7033_/CLK _6591_/D fanout504/X VGND VGND VPWR VPWR _6591_/Q sky130_fd_sc_hd__dfrtp_1
X_5542_ hold902/X _5587_/A0 _5543_/S VGND VGND VPWR VPWR _5542_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5473_ hold910/X _5587_/A0 _5474_/S VGND VGND VPWR VPWR _5473_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4424_ _4758_/A _4758_/B _4758_/C VGND VGND VPWR VPWR _4424_/Y sky130_fd_sc_hd__nand3_4
XFILLER_132_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7143_ _7181_/CLK _7143_/D fanout499/X VGND VGND VPWR VPWR _7143_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_99_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4355_ _4819_/C _4781_/A _4935_/A VGND VGND VPWR VPWR _4355_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_113_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout427 _5203_/B VGND VGND VPWR VPWR _5535_/B sky130_fd_sc_hd__buf_12
X_3306_ _3546_/A hold68/X VGND VGND VPWR VPWR hold69/A sky130_fd_sc_hd__nor2_8
X_7074_ _7074_/CLK _7074_/D fanout501/X VGND VGND VPWR VPWR _7074_/Q sky130_fd_sc_hd__dfstp_1
Xfanout438 _5569_/A0 VGND VGND VPWR VPWR _5578_/A0 sky130_fd_sc_hd__clkbuf_4
X_4286_ _6396_/A0 hold540/X _4287_/S VGND VGND VPWR VPWR _4286_/X sky130_fd_sc_hd__mux2_1
Xfanout449 _5539_/A1 VGND VGND VPWR VPWR _6396_/A0 sky130_fd_sc_hd__buf_8
XFILLER_113_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6025_ _6025_/A _6025_/B _6025_/C _6025_/D VGND VGND VPWR VPWR _6026_/D sky130_fd_sc_hd__or4_1
X_3237_ _4570_/B VGND VGND VPWR VPWR _4667_/C sky130_fd_sc_hd__inv_4
XFILLER_86_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6927_ _7079_/CLK _6927_/D fanout517/X VGND VGND VPWR VPWR _6927_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_81_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6858_ _7110_/CLK _6858_/D fanout506/X VGND VGND VPWR VPWR _6858_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_120_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5809_ _6887_/Q _5846_/A2 _5848_/B1 _7047_/Q VGND VGND VPWR VPWR _5809_/X sky130_fd_sc_hd__a22o_1
X_6789_ _3927_/A1 _6789_/D _6440_/X VGND VGND VPWR VPWR _6789_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold470 _3981_/X VGND VGND VPWR VPWR hold39/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold481 _4299_/X VGND VGND VPWR VPWR _6745_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold492 _7045_/Q VGND VGND VPWR VPWR hold492/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1170 _4333_/X VGND VGND VPWR VPWR _6773_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1181 _5536_/X VGND VGND VPWR VPWR _7095_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1192 _5422_/X VGND VGND VPWR VPWR _6994_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_728 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4140_ hold484/X _6397_/A0 _4140_/S VGND VGND VPWR VPWR _4140_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4071_ hold977/X _6393_/A0 _4083_/S VGND VGND VPWR VPWR _4071_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4973_ _5140_/A _4973_/B VGND VGND VPWR VPWR _4979_/C sky130_fd_sc_hd__or2_1
X_6712_ _6725_/CLK _6712_/D fanout509/X VGND VGND VPWR VPWR _6712_/Q sky130_fd_sc_hd__dfrtp_4
X_3924_ _6575_/Q input78/X _3958_/B VGND VGND VPWR VPWR _3924_/X sky130_fd_sc_hd__mux2_8
XFILLER_20_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6643_ _7193_/CLK _6643_/D VGND VGND VPWR VPWR _6643_/Q sky130_fd_sc_hd__dfxtp_1
X_3855_ _6455_/Q _3856_/B _3854_/Y _3855_/B2 VGND VGND VPWR VPWR _3855_/X sky130_fd_sc_hd__o22a_1
XFILLER_164_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3786_ _6986_/Q _3298_/Y _3471_/Y _6761_/Q _3785_/X VGND VGND VPWR VPWR _3788_/C
+ sky130_fd_sc_hd__a221o_1
X_6574_ _6764_/CLK _6574_/D _6426_/A VGND VGND VPWR VPWR _6574_/Q sky130_fd_sc_hd__dfrtp_1
X_5525_ _5549_/A0 hold625/X _5528_/S VGND VGND VPWR VPWR _5525_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5456_ hold40/X hold119/X _5456_/S VGND VGND VPWR VPWR _5456_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4407_ _4621_/B _4538_/B VGND VGND VPWR VPWR _4436_/B sky130_fd_sc_hd__xnor2_2
XFILLER_160_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5387_ _5459_/A0 hold315/X _5393_/S VGND VGND VPWR VPWR _5387_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7126_ _7126_/CLK _7126_/D fanout524/X VGND VGND VPWR VPWR _7126_/Q sky130_fd_sc_hd__dfrtp_1
X_4338_ _4338_/A _4338_/B _4338_/C _4338_/D VGND VGND VPWR VPWR _4348_/B sky130_fd_sc_hd__and4_1
XFILLER_59_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4269_ hold785/X _6397_/A0 _4269_/S VGND VGND VPWR VPWR _4269_/X sky130_fd_sc_hd__mux2_1
X_7057_ _7102_/CLK _7057_/D fanout503/X VGND VGND VPWR VPWR _7057_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6008_ _6033_/A _6020_/C _6030_/C VGND VGND VPWR VPWR _6023_/C sky130_fd_sc_hd__and3_4
XFILLER_67_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_140 _3961_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_151 _6496_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_162 _6027_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_173 _5212_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_184 _3927_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_195 _5205_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3640_ _7012_/Q _5439_/A _4282_/A _6733_/Q VGND VGND VPWR VPWR _3640_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3571_ _6869_/Q _5277_/A _4159_/A _6624_/Q VGND VGND VPWR VPWR _3571_/X sky130_fd_sc_hd__a22o_1
X_5310_ _5550_/A0 hold573/X _5312_/S VGND VGND VPWR VPWR _5310_/X sky130_fd_sc_hd__mux2_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6290_ _6613_/Q _6023_/C _6020_/X _6708_/Q _6289_/X VGND VGND VPWR VPWR _6291_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_154_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5241_ hold96/A _5241_/B _6407_/B hold13/X VGND VGND VPWR VPWR hold14/A sky130_fd_sc_hd__or4_4
XFILLER_130_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5172_ _5172_/A _5172_/B _5172_/C _5172_/D VGND VGND VPWR VPWR _5183_/A sky130_fd_sc_hd__nor4_1
XFILLER_68_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4123_ _5583_/A0 hold329/X _4128_/S VGND VGND VPWR VPWR _4123_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput2 debug_oeb VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__clkbuf_1
X_4054_ hold793/X _5581_/A0 _4068_/S VGND VGND VPWR VPWR _4054_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_opt_1_0_csclk _7018_/CLK VGND VGND VPWR VPWR clkbuf_leaf_4_csclk/A sky130_fd_sc_hd__clkbuf_16
XFILLER_37_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4956_ _4997_/A _5035_/B _4935_/C _4944_/X _4916_/B VGND VGND VPWR VPWR _5163_/A
+ sky130_fd_sc_hd__o221a_1
X_3907_ _6318_/S _5592_/B VGND VGND VPWR VPWR _5651_/A sky130_fd_sc_hd__nor2_1
XFILLER_177_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4887_ _4885_/X _4887_/B _4887_/C _4887_/D VGND VGND VPWR VPWR _4890_/B sky130_fd_sc_hd__nand4b_1
XFILLER_165_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6626_ _7193_/CLK _6626_/D VGND VGND VPWR VPWR _6626_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3838_ _6541_/Q _3838_/B VGND VGND VPWR VPWR _3839_/B sky130_fd_sc_hd__nand2_1
XFILLER_192_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6557_ _7141_/CLK _6557_/D fanout504/X VGND VGND VPWR VPWR _6557_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_180_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3769_ _6490_/Q _3992_/A _5466_/A _7034_/Q _3768_/X VGND VGND VPWR VPWR _3769_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5508_ _5550_/A0 hold679/X _5510_/S VGND VGND VPWR VPWR _5508_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6488_ _7002_/CLK _6488_/D fanout498/X VGND VGND VPWR VPWR _6488_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_105_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5439_ _5439_/A _5571_/B VGND VGND VPWR VPWR _5447_/S sky130_fd_sc_hd__nand2_8
XFILLER_161_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7109_ _7133_/CLK _7109_/D fanout506/X VGND VGND VPWR VPWR _7109_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4810_ _4806_/X _4810_/B _4810_/C _4810_/D VGND VGND VPWR VPWR _4810_/X sky130_fd_sc_hd__and4b_1
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5790_ _6998_/Q _5656_/X _5671_/X _7062_/Q VGND VGND VPWR VPWR _5790_/X sky130_fd_sc_hd__a22o_1
XFILLER_178_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4741_ _4931_/B _4742_/C _4741_/C VGND VGND VPWR VPWR _4741_/X sky130_fd_sc_hd__and3_1
XFILLER_193_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4672_ _4672_/A _5021_/B VGND VGND VPWR VPWR _5128_/B sky130_fd_sc_hd__or2_1
XFILLER_186_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6411_ _6433_/A _6441_/B VGND VGND VPWR VPWR _6411_/X sky130_fd_sc_hd__and2_1
X_3623_ _3958_/A _4104_/A _4210_/A _6667_/Q _3612_/X VGND VGND VPWR VPWR _3627_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_174_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6342_ _6600_/Q _6046_/B _6332_/X _6341_/X _3195_/Y VGND VGND VPWR VPWR _6342_/X
+ sky130_fd_sc_hd__o221a_2
X_3554_ _6744_/Q _4294_/A _4034_/A _6529_/Q VGND VGND VPWR VPWR _3554_/X sky130_fd_sc_hd__a22o_1
XFILLER_142_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6273_ _6703_/Q _6336_/A2 _6033_/X _7209_/Q VGND VGND VPWR VPWR _6273_/X sky130_fd_sc_hd__a22o_1
X_3485_ _3525_/A _3538_/B VGND VGND VPWR VPWR _6392_/A sky130_fd_sc_hd__nor2_8
XFILLER_143_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5224_ _5521_/A0 _5224_/A1 _5224_/S VGND VGND VPWR VPWR _5224_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5155_ _5155_/A _5155_/B _5155_/C _4681_/X VGND VGND VPWR VPWR _5178_/C sky130_fd_sc_hd__or4b_1
XFILLER_84_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4106_ _6394_/A0 _4106_/A1 _4110_/S VGND VGND VPWR VPWR _4106_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5086_ _5156_/B _5178_/A _5106_/C _5086_/D VGND VGND VPWR VPWR _5087_/B sky130_fd_sc_hd__or4_1
XFILLER_110_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4037_ _4037_/A0 _6395_/A0 _4039_/S VGND VGND VPWR VPWR _4037_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5988_ _6014_/A _6040_/B _6040_/C VGND VGND VPWR VPWR _5988_/X sky130_fd_sc_hd__and3_4
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4939_ _5065_/D _5124_/C _4939_/C VGND VGND VPWR VPWR _4961_/A sky130_fd_sc_hd__or3_1
XFILLER_178_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_40 _3580_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_51 _5016_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_62 _5667_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_73 _5968_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_84 _6930_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6609_ _6725_/CLK _6609_/D fanout509/X VGND VGND VPWR VPWR _6609_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_192_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_95 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput180 _3220_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[14] sky130_fd_sc_hd__buf_12
XFILLER_121_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput191 _3210_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[24] sky130_fd_sc_hd__buf_12
XFILLER_0_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_44_csclk _6931_/CLK VGND VGND VPWR VPWR _7031_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_140_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3270_ hold18/X _3301_/C VGND VGND VPWR VPWR hold19/A sky130_fd_sc_hd__nand2_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_59_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7080_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_97_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6960_ _7141_/CLK _6960_/D fanout504/X VGND VGND VPWR VPWR _6960_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_54_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5911_ _6636_/Q _5655_/X _5656_/X _6743_/Q VGND VGND VPWR VPWR _5911_/X sky130_fd_sc_hd__a22o_1
XFILLER_46_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6891_ _7012_/CLK _6891_/D fanout505/X VGND VGND VPWR VPWR _6891_/Q sky130_fd_sc_hd__dfstp_1
X_5842_ _6865_/Q _5688_/X _5696_/X _7041_/Q _5841_/X VGND VGND VPWR VPWR _5847_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5773_ _5650_/A _7164_/Q _5772_/X VGND VGND VPWR VPWR _5773_/X sky130_fd_sc_hd__a21o_1
XFILLER_166_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4724_ _4724_/A _4724_/B VGND VGND VPWR VPWR _4742_/C sky130_fd_sc_hd__nor2_1
XFILLER_147_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4655_ _4832_/B _4659_/B VGND VGND VPWR VPWR _5177_/B sky130_fd_sc_hd__nor2_2
XFILLER_135_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput60 mgmt_gpio_in[31] VGND VGND VPWR VPWR input60/X sky130_fd_sc_hd__clkbuf_1
X_3606_ _6892_/Q _5304_/A _5268_/A _6860_/Q VGND VGND VPWR VPWR _3606_/X sky130_fd_sc_hd__a22o_1
Xhold800 _4109_/X VGND VGND VPWR VPWR _6578_/D sky130_fd_sc_hd__dlygate4sd3_1
Xinput71 mgmt_gpio_in[8] VGND VGND VPWR VPWR input71/X sky130_fd_sc_hd__buf_2
Xhold811 _6868_/Q VGND VGND VPWR VPWR hold811/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput82 spi_sdoenb VGND VGND VPWR VPWR input82/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4586_ _4814_/A _5018_/C VGND VGND VPWR VPWR _4677_/B sky130_fd_sc_hd__or2_4
XFILLER_190_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput93 trap VGND VGND VPWR VPWR input93/X sky130_fd_sc_hd__buf_4
Xhold822 _5446_/X VGND VGND VPWR VPWR _7016_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold833 _5356_/X VGND VGND VPWR VPWR _6936_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6325_ _6659_/Q _6022_/B _6016_/X _6685_/Q VGND VGND VPWR VPWR _6325_/X sky130_fd_sc_hd__a22o_1
Xhold844 _7043_/Q VGND VGND VPWR VPWR hold844/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3537_ _7038_/Q _5466_/A _4312_/A _6760_/Q _3535_/X VGND VGND VPWR VPWR _3541_/C
+ sky130_fd_sc_hd__a221o_2
Xhold855 _5307_/X VGND VGND VPWR VPWR _6892_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold866 hold866/A VGND VGND VPWR VPWR hold866/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold877 _5219_/X VGND VGND VPWR VPWR _6817_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 _6915_/Q VGND VGND VPWR VPWR hold888/X sky130_fd_sc_hd__dlygate4sd3_1
X_6256_ _6712_/Q _6009_/X _6038_/Y _6722_/Q _6255_/X VGND VGND VPWR VPWR _6257_/D
+ sky130_fd_sc_hd__a221o_1
Xhold899 _4003_/X VGND VGND VPWR VPWR _6499_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3468_ _3468_/A _3468_/B _3468_/C _3468_/D VGND VGND VPWR VPWR _3543_/A sky130_fd_sc_hd__or4_1
X_5207_ hold391/X _5555_/A0 _5209_/S VGND VGND VPWR VPWR _5207_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6187_ _7016_/Q _5998_/Y wire412/X _6920_/Q _6186_/X VGND VGND VPWR VPWR _6192_/B
+ sky130_fd_sc_hd__a221o_1
X_3399_ _7101_/Q _5535_/A hold69/A _7141_/Q _3398_/X VGND VGND VPWR VPWR _3399_/X
+ sky130_fd_sc_hd__a221o_1
Xhold1500 _7160_/Q VGND VGND VPWR VPWR _5647_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_191_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1511 _7181_/Q VGND VGND VPWR VPWR _6196_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1522 _3861_/X VGND VGND VPWR VPWR _6451_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1533 _6457_/Q VGND VGND VPWR VPWR _3845_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5138_ _5148_/C _5138_/B VGND VGND VPWR VPWR _5139_/D sky130_fd_sc_hd__and2b_1
Xhold1544 _6825_/Q VGND VGND VPWR VPWR hold1544/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1555 _6473_/Q VGND VGND VPWR VPWR _3798_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1566 _6583_/Q VGND VGND VPWR VPWR hold472/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1577 _6588_/Q VGND VGND VPWR VPWR hold977/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1588 _6554_/Q VGND VGND VPWR VPWR hold1588/X sky130_fd_sc_hd__dlygate4sd3_1
X_5069_ _5069_/A _5160_/A VGND VGND VPWR VPWR _5104_/B sky130_fd_sc_hd__nor2_1
Xhold1599 _7148_/Q VGND VGND VPWR VPWR _5611_/S sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_40_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4440_ _4441_/A _4453_/C VGND VGND VPWR VPWR _4516_/B sky130_fd_sc_hd__nor2_4
XFILLER_156_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold107 _3329_/Y VGND VGND VPWR VPWR hold107/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold118 _5293_/X VGND VGND VPWR VPWR _6880_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 _6567_/Q VGND VGND VPWR VPWR hold129/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4371_ _4846_/A _4570_/B VGND VGND VPWR VPWR _4781_/B sky130_fd_sc_hd__nand2_2
XFILLER_171_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6110_ _6110_/A _6110_/B VGND VGND VPWR VPWR _6110_/X sky130_fd_sc_hd__or2_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3322_ _5241_/B _3530_/B VGND VGND VPWR VPWR _5385_/A sky130_fd_sc_hd__nor2_8
XFILLER_140_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7090_ _7209_/CLK _7090_/D fanout485/X VGND VGND VPWR VPWR _7090_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6041_ _6962_/Q _6025_/D _6212_/B1 _7042_/Q VGND VGND VPWR VPWR _6041_/X sky130_fd_sc_hd__a22o_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3253_ _3248_/A hold72/X _3818_/A VGND VGND VPWR VPWR _3253_/X sky130_fd_sc_hd__a21bo_1
XFILLER_98_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3184_ _6472_/Q VGND VGND VPWR VPWR _3184_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6943_ _7049_/CLK _6943_/D fanout522/X VGND VGND VPWR VPWR _6943_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6874_ _7135_/CLK _6874_/D fanout519/X VGND VGND VPWR VPWR _6874_/Q sky130_fd_sc_hd__dfstp_2
X_5825_ _5825_/A _5825_/B _5825_/C _5825_/D VGND VGND VPWR VPWR _5825_/X sky130_fd_sc_hd__or4_1
XFILLER_50_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5756_ _6885_/Q _5846_/A2 _5848_/B1 _7045_/Q VGND VGND VPWR VPWR _5756_/X sky130_fd_sc_hd__a22o_1
X_4707_ _4707_/A _4707_/B VGND VGND VPWR VPWR _4850_/B sky130_fd_sc_hd__or2_1
XFILLER_148_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5687_ _6906_/Q _5685_/X _5686_/X _7010_/Q _5684_/X VGND VGND VPWR VPWR _5708_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_162_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4638_ _4814_/A _4638_/B VGND VGND VPWR VPWR _4689_/B sky130_fd_sc_hd__or2_4
XFILLER_116_550 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold630 _4281_/X VGND VGND VPWR VPWR _6730_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4569_ _4846_/B _4569_/B VGND VGND VPWR VPWR _4569_/Y sky130_fd_sc_hd__nor2_1
XFILLER_150_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold641 _6918_/Q VGND VGND VPWR VPWR hold641/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold652 _5504_/X VGND VGND VPWR VPWR _7067_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap371 _5484_/A VGND VGND VPWR VPWR _3684_/B1 sky130_fd_sc_hd__buf_6
Xhold663 _6894_/Q VGND VGND VPWR VPWR hold663/X sky130_fd_sc_hd__dlygate4sd3_1
X_6308_ _6719_/Q _6308_/A2 _6338_/B1 _6769_/Q _6296_/X VGND VGND VPWR VPWR _6308_/X
+ sky130_fd_sc_hd__a221o_1
Xmax_cap382 hold49/X VGND VGND VPWR VPWR _3530_/B sky130_fd_sc_hd__buf_12
Xhold674 _5463_/X VGND VGND VPWR VPWR _7031_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap393 _6025_/C VGND VGND VPWR VPWR _6322_/B1 sky130_fd_sc_hd__buf_8
Xhold685 _6674_/Q VGND VGND VPWR VPWR hold685/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold696 _5534_/X VGND VGND VPWR VPWR _7094_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6239_ _7090_/Q _5642_/X _5992_/X _6675_/Q VGND VGND VPWR VPWR _6239_/X sky130_fd_sc_hd__a22o_1
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1330 hold1330/A VGND VGND VPWR VPWR wb_dat_o[13] sky130_fd_sc_hd__buf_12
Xhold1341 _4184_/A0 VGND VGND VPWR VPWR hold1341/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1352 hold1352/A VGND VGND VPWR VPWR wb_dat_o[4] sky130_fd_sc_hd__buf_12
XFILLER_85_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1363 _4166_/A0 VGND VGND VPWR VPWR hold1363/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1374 _5243_/X VGND VGND VPWR VPWR hold15/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1385 _6609_/Q VGND VGND VPWR VPWR _4145_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1396 _6632_/Q VGND VGND VPWR VPWR hold1396/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3940_ _7161_/Q _6814_/Q _6818_/Q VGND VGND VPWR VPWR _3940_/X sky130_fd_sc_hd__mux2_2
XFILLER_63_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3871_ input58/X _3840_/S _3870_/X _3914_/A1 VGND VGND VPWR VPWR _6444_/D sky130_fd_sc_hd__a22o_1
XFILLER_176_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5610_ _6562_/Q _6564_/Q VGND VGND VPWR VPWR _5610_/X sky130_fd_sc_hd__or2_1
XFILLER_177_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6590_ _7141_/CLK _6590_/D fanout504/X VGND VGND VPWR VPWR _6590_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_31_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5541_ hold261/X hold127/X _5543_/S VGND VGND VPWR VPWR _5541_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5472_ hold609/X _5550_/A0 _5474_/S VGND VGND VPWR VPWR _5472_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7211_ _7211_/CLK _7211_/D fanout485/X VGND VGND VPWR VPWR _7211_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_160_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4423_ _4758_/A _4758_/B _4758_/C VGND VGND VPWR VPWR _4485_/A sky130_fd_sc_hd__and3_4
X_7142_ _7142_/CLK hold71/X fanout525/X VGND VGND VPWR VPWR _7142_/Q sky130_fd_sc_hd__dfrtp_1
X_4354_ _4354_/A _4354_/B VGND VGND VPWR VPWR _4935_/B sky130_fd_sc_hd__nand2_1
XFILLER_99_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3305_ hold67/X _3330_/B VGND VGND VPWR VPWR hold68/A sky130_fd_sc_hd__nand2_8
Xfanout428 _5385_/B VGND VGND VPWR VPWR _5313_/B sky130_fd_sc_hd__buf_12
XFILLER_59_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7073_ _7134_/CLK _7073_/D fanout525/X VGND VGND VPWR VPWR _7073_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout439 hold101/X VGND VGND VPWR VPWR _5569_/A0 sky130_fd_sc_hd__buf_12
X_4285_ _6395_/A0 _4285_/A1 _4287_/S VGND VGND VPWR VPWR _4285_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6024_ _6024_/A _6024_/B _6024_/C _6024_/D VGND VGND VPWR VPWR _6026_/C sky130_fd_sc_hd__or4_1
XFILLER_100_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3236_ _4846_/A VGND VGND VPWR VPWR _4420_/A sky130_fd_sc_hd__clkinv_2
XFILLER_39_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6926_ _7082_/CLK _6926_/D _3873_/A VGND VGND VPWR VPWR _6926_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_81_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6857_ _6992_/CLK _6857_/D fanout517/X VGND VGND VPWR VPWR _6857_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5808_ _7055_/Q _5699_/X _5702_/X _6983_/Q _5807_/X VGND VGND VPWR VPWR _5813_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_167_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6788_ _3487_/B2 _6788_/D _6439_/X VGND VGND VPWR VPWR _6788_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_183_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5739_ _6892_/Q _5655_/X _5663_/X _7020_/Q _5738_/X VGND VGND VPWR VPWR _5740_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold460 _4334_/X VGND VGND VPWR VPWR _6774_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold471 _3991_/X VGND VGND VPWR VPWR _6489_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold482 _6478_/Q VGND VGND VPWR VPWR hold482/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold493 _5479_/X VGND VGND VPWR VPWR _7045_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1160 _3986_/X VGND VGND VPWR VPWR _6484_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1171 _6807_/Q VGND VGND VPWR VPWR _5206_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1182 _6483_/Q VGND VGND VPWR VPWR _3985_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1193 _6500_/Q VGND VGND VPWR VPWR _4004_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_2__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR _3487_/B2
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_154_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4070_ _4120_/B _6407_/B _4052_/X _4085_/S _4330_/B VGND VGND VPWR VPWR _4086_/S
+ sky130_fd_sc_hd__o221a_4
XFILLER_110_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4972_ _4783_/A _4794_/C _4971_/Y _4781_/Y _5013_/A VGND VGND VPWR VPWR _4973_/B
+ sky130_fd_sc_hd__o32ai_4
XFILLER_17_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6711_ _6725_/CLK _6711_/D fanout509/X VGND VGND VPWR VPWR _6711_/Q sky130_fd_sc_hd__dfrtp_4
X_3923_ _6574_/Q input80/X _3958_/B VGND VGND VPWR VPWR _3923_/X sky130_fd_sc_hd__mux2_8
XFILLER_20_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6642_ _7193_/CLK _6642_/D VGND VGND VPWR VPWR _6642_/Q sky130_fd_sc_hd__dfxtp_1
X_3854_ _3856_/B _3858_/B VGND VGND VPWR VPWR _3854_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6573_ _7140_/CLK _6573_/D fanout522/X VGND VGND VPWR VPWR _6573_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3785_ input93/X _3256_/Y _3286_/Y _4282_/A _6731_/Q VGND VGND VPWR VPWR _3785_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_164_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5524_ _5584_/A0 hold439/X _5528_/S VGND VGND VPWR VPWR _5524_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5455_ _5587_/A0 hold936/X _5456_/S VGND VGND VPWR VPWR _5455_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4406_ _4560_/A _4731_/C _4731_/B VGND VGND VPWR VPWR _4453_/A sky130_fd_sc_hd__nand3_2
X_5386_ _5521_/A0 _5386_/A1 _5393_/S VGND VGND VPWR VPWR _5386_/X sky130_fd_sc_hd__mux2_1
XFILLER_120_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7125_ _7134_/CLK _7125_/D fanout524/X VGND VGND VPWR VPWR _7125_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_101_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4337_ _4337_/A _4337_/B _4337_/C _4337_/D VGND VGND VPWR VPWR _4348_/A sky130_fd_sc_hd__and4_1
XFILLER_101_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7056_ _7102_/CLK _7056_/D fanout503/X VGND VGND VPWR VPWR _7056_/Q sky130_fd_sc_hd__dfrtp_2
X_4268_ hold577/X _6396_/A0 _4269_/S VGND VGND VPWR VPWR _4268_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6007_ _6019_/A _6038_/B VGND VGND VPWR VPWR _6007_/Y sky130_fd_sc_hd__nor2_8
X_3219_ _6965_/Q VGND VGND VPWR VPWR _3219_/Y sky130_fd_sc_hd__inv_2
X_4199_ _4199_/A0 _5476_/A0 _4203_/S VGND VGND VPWR VPWR _4199_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6909_ _7138_/CLK _6909_/D fanout520/X VGND VGND VPWR VPWR _6909_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold290 _4143_/X VGND VGND VPWR VPWR _6607_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_130 input84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_141 input38/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_152 _6497_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_163 _6329_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_174 _3937_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_185 _3927_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_196 _3573_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3570_ _6973_/Q _5394_/A hold31/A _6877_/Q _3569_/X VGND VGND VPWR VPWR _3573_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5240_ _5579_/A0 hold399/X _5240_/S VGND VGND VPWR VPWR _5240_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5171_ _5171_/A _5171_/B VGND VGND VPWR VPWR _5172_/D sky130_fd_sc_hd__nor2_1
X_4122_ _5531_/A1 hold922/X _4128_/S VGND VGND VPWR VPWR _4122_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4053_ _4111_/B _6407_/B _4052_/X _3308_/Y _5580_/B VGND VGND VPWR VPWR _4069_/S
+ sky130_fd_sc_hd__o221a_4
Xinput3 debug_out VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4955_ _4462_/Y _4933_/Y _4828_/X VGND VGND VPWR VPWR _5123_/A sky130_fd_sc_hd__a21oi_1
XFILLER_51_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3906_ _6019_/A _6018_/A VGND VGND VPWR VPWR _3906_/X sky130_fd_sc_hd__or2_1
XFILLER_189_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4886_ _4424_/Y _4872_/B _4758_/Y _4504_/B VGND VGND VPWR VPWR _4887_/B sky130_fd_sc_hd__o211a_1
X_6625_ _6679_/CLK _6625_/D fanout511/X VGND VGND VPWR VPWR _6625_/Q sky130_fd_sc_hd__dfrtp_2
X_3837_ _3850_/B _3837_/A2 _3836_/Y _6461_/Q VGND VGND VPWR VPWR _6461_/D sky130_fd_sc_hd__a31o_1
X_6556_ _7141_/CLK _6556_/D fanout504/X VGND VGND VPWR VPWR _6556_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3768_ _6506_/Q _4010_/A _4022_/A _6516_/Q VGND VGND VPWR VPWR _3768_/X sky130_fd_sc_hd__a22o_1
X_5507_ _5549_/A0 hold643/X _5510_/S VGND VGND VPWR VPWR _5507_/X sky130_fd_sc_hd__mux2_1
XFILLER_180_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6487_ _6825_/CLK _6487_/D fanout498/X VGND VGND VPWR VPWR _6487_/Q sky130_fd_sc_hd__dfstp_1
X_3699_ _6979_/Q _5403_/A _6392_/A _7208_/Q VGND VGND VPWR VPWR _3699_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5438_ _5552_/A0 hold779/X _5438_/S VGND VGND VPWR VPWR _5438_/X sky130_fd_sc_hd__mux2_1
Xoutput340 hold1355/X VGND VGND VPWR VPWR hold1356/A sky130_fd_sc_hd__buf_12
XFILLER_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5369_ _5573_/A0 hold838/X _5375_/S VGND VGND VPWR VPWR _5369_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7108_ _7108_/CLK _7108_/D fanout523/X VGND VGND VPWR VPWR _7108_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7039_ _7079_/CLK _7039_/D fanout516/X VGND VGND VPWR VPWR _7039_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_28_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire412 _6027_/C VGND VGND VPWR VPWR wire412/X sky130_fd_sc_hd__buf_12
XFILLER_183_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4740_ _4931_/B _4742_/C VGND VGND VPWR VPWR _4740_/Y sky130_fd_sc_hd__nand2_1
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4671_ _4672_/A _5021_/B VGND VGND VPWR VPWR _5158_/A sky130_fd_sc_hd__nor2_2
XFILLER_186_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6410_ _6433_/A _6440_/B VGND VGND VPWR VPWR _6410_/X sky130_fd_sc_hd__and2_1
X_3622_ _6728_/Q _4276_/A _3616_/X _3620_/X _3621_/X VGND VGND VPWR VPWR _3633_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_147_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6341_ _6341_/A _6341_/B _6341_/C _6341_/D VGND VGND VPWR VPWR _6341_/X sky130_fd_sc_hd__or4_1
X_3553_ _7005_/Q _5430_/A _4282_/A _6734_/Q VGND VGND VPWR VPWR _3553_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6272_ _6533_/Q _6272_/B VGND VGND VPWR VPWR _6272_/X sky130_fd_sc_hd__and2_1
X_3484_ _3484_/A _3484_/B _3484_/C _3484_/D VGND VGND VPWR VPWR _3543_/B sky130_fd_sc_hd__or4_1
XFILLER_170_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5223_ _5223_/A _5580_/B VGND VGND VPWR VPWR _5224_/S sky130_fd_sc_hd__nand2_1
XFILLER_102_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5154_ _5076_/B _5021_/B _5017_/A VGND VGND VPWR VPWR _5155_/C sky130_fd_sc_hd__a21oi_1
X_4105_ _6393_/A0 _4105_/A1 _4110_/S VGND VGND VPWR VPWR _4105_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5085_ _4420_/A _5106_/A _5109_/C _5107_/B _5153_/B VGND VGND VPWR VPWR _5086_/D
+ sky130_fd_sc_hd__a2111o_1
XFILLER_56_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4036_ _4036_/A0 _6394_/A0 _4039_/S VGND VGND VPWR VPWR _4036_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5987_ _7155_/Q _7156_/Q VGND VGND VPWR VPWR _6040_/C sky130_fd_sc_hd__and2b_2
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4938_ _4605_/A _4428_/B _4957_/B _5177_/B _4506_/Y VGND VGND VPWR VPWR _4939_/C
+ sky130_fd_sc_hd__a311o_1
XFILLER_178_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_30 _3481_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_41 _3620_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4869_ _4930_/C _4868_/X _4930_/A VGND VGND VPWR VPWR _4928_/B sky130_fd_sc_hd__o21ba_1
XFILLER_20_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_52 _5285_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_63 _5671_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6608_ _6725_/CLK _6608_/D fanout509/X VGND VGND VPWR VPWR _6608_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA_74 _6045_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_85 _6957_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_96 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6539_ _6707_/CLK _6539_/D _6432_/A VGND VGND VPWR VPWR _6539_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_106_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput181 _3219_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[15] sky130_fd_sc_hd__buf_12
Xoutput192 _3209_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[25] sky130_fd_sc_hd__buf_12
XFILLER_153_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5910_ _6608_/Q _5688_/X _5909_/X VGND VGND VPWR VPWR _5913_/C sky130_fd_sc_hd__a21o_1
X_6890_ _7123_/CLK _6890_/D fanout519/X VGND VGND VPWR VPWR _6890_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5841_ _6961_/Q _5659_/X _5705_/X _6945_/Q VGND VGND VPWR VPWR _5841_/X sky130_fd_sc_hd__a22o_1
XFILLER_62_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5772_ _6845_/Q _5691_/Y _5770_/X _5771_/X _6318_/S VGND VGND VPWR VPWR _5772_/X
+ sky130_fd_sc_hd__o221a_2
X_4723_ _4650_/Y _4722_/X _6362_/A _4648_/Y VGND VGND VPWR VPWR _4723_/X sky130_fd_sc_hd__a211o_1
XFILLER_175_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4654_ _4654_/A _4654_/B _4390_/A VGND VGND VPWR VPWR _5021_/C sky130_fd_sc_hd__or3b_4
X_3605_ _7097_/Q _5535_/A _5250_/A _6844_/Q VGND VGND VPWR VPWR _3605_/X sky130_fd_sc_hd__a22o_1
XFILLER_174_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput50 mgmt_gpio_in[22] VGND VGND VPWR VPWR input50/X sky130_fd_sc_hd__buf_2
XFILLER_190_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput61 mgmt_gpio_in[32] VGND VGND VPWR VPWR input61/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold801 _6848_/Q VGND VGND VPWR VPWR hold801/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput72 mgmt_gpio_in[9] VGND VGND VPWR VPWR input72/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4585_ _4588_/A _4935_/A _4341_/X VGND VGND VPWR VPWR _5018_/C sky130_fd_sc_hd__or3b_4
Xhold812 _5280_/X VGND VGND VPWR VPWR _6868_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_174_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold823 _6856_/Q VGND VGND VPWR VPWR hold823/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput83 spimemio_flash_clk VGND VGND VPWR VPWR input83/X sky130_fd_sc_hd__buf_2
Xinput94 uart_enabled VGND VGND VPWR VPWR _3957_/B sky130_fd_sc_hd__clkbuf_1
Xhold834 _7072_/Q VGND VGND VPWR VPWR hold834/X sky130_fd_sc_hd__dlygate4sd3_1
X_6324_ _6525_/Q _5994_/X _5998_/Y _6765_/Q _6323_/X VGND VGND VPWR VPWR _6331_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3536_ _3536_/A _3726_/B VGND VGND VPWR VPWR _4312_/A sky130_fd_sc_hd__nor2_2
Xhold845 _5477_/X VGND VGND VPWR VPWR _7043_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold856 _6667_/Q VGND VGND VPWR VPWR hold856/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold867 _5560_/X VGND VGND VPWR VPWR _7117_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold878 _7120_/Q VGND VGND VPWR VPWR hold878/X sky130_fd_sc_hd__dlygate4sd3_1
X_6255_ _6702_/Q _6336_/A2 _6033_/X _7208_/Q VGND VGND VPWR VPWR _6255_/X sky130_fd_sc_hd__a22o_1
Xhold889 _5333_/X VGND VGND VPWR VPWR _6915_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3467_ _6685_/Q hold58/A _4210_/A _6669_/Q _3464_/X VGND VGND VPWR VPWR _3468_/D
+ sky130_fd_sc_hd__a221o_1
X_5206_ _5206_/A0 _5536_/A1 _5209_/S VGND VGND VPWR VPWR _5206_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6186_ _7032_/Q _6049_/B _6272_/B _7072_/Q VGND VGND VPWR VPWR _6186_/X sky130_fd_sc_hd__a22o_1
X_3398_ _7000_/Q _3300_/Y _3992_/A _6496_/Q VGND VGND VPWR VPWR _3398_/X sky130_fd_sc_hd__a22o_1
Xhold1501 _7165_/Q VGND VGND VPWR VPWR _5794_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1512 _6446_/Q VGND VGND VPWR VPWR _3866_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5137_ _5148_/A _5151_/B _5148_/D _5137_/D VGND VGND VPWR VPWR _5138_/B sky130_fd_sc_hd__or4_1
Xhold1523 _7166_/Q VGND VGND VPWR VPWR _5795_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1534 _6444_/Q VGND VGND VPWR VPWR _3914_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1545 hold91/A VGND VGND VPWR VPWR _3810_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1556 _7171_/Q VGND VGND VPWR VPWR _5904_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1567 _6589_/Q VGND VGND VPWR VPWR hold922/A sky130_fd_sc_hd__dlygate4sd3_1
X_5068_ _5068_/A _5068_/B VGND VGND VPWR VPWR _5160_/A sky130_fd_sc_hd__or2_1
XFILLER_84_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1578 _6840_/Q VGND VGND VPWR VPWR hold123/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1589 _7147_/Q VGND VGND VPWR VPWR _5608_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4019_ _4327_/A1 hold870/X _4021_/S VGND VGND VPWR VPWR _4019_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold108 _5493_/Y VGND VGND VPWR VPWR _5501_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_156_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold119 _7025_/Q VGND VGND VPWR VPWR hold119/X sky130_fd_sc_hd__dlygate4sd3_1
X_4370_ _4745_/A _5076_/A _6700_/Q VGND VGND VPWR VPWR _4930_/A sky130_fd_sc_hd__o21ai_1
XFILLER_125_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3321_ _3536_/A hold68/X VGND VGND VPWR VPWR _5511_/A sky130_fd_sc_hd__nor2_8
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ _6040_/A _6040_/B _6040_/C VGND VGND VPWR VPWR _6040_/X sky130_fd_sc_hd__and3_4
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3252_ _6468_/Q _3252_/B VGND VGND VPWR VPWR _3818_/A sky130_fd_sc_hd__nand2_1
XFILLER_140_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6942_ _7123_/CLK _6942_/D _6407_/A VGND VGND VPWR VPWR _6942_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6873_ _6992_/CLK _6873_/D fanout517/X VGND VGND VPWR VPWR _6873_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_62_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5824_ _6896_/Q _5655_/X _5671_/X _7064_/Q _5823_/X VGND VGND VPWR VPWR _5825_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_179_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5755_ _6981_/Q _5702_/X _5706_/X _6501_/Q VGND VGND VPWR VPWR _5755_/X sky130_fd_sc_hd__a22o_1
X_4706_ _4707_/A _4683_/B _4863_/B _4705_/X VGND VGND VPWR VPWR _4708_/C sky130_fd_sc_hd__o211a_1
X_5686_ _7152_/Q _5700_/C _5703_/C VGND VGND VPWR VPWR _5686_/X sky130_fd_sc_hd__and3_4
XFILLER_148_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4637_ _5013_/A _5036_/A _5076_/B _5027_/A _4636_/X VGND VGND VPWR VPWR _4642_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_190_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold620 _5416_/X VGND VGND VPWR VPWR _6989_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 _6740_/Q VGND VGND VPWR VPWR hold631/X sky130_fd_sc_hd__dlygate4sd3_1
X_4568_ _4666_/B _5016_/A VGND VGND VPWR VPWR _4568_/X sky130_fd_sc_hd__or2_1
XFILLER_162_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap350 hold30/X VGND VGND VPWR VPWR hold31/A sky130_fd_sc_hd__buf_8
XFILLER_116_562 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold642 _5336_/X VGND VGND VPWR VPWR _6918_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold653 hold653/A VGND VGND VPWR VPWR hold653/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap361 _6168_/A VGND VGND VPWR VPWR _6217_/A sky130_fd_sc_hd__clkbuf_2
Xmax_cap372 _3326_/Y VGND VGND VPWR VPWR _5457_/A sky130_fd_sc_hd__buf_6
X_6307_ _6534_/Q _6272_/B _6302_/X _6304_/X _6306_/X VGND VGND VPWR VPWR _6307_/X
+ sky130_fd_sc_hd__a2111o_1
X_3519_ hold21/X _3525_/B VGND VGND VPWR VPWR _4141_/A sky130_fd_sc_hd__nor2_4
Xhold664 _5309_/X VGND VGND VPWR VPWR _6894_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold675 _6942_/Q VGND VGND VPWR VPWR hold675/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 _4221_/X VGND VGND VPWR VPWR _6674_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4499_ _4420_/A _4570_/B _4498_/X _4489_/X _4484_/X VGND VGND VPWR VPWR _4503_/D
+ sky130_fd_sc_hd__o311a_1
Xhold697 _6690_/Q VGND VGND VPWR VPWR hold697/X sky130_fd_sc_hd__dlygate4sd3_1
X_6238_ _6606_/Q _6326_/A2 _6021_/Y _6621_/Q _6237_/X VGND VGND VPWR VPWR _6241_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6169_ _6847_/Q _6046_/B _6156_/X _6168_/X _6318_/S VGND VGND VPWR VPWR _6169_/X
+ sky130_fd_sc_hd__o221a_2
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1320 hold1320/A VGND VGND VPWR VPWR wb_dat_o[23] sky130_fd_sc_hd__buf_12
Xhold1331 hold1411/X VGND VGND VPWR VPWR hold1331/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1342 hold1342/A VGND VGND VPWR VPWR wb_dat_o[11] sky130_fd_sc_hd__buf_12
XFILLER_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1353 _6351_/A0 VGND VGND VPWR VPWR hold1353/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1364 hold1364/A VGND VGND VPWR VPWR wb_dat_o[16] sky130_fd_sc_hd__buf_12
XFILLER_57_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1375 _7142_/Q VGND VGND VPWR VPWR _5588_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1386 _7049_/Q VGND VGND VPWR VPWR _5483_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1397 _6646_/Q VGND VGND VPWR VPWR hold1397/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_43_csclk _6931_/CLK VGND VGND VPWR VPWR _7065_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_58_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7102_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_185_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3870_ _6471_/Q _6445_/Q _3839_/B VGND VGND VPWR VPWR _3870_/X sky130_fd_sc_hd__a21o_1
XFILLER_177_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5540_ hold259/X _5558_/A0 _5543_/S VGND VGND VPWR VPWR _5540_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5471_ hold201/X _5558_/A0 _5474_/S VGND VGND VPWR VPWR _5471_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7210_ _7211_/CLK _7210_/D fanout485/X VGND VGND VPWR VPWR _7210_/Q sky130_fd_sc_hd__dfrtp_4
X_4422_ _4758_/A _4758_/C VGND VGND VPWR VPWR _4441_/A sky130_fd_sc_hd__nand2_1
X_7141_ _7141_/CLK _7141_/D fanout504/X VGND VGND VPWR VPWR _7141_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_132_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4353_ _4341_/X _4781_/A _4588_/A VGND VGND VPWR VPWR _4354_/B sky130_fd_sc_hd__a21o_1
X_3304_ _3731_/A _3528_/B VGND VGND VPWR VPWR _3304_/Y sky130_fd_sc_hd__nor2_4
X_7072_ _7098_/CLK _7072_/D fanout506/X VGND VGND VPWR VPWR _7072_/Q sky130_fd_sc_hd__dfrtp_1
X_4284_ _6394_/A0 _4284_/A1 _4287_/S VGND VGND VPWR VPWR _4284_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout429 _5203_/B VGND VGND VPWR VPWR _5580_/B sky130_fd_sc_hd__buf_12
XFILLER_140_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6023_ _6023_/A _6023_/B _6023_/C _6023_/D VGND VGND VPWR VPWR _6026_/B sky130_fd_sc_hd__or4_1
X_3235_ _7152_/Q VGND VGND VPWR VPWR _5960_/B sky130_fd_sc_hd__clkinv_8
XFILLER_101_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6925_ _6925_/CLK _6925_/D fanout516/X VGND VGND VPWR VPWR _6925_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_82_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6856_ _6977_/CLK _6856_/D fanout506/X VGND VGND VPWR VPWR _6856_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_120_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5807_ _6879_/Q _5667_/X _5675_/X _6967_/Q VGND VGND VPWR VPWR _5807_/X sky130_fd_sc_hd__a22o_1
XFILLER_167_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3999_ hold243/X _5569_/A0 _4000_/S VGND VGND VPWR VPWR _3999_/X sky130_fd_sc_hd__mux2_1
X_6787_ _3487_/B2 _6787_/D _6438_/X VGND VGND VPWR VPWR _6787_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_183_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5738_ _6988_/Q _5697_/X _5705_/X _6940_/Q VGND VGND VPWR VPWR _5738_/X sky130_fd_sc_hd__a22o_1
XFILLER_129_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5669_ _7150_/Q _7151_/Q VGND VGND VPWR VPWR _5699_/C sky130_fd_sc_hd__and2b_2
XFILLER_136_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold450 _5362_/X VGND VGND VPWR VPWR _6941_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 _6664_/Q VGND VGND VPWR VPWR hold461/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold472 hold472/A VGND VGND VPWR VPWR hold472/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold483 _3976_/X VGND VGND VPWR VPWR _6478_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 _6663_/Q VGND VGND VPWR VPWR hold494/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1150 _5190_/X VGND VGND VPWR VPWR _6795_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_161_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1161 _6732_/Q VGND VGND VPWR VPWR _4284_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1172 _5206_/X VGND VGND VPWR VPWR _6807_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1183 _3985_/X VGND VGND VPWR VPWR _6483_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1194 _4004_/X VGND VGND VPWR VPWR _6500_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_1_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_68_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4971_ _4971_/A _4971_/B VGND VGND VPWR VPWR _4971_/Y sky130_fd_sc_hd__nor2_1
XFILLER_64_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6710_ _7094_/CLK _6710_/D fanout494/X VGND VGND VPWR VPWR _6710_/Q sky130_fd_sc_hd__dfrtp_2
X_3922_ _3199_/Y input82/X _3958_/B VGND VGND VPWR VPWR _3922_/X sky130_fd_sc_hd__mux2_8
XFILLER_51_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3853_ _6453_/Q _3853_/B VGND VGND VPWR VPWR _3858_/B sky130_fd_sc_hd__nor2_1
X_6641_ _7193_/CLK _6641_/D VGND VGND VPWR VPWR _6641_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3784_ _7042_/Q hold77/A _4034_/A _6526_/Q _3783_/X VGND VGND VPWR VPWR _3788_/B
+ sky130_fd_sc_hd__a221o_1
X_6572_ _7108_/CLK _6572_/D fanout523/X VGND VGND VPWR VPWR _6572_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5523_ _5583_/A0 hold213/X _5528_/S VGND VGND VPWR VPWR _5523_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5454_ hold127/X hold291/X _5456_/S VGND VGND VPWR VPWR _5454_/X sky130_fd_sc_hd__mux2_1
X_4405_ _4560_/A _4731_/C _4731_/B VGND VGND VPWR VPWR _4758_/A sky130_fd_sc_hd__and3_4
X_5385_ _5385_/A _5385_/B VGND VGND VPWR VPWR _5393_/S sky130_fd_sc_hd__nand2_8
XFILLER_99_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7124_ _7126_/CLK _7124_/D fanout524/X VGND VGND VPWR VPWR _7124_/Q sky130_fd_sc_hd__dfrtp_1
X_4336_ _4390_/A _4390_/C _4390_/D VGND VGND VPWR VPWR _4547_/A sky130_fd_sc_hd__or3_4
XFILLER_59_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7055_ _7055_/CLK _7055_/D fanout522/X VGND VGND VPWR VPWR _7055_/Q sky130_fd_sc_hd__dfrtp_2
X_4267_ hold211/X _5583_/A0 _4269_/S VGND VGND VPWR VPWR _4267_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6006_ _6038_/A _6006_/B VGND VGND VPWR VPWR _6006_/Y sky130_fd_sc_hd__nor2_8
X_3218_ _6973_/Q VGND VGND VPWR VPWR _3218_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4198_ _4198_/A _5580_/B VGND VGND VPWR VPWR _4203_/S sky130_fd_sc_hd__and2_2
XFILLER_39_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_614 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6908_ _7123_/CLK _6908_/D fanout519/X VGND VGND VPWR VPWR _6908_/Q sky130_fd_sc_hd__dfrtp_4
X_6839_ _7053_/CLK _6839_/D fanout520/X VGND VGND VPWR VPWR _6839_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold280 _5425_/X VGND VGND VPWR VPWR _6997_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 _7023_/Q VGND VGND VPWR VPWR hold291/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_120 _3949_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_131 input84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_142 _3959_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_153 _6497_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_164 _6329_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_175 _3937_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_186 hold79/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_197 _3682_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5170_ _5170_/A _5170_/B _5170_/C _5169_/X VGND VGND VPWR VPWR _5171_/B sky130_fd_sc_hd__or4b_1
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4121_ _6393_/A0 hold977/X _4128_/S VGND VGND VPWR VPWR _4121_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4052_ _6407_/B _5232_/A VGND VGND VPWR VPWR _4052_/X sky130_fd_sc_hd__and2b_4
Xinput4 mask_rev_in[0] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4954_ _5158_/B _4954_/B _4954_/C _5158_/C VGND VGND VPWR VPWR _4960_/B sky130_fd_sc_hd__or4_1
X_3905_ _6014_/A _6000_/A VGND VGND VPWR VPWR _6018_/A sky130_fd_sc_hd__nand2_4
XFILLER_20_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4885_ _5039_/A _4885_/B _4885_/C _4885_/D VGND VGND VPWR VPWR _4885_/X sky130_fd_sc_hd__or4_1
XFILLER_20_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6624_ _6679_/CLK _6624_/D fanout511/X VGND VGND VPWR VPWR _6624_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_165_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3836_ hold72/A _6541_/Q _6545_/Q VGND VGND VPWR VPWR _3836_/Y sky130_fd_sc_hd__nor3_1
XFILLER_177_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3767_ _6766_/Q _4324_/A _4046_/A _6536_/Q VGND VGND VPWR VPWR _3767_/X sky130_fd_sc_hd__a22o_1
X_6555_ _6707_/CLK _6555_/D _6433_/A VGND VGND VPWR VPWR _6555_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5506_ _5584_/A0 hold476/X _5510_/S VGND VGND VPWR VPWR _5506_/X sky130_fd_sc_hd__mux2_1
X_6486_ _6760_/CLK _6486_/D fanout490/X VGND VGND VPWR VPWR _6486_/Q sky130_fd_sc_hd__dfrtp_1
X_3698_ _6499_/Q _3778_/A2 _5448_/A _7019_/Q _3697_/X VGND VGND VPWR VPWR _3701_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_106_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5437_ _5587_/A0 hold938/X _5438_/S VGND VGND VPWR VPWR _5437_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput330 hold1359/X VGND VGND VPWR VPWR hold1360/A sky130_fd_sc_hd__buf_12
XFILLER_133_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput341 hold1317/X VGND VGND VPWR VPWR hold1318/A sky130_fd_sc_hd__buf_12
X_5368_ _5581_/A0 _5368_/A1 _5375_/S VGND VGND VPWR VPWR _5368_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7107_ _7107_/CLK _7107_/D fanout511/X VGND VGND VPWR VPWR _7107_/Q sky130_fd_sc_hd__dfrtp_1
X_4319_ _4319_/A0 _6393_/A0 _4323_/S VGND VGND VPWR VPWR _4319_/X sky130_fd_sc_hd__mux2_1
X_5299_ _5584_/A0 hold465/X _5303_/S VGND VGND VPWR VPWR _5299_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7038_ _7050_/CLK _7038_/D fanout498/X VGND VGND VPWR VPWR _7038_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_28_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4670_ _4739_/A _4672_/A VGND VGND VPWR VPWR _4670_/Y sky130_fd_sc_hd__nor2_1
XFILLER_159_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3621_ _6688_/Q _4240_/A _4270_/A _6723_/Q _3615_/X VGND VGND VPWR VPWR _3621_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_174_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3552_ _7098_/Q _5535_/A _5221_/B _6814_/Q VGND VGND VPWR VPWR _3552_/X sky130_fd_sc_hd__a22o_1
X_6340_ _6674_/Q _6340_/A2 _6337_/X _6339_/X VGND VGND VPWR VPWR _6341_/D sky130_fd_sc_hd__a211o_1
XFILLER_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6271_ _6728_/Q _6320_/A2 _6320_/B1 _6618_/Q VGND VGND VPWR VPWR _6271_/X sky130_fd_sc_hd__a22o_2
XFILLER_142_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3483_ _7070_/Q _5502_/A _4022_/A _6520_/Q _3481_/X VGND VGND VPWR VPWR _3484_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5222_ _3714_/B _3538_/B _5536_/A1 hold967/X _5535_/B VGND VGND VPWR VPWR _5222_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_130_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5153_ _5153_/A _5153_/B _5152_/X VGND VGND VPWR VPWR _5153_/X sky130_fd_sc_hd__or3b_1
XFILLER_96_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4104_ _4104_/A _5580_/B VGND VGND VPWR VPWR _4110_/S sky130_fd_sc_hd__nand2_8
X_5084_ _5108_/A _5027_/B _5108_/B _4677_/B _4909_/Y VGND VGND VPWR VPWR _5153_/B
+ sky130_fd_sc_hd__o221ai_2
XFILLER_84_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_696 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4035_ _4035_/A0 _6393_/A0 _4039_/S VGND VGND VPWR VPWR _4035_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5986_ _7127_/Q _6320_/A2 _6320_/B1 _6874_/Q _5985_/X VGND VGND VPWR VPWR _6045_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_24_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4937_ _4462_/Y _4957_/B _4864_/D VGND VGND VPWR VPWR _5124_/C sky130_fd_sc_hd__a21o_1
XFILLER_33_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_20 _3410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_31 _3515_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4868_ _4868_/A _5068_/A _4868_/C _4868_/D VGND VGND VPWR VPWR _4868_/X sky130_fd_sc_hd__or4_1
XANTENNA_42 _3632_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_53 _5492_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_64 _5682_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6607_ _6725_/CLK _6607_/D fanout509/X VGND VGND VPWR VPWR _6607_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_75 _6045_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3819_ _3818_/Y _6468_/Q _3833_/S VGND VGND VPWR VPWR _6468_/D sky130_fd_sc_hd__mux2_1
X_4799_ _4996_/A _4802_/A _5076_/B _4659_/B VGND VGND VPWR VPWR _4799_/X sky130_fd_sc_hd__o22a_1
XANTENNA_86 _6708_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_97 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6538_ _6764_/CLK _6538_/D _3946_/B VGND VGND VPWR VPWR _6538_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_21_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6469_ _3927_/A1 _6469_/D _6424_/X VGND VGND VPWR VPWR hold46/A sky130_fd_sc_hd__dfrtp_1
XFILLER_161_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput171 _3959_/X VGND VGND VPWR VPWR debug_in sky130_fd_sc_hd__buf_12
XFILLER_133_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput182 _3218_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[16] sky130_fd_sc_hd__buf_12
Xoutput193 _3208_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[26] sky130_fd_sc_hd__buf_12
XFILLER_121_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_506 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5840_ _6929_/Q _5672_/X _5694_/X _7081_/Q _5839_/X VGND VGND VPWR VPWR _5847_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_34_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5771_ _5771_/A _5771_/B _5771_/C VGND VGND VPWR VPWR _5771_/X sky130_fd_sc_hd__or3_1
X_4722_ _5130_/A _4722_/B _4722_/C VGND VGND VPWR VPWR _4722_/X sky130_fd_sc_hd__or3_1
XFILLER_187_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4653_ _4814_/A _4832_/B _4653_/C VGND VGND VPWR VPWR _4653_/X sky130_fd_sc_hd__or3_1
Xinput40 mgmt_gpio_in[13] VGND VGND VPWR VPWR input40/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3604_ _7137_/Q hold69/A _5205_/A _6809_/Q VGND VGND VPWR VPWR _3604_/X sky130_fd_sc_hd__a22o_1
XFILLER_175_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput51 mgmt_gpio_in[23] VGND VGND VPWR VPWR input51/X sky130_fd_sc_hd__buf_2
Xhold802 _5257_/X VGND VGND VPWR VPWR _6848_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4584_ _4672_/A _5036_/A _4646_/A _4784_/B VGND VGND VPWR VPWR _4584_/X sky130_fd_sc_hd__o22a_1
Xinput62 mgmt_gpio_in[33] VGND VGND VPWR VPWR input62/X sky130_fd_sc_hd__clkbuf_2
Xinput73 pad_flash_io0_di VGND VGND VPWR VPWR _3952_/B sky130_fd_sc_hd__clkbuf_1
Xhold813 _6928_/Q VGND VGND VPWR VPWR hold813/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput84 spimemio_flash_csb VGND VGND VPWR VPWR input84/X sky130_fd_sc_hd__buf_2
Xhold824 _5266_/X VGND VGND VPWR VPWR _6856_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6323_ _7094_/Q _6323_/A2 _6323_/B1 _6740_/Q VGND VGND VPWR VPWR _6323_/X sky130_fd_sc_hd__a22o_1
XFILLER_155_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput95 usr1_vcc_pwrgood VGND VGND VPWR VPWR input95/X sky130_fd_sc_hd__buf_2
Xhold835 _5509_/X VGND VGND VPWR VPWR _7072_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3535_ _6942_/Q _5358_/A _4330_/A _6775_/Q VGND VGND VPWR VPWR _3535_/X sky130_fd_sc_hd__a22o_1
XFILLER_143_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold846 _6896_/Q VGND VGND VPWR VPWR hold846/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold857 _4213_/X VGND VGND VPWR VPWR _6667_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold868 _6836_/Q VGND VGND VPWR VPWR hold868/X sky130_fd_sc_hd__dlygate4sd3_1
X_6254_ _6772_/Q _6002_/Y _6007_/Y _6757_/Q _6253_/X VGND VGND VPWR VPWR _6257_/C
+ sky130_fd_sc_hd__a221o_1
X_3466_ hold21/X _3726_/B VGND VGND VPWR VPWR _4210_/A sky130_fd_sc_hd__nor2_4
XFILLER_130_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold879 _5564_/X VGND VGND VPWR VPWR _7120_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5205_ _5205_/A _5535_/B VGND VGND VPWR VPWR _5209_/S sky130_fd_sc_hd__and2_1
XFILLER_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3397_ _7117_/Q _3278_/Y _5268_/A _6864_/Q VGND VGND VPWR VPWR _3397_/X sky130_fd_sc_hd__a22o_1
X_6185_ _6856_/Q _6027_/A _6025_/A _6864_/Q _6184_/X VGND VGND VPWR VPWR _6192_/A
+ sky130_fd_sc_hd__a221o_1
Xhold1502 _5774_/X VGND VGND VPWR VPWR _7165_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1513 _6640_/Q VGND VGND VPWR VPWR _4182_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5136_ _5136_/A _5136_/B _4759_/Y VGND VGND VPWR VPWR _5137_/D sky130_fd_sc_hd__or3b_1
Xhold1524 _6654_/Q VGND VGND VPWR VPWR _4197_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1535 _7182_/Q VGND VGND VPWR VPWR _6220_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1546 _6639_/Q VGND VGND VPWR VPWR _4181_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1557 _6783_/Q VGND VGND VPWR VPWR _3792_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5067_ _5067_/A _5067_/B _5067_/C VGND VGND VPWR VPWR _5069_/A sky130_fd_sc_hd__nor3_1
Xhold1568 _6581_/Q VGND VGND VPWR VPWR hold237/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1579 _6580_/Q VGND VGND VPWR VPWR hold793/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4018_ _5531_/A1 hold946/X _4021_/S VGND VGND VPWR VPWR _4018_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_550 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5969_ _6563_/Q _7173_/Q _5968_/X VGND VGND VPWR VPWR _5969_/X sky130_fd_sc_hd__a21o_1
XFILLER_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold109 _5500_/X VGND VGND VPWR VPWR _7064_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3320_ _5212_/B _3334_/A VGND VGND VPWR VPWR _3320_/Y sky130_fd_sc_hd__nor2_8
XFILLER_98_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ _3971_/S hold17/X _3250_/Y VGND VGND VPWR VPWR hold18/A sky130_fd_sc_hd__o21ai_2
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6941_ _7138_/CLK _6941_/D fanout520/X VGND VGND VPWR VPWR _6941_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_81_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6872_ _6925_/CLK _6872_/D fanout516/X VGND VGND VPWR VPWR _6872_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5823_ _6968_/Q _5675_/X _5702_/X _6984_/Q VGND VGND VPWR VPWR _5823_/X sky130_fd_sc_hd__a22o_1
XFILLER_62_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5754_ _6901_/Q _5693_/X _5703_/X _6853_/Q VGND VGND VPWR VPWR _5754_/X sky130_fd_sc_hd__a22o_1
XFILLER_147_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4705_ _4814_/C _4707_/B _4703_/X _4704_/X VGND VGND VPWR VPWR _4705_/X sky130_fd_sc_hd__o211a_1
XFILLER_148_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5685_ _5938_/B _5705_/B _5699_/C VGND VGND VPWR VPWR _5685_/X sky130_fd_sc_hd__and3_4
XFILLER_8_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4636_ _5027_/A _5021_/B _4679_/B _5076_/B VGND VGND VPWR VPWR _4636_/X sky130_fd_sc_hd__o22a_1
XFILLER_175_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold610 _5472_/X VGND VGND VPWR VPWR _7039_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold621 _6847_/Q VGND VGND VPWR VPWR hold621/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4567_ _4846_/C _5023_/C VGND VGND VPWR VPWR _5016_/A sky130_fd_sc_hd__or2_4
Xhold632 _4293_/X VGND VGND VPWR VPWR _6740_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap351 _4083_/S VGND VGND VPWR VPWR _4085_/S sky130_fd_sc_hd__buf_8
Xhold643 _7070_/Q VGND VGND VPWR VPWR hold643/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6306_ _6714_/Q _6009_/X _6038_/Y _6724_/Q _6305_/X VGND VGND VPWR VPWR _6306_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_116_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold654 _5549_/X VGND VGND VPWR VPWR _7107_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold665 _6540_/Q VGND VGND VPWR VPWR hold665/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap373 _3320_/Y VGND VGND VPWR VPWR _5376_/A sky130_fd_sc_hd__buf_8
XFILLER_104_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3518_ hold57/X hold96/X VGND VGND VPWR VPWR _4276_/A sky130_fd_sc_hd__nor2_4
Xmax_cap384 _3476_/A VGND VGND VPWR VPWR _3507_/B sky130_fd_sc_hd__buf_12
Xhold676 _5363_/X VGND VGND VPWR VPWR _6942_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4498_ _4947_/A _4944_/B _4933_/A _4846_/B _4932_/A VGND VGND VPWR VPWR _4498_/X
+ sky130_fd_sc_hd__a2111o_1
Xmax_cap395 _6007_/Y VGND VGND VPWR VPWR _6025_/B sky130_fd_sc_hd__buf_8
Xhold687 _6710_/Q VGND VGND VPWR VPWR hold687/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold698 _4245_/X VGND VGND VPWR VPWR _6690_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6237_ _6686_/Q _5982_/X _6040_/X _6526_/Q VGND VGND VPWR VPWR _6237_/X sky130_fd_sc_hd__a22o_1
XFILLER_77_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3449_ _3448_/X _3449_/A1 _3917_/A VGND VGND VPWR VPWR _3449_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_588 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6168_ _6168_/A _6168_/B _6168_/C VGND VGND VPWR VPWR _6168_/X sky130_fd_sc_hd__or3_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1310 hold1310/A VGND VGND VPWR VPWR wb_dat_o[21] sky130_fd_sc_hd__buf_12
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1321 hold1407/X VGND VGND VPWR VPWR hold1321/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1332 hold1332/A VGND VGND VPWR VPWR wb_dat_o[7] sky130_fd_sc_hd__buf_12
Xhold1343 _4193_/A0 VGND VGND VPWR VPWR hold1343/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5119_ _5119_/A _5119_/B _5119_/C VGND VGND VPWR VPWR _5119_/Y sky130_fd_sc_hd__nor3_1
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1354 hold1354/A VGND VGND VPWR VPWR wb_dat_o[26] sky130_fd_sc_hd__buf_12
X_6099_ _7106_/Q _6025_/B _6272_/B _7069_/Q _6098_/X VGND VGND VPWR VPWR _6099_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_84_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1365 _6350_/A0 VGND VGND VPWR VPWR hold1365/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1376 _6830_/Q VGND VGND VPWR VPWR _5237_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1387 _6912_/Q VGND VGND VPWR VPWR _5329_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1398 _6631_/Q VGND VGND VPWR VPWR hold1398/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_3_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A VGND VGND VPWR VPWR _7181_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_53_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5470_ hold277/X hold36/X _5474_/S VGND VGND VPWR VPWR _5470_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4421_ _4605_/A _4436_/B VGND VGND VPWR VPWR _4758_/C sky130_fd_sc_hd__nor2_2
XFILLER_172_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7140_ _7140_/CLK _7140_/D fanout523/X VGND VGND VPWR VPWR _7140_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_172_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4352_ _4547_/A _4352_/B VGND VGND VPWR VPWR _4474_/A sky130_fd_sc_hd__or2_2
XFILLER_98_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3303_ _3303_/A _3378_/B VGND VGND VPWR VPWR _3528_/B sky130_fd_sc_hd__nand2_8
X_4283_ _6393_/A0 _4283_/A1 _4287_/S VGND VGND VPWR VPWR _4283_/X sky130_fd_sc_hd__mux2_1
X_7071_ _7071_/CLK _7071_/D fanout526/X VGND VGND VPWR VPWR _7071_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6022_ _6022_/A _6022_/B _6022_/C _6022_/D VGND VGND VPWR VPWR _6026_/A sky130_fd_sc_hd__or4_1
XFILLER_39_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6924_ _7136_/CLK _6924_/D fanout520/X VGND VGND VPWR VPWR _6924_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6855_ _7140_/CLK _6855_/D fanout522/X VGND VGND VPWR VPWR _6855_/Q sky130_fd_sc_hd__dfrtp_2
X_5806_ _6871_/Q _5683_/X _5706_/X _6503_/Q _5805_/X VGND VGND VPWR VPWR _5813_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_50_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6786_ _3487_/B2 _6786_/D _6437_/X VGND VGND VPWR VPWR _6786_/Q sky130_fd_sc_hd__dfrtn_1
X_3998_ _3998_/A0 hold127/X _4000_/S VGND VGND VPWR VPWR _3998_/X sky130_fd_sc_hd__mux2_1
X_5737_ _6868_/Q _5683_/X _5736_/X VGND VGND VPWR VPWR _5740_/C sky130_fd_sc_hd__a21o_1
XFILLER_13_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5668_ _6946_/Q _5666_/X _5667_/X _6874_/Q _5665_/X VGND VGND VPWR VPWR _5681_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_135_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4619_ _5016_/A _4659_/B VGND VGND VPWR VPWR _4986_/A sky130_fd_sc_hd__nor2_1
XFILLER_136_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5599_ _5606_/A _5599_/B _5599_/C VGND VGND VPWR VPWR _7144_/D sky130_fd_sc_hd__and3_1
XFILLER_151_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold440 _5524_/X VGND VGND VPWR VPWR _7085_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_151_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold451 _6829_/Q VGND VGND VPWR VPWR hold451/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 _4209_/X VGND VGND VPWR VPWR _6664_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold473 _4115_/X VGND VGND VPWR VPWR _6583_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 _6605_/Q VGND VGND VPWR VPWR hold484/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold495 _4208_/X VGND VGND VPWR VPWR _6663_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1140 _4149_/X VGND VGND VPWR VPWR _6612_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1151 _6602_/Q VGND VGND VPWR VPWR _4137_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1162 _4284_/X VGND VGND VPWR VPWR _6732_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1173 _6794_/Q VGND VGND VPWR VPWR _5189_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1184 hold1430/X VGND VGND VPWR VPWR _5467_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1195 hold1416/X VGND VGND VPWR VPWR _3994_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4970_ _4759_/A _4838_/B _5148_/A _5158_/A VGND VGND VPWR VPWR _5140_/A sky130_fd_sc_hd__a211o_1
XFILLER_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3921_ _3198_/Y input90/X _3921_/S VGND VGND VPWR VPWR _3921_/X sky130_fd_sc_hd__mux2_2
X_6640_ _7193_/CLK _6640_/D VGND VGND VPWR VPWR _6640_/Q sky130_fd_sc_hd__dfxtp_1
X_3852_ _3866_/S _3851_/Y _3856_/B VGND VGND VPWR VPWR _3853_/B sky130_fd_sc_hd__o21ba_1
XFILLER_149_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6571_ _7053_/CLK _6571_/D fanout518/X VGND VGND VPWR VPWR _6571_/Q sky130_fd_sc_hd__dfrtp_1
X_3783_ _6842_/Q _5250_/A _5225_/A _6823_/Q VGND VGND VPWR VPWR _3783_/X sky130_fd_sc_hd__a22o_1
XFILLER_192_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5522_ _5573_/A0 hold862/X _5528_/S VGND VGND VPWR VPWR _5522_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5453_ _5567_/A0 hold771/X _5456_/S VGND VGND VPWR VPWR _5453_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4404_ _4546_/A _4404_/B _4415_/A VGND VGND VPWR VPWR _4731_/B sky130_fd_sc_hd__nand3_2
XFILLER_99_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5384_ hold40/X hold183/X _5384_/S VGND VGND VPWR VPWR _5384_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7123_ _7123_/CLK _7123_/D fanout519/X VGND VGND VPWR VPWR _7123_/Q sky130_fd_sc_hd__dfrtp_1
X_4335_ _6397_/A0 hold530/X _4335_/S VGND VGND VPWR VPWR _4335_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7054_ _7139_/CLK _7054_/D fanout518/X VGND VGND VPWR VPWR _7054_/Q sky130_fd_sc_hd__dfrtp_4
X_4266_ hold405/X _5555_/A0 _4269_/S VGND VGND VPWR VPWR _4266_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_57_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7033_/CLK sky130_fd_sc_hd__clkbuf_16
X_6005_ _7026_/Q _6049_/B _6326_/A2 _6858_/Q _6004_/X VGND VGND VPWR VPWR _6012_/C
+ sky130_fd_sc_hd__a221o_1
X_3217_ _6981_/Q VGND VGND VPWR VPWR _3217_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4197_ _4197_/A0 _3373_/X _4197_/S VGND VGND VPWR VPWR _6654_/D sky130_fd_sc_hd__mux2_1
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6907_ _7123_/CLK _6907_/D _6407_/A VGND VGND VPWR VPWR _6907_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_23_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6838_ _6925_/CLK _6838_/D fanout516/X VGND VGND VPWR VPWR _6838_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6769_ _7050_/CLK _6769_/D fanout498/X VGND VGND VPWR VPWR _6769_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_109_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold270 _5419_/X VGND VGND VPWR VPWR _6992_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 _6576_/Q VGND VGND VPWR VPWR hold281/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 _5454_/X VGND VGND VPWR VPWR _7023_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_110 _3949_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_121 _3949_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_132 input84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_143 input35/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_154 _6292_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_165 _6329_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_176 _3927_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_187 hold85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_198 _3715_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4120_ hold96/X _4120_/B _6407_/B hold13/X VGND VGND VPWR VPWR _4128_/S sky130_fd_sc_hd__or4_4
XFILLER_69_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4051_ _6397_/A0 hold665/X _4051_/S VGND VGND VPWR VPWR _4051_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput5 mask_rev_in[10] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_615 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4953_ _4999_/B _4475_/A _4846_/D VGND VGND VPWR VPWR _5158_/C sky130_fd_sc_hd__o21a_1
X_3904_ _7156_/Q _7155_/Q VGND VGND VPWR VPWR _6000_/A sky130_fd_sc_hd__and2b_4
XFILLER_51_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4884_ _4931_/B _4870_/B _4971_/B _4744_/X VGND VGND VPWR VPWR _4885_/D sky130_fd_sc_hd__o31a_1
X_6623_ _6679_/CLK _6623_/D fanout511/X VGND VGND VPWR VPWR _6623_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_138_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3835_ _3914_/A1 _6462_/Q _3835_/S VGND VGND VPWR VPWR _6462_/D sky130_fd_sc_hd__mux2_1
XFILLER_192_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6554_ _6664_/CLK _6554_/D _6426_/A VGND VGND VPWR VPWR _6554_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3766_ _7095_/Q _5535_/A _4016_/A _6511_/Q _3736_/X VGND VGND VPWR VPWR _3789_/A
+ sky130_fd_sc_hd__a221o_1
X_5505_ _5583_/A0 hold249/X _5510_/S VGND VGND VPWR VPWR _5505_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6485_ _6760_/CLK _6485_/D fanout490/X VGND VGND VPWR VPWR _6485_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_146_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3697_ input15/X _3304_/Y _5225_/A _6822_/Q VGND VGND VPWR VPWR _3697_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5436_ _5550_/A0 hold677/X _5438_/S VGND VGND VPWR VPWR _5436_/X sky130_fd_sc_hd__mux2_1
Xoutput320 hold1341/X VGND VGND VPWR VPWR hold1342/A sky130_fd_sc_hd__buf_12
XFILLER_160_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput331 hold1309/X VGND VGND VPWR VPWR hold1310/A sky130_fd_sc_hd__buf_12
Xoutput342 hold1339/X VGND VGND VPWR VPWR hold1340/A sky130_fd_sc_hd__buf_12
X_5367_ _5367_/A _5571_/B VGND VGND VPWR VPWR _5375_/S sky130_fd_sc_hd__nand2_8
X_7106_ _7138_/CLK _7106_/D fanout525/X VGND VGND VPWR VPWR _7106_/Q sky130_fd_sc_hd__dfrtp_1
X_4318_ _4318_/A _6392_/B VGND VGND VPWR VPWR _4323_/S sky130_fd_sc_hd__and2_2
XFILLER_59_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5298_ _5574_/A0 _5298_/A1 _5303_/S VGND VGND VPWR VPWR _5298_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7037_ _7037_/CLK _7037_/D fanout515/X VGND VGND VPWR VPWR _7037_/Q sky130_fd_sc_hd__dfrtp_4
X_4249_ _4327_/A1 hold874/X _4251_/S VGND VGND VPWR VPWR _4249_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3620_ _6703_/Q _4246_/A _4198_/A _6657_/Q _3604_/X VGND VGND VPWR VPWR _3620_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_186_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3551_ _7037_/Q _5466_/A _4022_/A _6519_/Q VGND VGND VPWR VPWR _3551_/X sky130_fd_sc_hd__a22o_1
XFILLER_128_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6270_ _6270_/A1 _6319_/S _6268_/X _6269_/X VGND VGND VPWR VPWR _7184_/D sky130_fd_sc_hd__o22a_1
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3482_ _3507_/B _4120_/B VGND VGND VPWR VPWR _4022_/A sky130_fd_sc_hd__nor2_8
XFILLER_170_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5221_ _5221_/A _5221_/B VGND VGND VPWR VPWR _5221_/X sky130_fd_sc_hd__or2_1
XFILLER_88_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5152_ _4677_/B _5027_/B _5108_/B _4689_/B VGND VGND VPWR VPWR _5152_/X sky130_fd_sc_hd__o22a_1
XFILLER_57_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4103_ hold271/X _4102_/X _4103_/S VGND VGND VPWR VPWR _4103_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5083_ _5083_/A _5083_/B _5083_/C _5083_/D VGND VGND VPWR VPWR _5107_/B sky130_fd_sc_hd__or4_1
XFILLER_56_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4034_ _4034_/A _6392_/B VGND VGND VPWR VPWR _4039_/S sky130_fd_sc_hd__and2_2
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5985_ _6946_/Q _6024_/A _6308_/A2 _7135_/Q _5981_/X VGND VGND VPWR VPWR _5985_/X
+ sky130_fd_sc_hd__a221o_1
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4936_ _4947_/B VGND VGND VPWR VPWR _4957_/B sky130_fd_sc_hd__inv_2
XFILLER_33_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_10 _5466_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_21 _3410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4867_ _4684_/A _5060_/A _5126_/B _4847_/Y _4866_/X VGND VGND VPWR VPWR _4868_/D
+ sky130_fd_sc_hd__a2111o_1
XANTENNA_32 _3515_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_43 _3651_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_54 _5519_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6606_ _6679_/CLK _6606_/D fanout509/X VGND VGND VPWR VPWR _6606_/Q sky130_fd_sc_hd__dfrtp_4
X_3818_ _3818_/A _3818_/B VGND VGND VPWR VPWR _3818_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_192_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_65 _5683_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_76 _5998_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4798_ _4846_/B _4563_/B _4684_/B _4759_/B _4971_/A VGND VGND VPWR VPWR _4984_/C
+ sky130_fd_sc_hd__a32o_1
XANTENNA_87 _6989_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_98 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6537_ _6764_/CLK _6537_/D _3946_/B VGND VGND VPWR VPWR _6537_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_119_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3749_ _3749_/A _3749_/B _3749_/C _3749_/D VGND VGND VPWR VPWR _3790_/A sky130_fd_sc_hd__or4_2
XFILLER_134_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6468_ _3487_/B2 _6468_/D _6423_/X VGND VGND VPWR VPWR _6468_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5419_ _5569_/A0 hold269/X _5420_/S VGND VGND VPWR VPWR _5419_/X sky130_fd_sc_hd__mux2_1
X_6399_ _6426_/A _6441_/B VGND VGND VPWR VPWR _6399_/X sky130_fd_sc_hd__and2_1
Xoutput172 _6812_/Q VGND VGND VPWR VPWR irq[0] sky130_fd_sc_hd__buf_12
XFILLER_161_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput183 _3217_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[17] sky130_fd_sc_hd__buf_12
Xoutput194 _3207_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[27] sky130_fd_sc_hd__buf_12
XFILLER_153_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5770_ _5770_/A _5770_/B _5770_/C _5770_/D VGND VGND VPWR VPWR _5770_/X sky130_fd_sc_hd__or4_1
XFILLER_21_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4721_ _5018_/A _5021_/A _5016_/A VGND VGND VPWR VPWR _4992_/B sky130_fd_sc_hd__or3_2
X_4652_ _4832_/B _4653_/C VGND VGND VPWR VPWR _4652_/X sky130_fd_sc_hd__or2_1
XFILLER_30_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput30 mask_rev_in[4] VGND VGND VPWR VPWR input30/X sky130_fd_sc_hd__clkbuf_1
X_3603_ _3602_/X _3603_/A1 _3917_/A VGND VGND VPWR VPWR _3603_/X sky130_fd_sc_hd__mux2_1
Xinput41 mgmt_gpio_in[14] VGND VGND VPWR VPWR input41/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput52 mgmt_gpio_in[24] VGND VGND VPWR VPWR input52/X sky130_fd_sc_hd__clkbuf_1
X_4583_ _4814_/A _4814_/B VGND VGND VPWR VPWR _4784_/B sky130_fd_sc_hd__or2_4
XFILLER_116_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput63 mgmt_gpio_in[34] VGND VGND VPWR VPWR _3958_/A sky130_fd_sc_hd__clkbuf_8
Xhold803 _7075_/Q VGND VGND VPWR VPWR hold803/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput74 pad_flash_io1_di VGND VGND VPWR VPWR _3953_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold814 _5347_/X VGND VGND VPWR VPWR _6928_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6322_ _6755_/Q _6006_/Y _6322_/B1 _6750_/Q _6321_/X VGND VGND VPWR VPWR _6332_/B
+ sky130_fd_sc_hd__a221o_1
X_3534_ _3534_/A _3729_/B VGND VGND VPWR VPWR _4330_/A sky130_fd_sc_hd__nor2_4
Xhold825 _6888_/Q VGND VGND VPWR VPWR hold825/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput85 spimemio_flash_io0_do VGND VGND VPWR VPWR input85/X sky130_fd_sc_hd__buf_2
Xinput96 usr1_vdd_pwrgood VGND VGND VPWR VPWR input96/X sky130_fd_sc_hd__buf_2
Xhold836 _6968_/Q VGND VGND VPWR VPWR hold836/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold847 _5311_/X VGND VGND VPWR VPWR _6896_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold858 _7133_/Q VGND VGND VPWR VPWR hold858/X sky130_fd_sc_hd__dlygate4sd3_1
X_6253_ _6732_/Q _5997_/Y _6015_/X _6661_/Q VGND VGND VPWR VPWR _6253_/X sky130_fd_sc_hd__a22o_1
Xhold869 _5244_/X VGND VGND VPWR VPWR _6836_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3465_ hold57/X _3530_/B VGND VGND VPWR VPWR hold58/A sky130_fd_sc_hd__nor2_4
XFILLER_170_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5204_ _5536_/A1 _5204_/A1 _5204_/S VGND VGND VPWR VPWR _5204_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6184_ _6936_/Q _6024_/B _6024_/C _6912_/Q VGND VGND VPWR VPWR _6184_/X sky130_fd_sc_hd__a22o_1
X_3396_ _6936_/Q _5349_/A _5277_/A _6872_/Q _3395_/X VGND VGND VPWR VPWR _3409_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_97_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5135_ _4424_/Y _5036_/B _4758_/Y _4860_/A _4504_/B VGND VGND VPWR VPWR _5136_/B
+ sky130_fd_sc_hd__o2111ai_1
Xhold1503 _7204_/Q VGND VGND VPWR VPWR _6386_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1514 hold34/A VGND VGND VPWR VPWR _3864_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1525 hold61/A VGND VGND VPWR VPWR _6371_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1536 _6777_/Q VGND VGND VPWR VPWR _4929_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1547 _6641_/Q VGND VGND VPWR VPWR _4183_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1558 _7183_/Q VGND VGND VPWR VPWR _6245_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5066_ _5066_/A _5125_/A _5066_/C VGND VGND VPWR VPWR _5067_/C sky130_fd_sc_hd__or3_1
Xhold1569 _6445_/Q VGND VGND VPWR VPWR _3913_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_4017_ _5476_/A0 _4017_/A1 _4021_/S VGND VGND VPWR VPWR _4017_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5968_ _6600_/Q _5691_/Y _5957_/X _5967_/X _6318_/S VGND VGND VPWR VPWR _5968_/X
+ sky130_fd_sc_hd__o221a_2
X_4919_ _5021_/A _4639_/A _4665_/Y VGND VGND VPWR VPWR _4919_/X sky130_fd_sc_hd__o21ba_1
XFILLER_21_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5899_ _6661_/Q _5685_/X _5705_/X hold89/A VGND VGND VPWR VPWR _5899_/X sky130_fd_sc_hd__a22o_1
XFILLER_166_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ hold1531/X _3971_/S VGND VGND VPWR VPWR _3250_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_112_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6940_ _7136_/CLK _6940_/D fanout521/X VGND VGND VPWR VPWR _6940_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_19_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6871_ _7049_/CLK _6871_/D fanout522/X VGND VGND VPWR VPWR _6871_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5822_ _6504_/Q _5706_/X _5821_/X VGND VGND VPWR VPWR _5825_/C sky130_fd_sc_hd__a21o_1
XFILLER_50_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5753_ _5753_/A0 _5752_/X _6319_/S VGND VGND VPWR VPWR _5753_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4704_ _4814_/C _4704_/B VGND VGND VPWR VPWR _4704_/X sky130_fd_sc_hd__or2_1
XFILLER_148_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5684_ _7082_/Q _5682_/X _5683_/X _6866_/Q VGND VGND VPWR VPWR _5684_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4635_ _5027_/A _5021_/B VGND VGND VPWR VPWR _4635_/Y sky130_fd_sc_hd__nor2_1
XFILLER_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold600 _5517_/X VGND VGND VPWR VPWR _7079_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4566_ _4846_/B _4596_/B VGND VGND VPWR VPWR _5023_/C sky130_fd_sc_hd__or2_2
Xhold611 _7019_/Q VGND VGND VPWR VPWR hold611/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold622 _5256_/X VGND VGND VPWR VPWR _6847_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold633 _6910_/Q VGND VGND VPWR VPWR hold633/X sky130_fd_sc_hd__dlygate4sd3_1
X_6305_ _6704_/Q _6336_/A2 _6033_/X _7210_/Q VGND VGND VPWR VPWR _6305_/X sky130_fd_sc_hd__a22o_1
Xmax_cap352 _3335_/Y VGND VGND VPWR VPWR _5571_/A sky130_fd_sc_hd__buf_8
Xhold644 _5507_/X VGND VGND VPWR VPWR _7070_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap363 _6341_/A VGND VGND VPWR VPWR _6069_/A sky130_fd_sc_hd__clkbuf_2
X_3517_ _7139_/Q hold69/A _5349_/A _6934_/Q _3516_/X VGND VGND VPWR VPWR _3524_/A
+ sky130_fd_sc_hd__a221o_1
Xhold655 _7123_/Q VGND VGND VPWR VPWR hold655/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap374 _3298_/Y VGND VGND VPWR VPWR _5412_/A sky130_fd_sc_hd__buf_6
XFILLER_1_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold666 _4051_/X VGND VGND VPWR VPWR _6540_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4497_ _5076_/A _5013_/A VGND VGND VPWR VPWR _4882_/A sky130_fd_sc_hd__or2_1
Xmax_cap385 _3534_/A VGND VGND VPWR VPWR _3476_/A sky130_fd_sc_hd__buf_12
Xhold677 _7007_/Q VGND VGND VPWR VPWR hold677/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap396 _6006_/Y VGND VGND VPWR VPWR _6202_/B1 sky130_fd_sc_hd__buf_8
Xhold688 _4257_/X VGND VGND VPWR VPWR _6710_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6236_ _6670_/Q _6340_/A2 _6023_/D _6634_/Q _6235_/X VGND VGND VPWR VPWR _6242_/C
+ sky130_fd_sc_hd__a221o_1
Xhold699 hold699/A VGND VGND VPWR VPWR hold699/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_170_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3448_ _3447_/X _6787_/Q _3791_/A VGND VGND VPWR VPWR _3448_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6167_ _6167_/A _6167_/B _6167_/C _6167_/D VGND VGND VPWR VPWR _6168_/C sky130_fd_sc_hd__or4_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1300 _3984_/X VGND VGND VPWR VPWR _6482_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3379_ _3714_/B _3538_/B VGND VGND VPWR VPWR _5221_/B sky130_fd_sc_hd__nor2_8
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1311 hold1400/X VGND VGND VPWR VPWR hold1311/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1322 hold1322/A VGND VGND VPWR VPWR wb_dat_o[5] sky130_fd_sc_hd__buf_12
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5118_ _4538_/B _4478_/Y _4644_/B _4829_/Y _5117_/X VGND VGND VPWR VPWR _5119_/C
+ sky130_fd_sc_hd__a2111o_1
Xhold1333 hold1412/X VGND VGND VPWR VPWR hold1333/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1344 hold1344/A VGND VGND VPWR VPWR wb_dat_o[3] sky130_fd_sc_hd__buf_12
X_6098_ _6957_/Q _6336_/A2 _6323_/B1 _7122_/Q VGND VGND VPWR VPWR _6098_/X sky130_fd_sc_hd__a22o_1
Xhold1355 _4192_/A0 VGND VGND VPWR VPWR hold1355/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1366 hold1366/A VGND VGND VPWR VPWR wb_dat_o[25] sky130_fd_sc_hd__buf_12
Xhold1377 _5237_/X VGND VGND VPWR VPWR hold86/A sky130_fd_sc_hd__dlygate4sd3_1
X_5049_ _5049_/A _5049_/B _5049_/C _5049_/D VGND VGND VPWR VPWR _5151_/A sky130_fd_sc_hd__or4_1
XTAP_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1388 _6899_/Q VGND VGND VPWR VPWR _5315_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1399 _6677_/Q VGND VGND VPWR VPWR _4225_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4420_ _4420_/A _4570_/B _4846_/B VGND VGND VPWR VPWR _4738_/A sky130_fd_sc_hd__or3_4
XFILLER_132_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4351_ _4351_/A _4351_/B VGND VGND VPWR VPWR _4352_/B sky130_fd_sc_hd__nand2_1
XFILLER_125_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3302_ _3546_/B _3714_/B VGND VGND VPWR VPWR _5250_/A sky130_fd_sc_hd__nor2_8
X_7070_ _7070_/CLK _7070_/D fanout510/X VGND VGND VPWR VPWR _7070_/Q sky130_fd_sc_hd__dfrtp_4
X_4282_ _4282_/A _6392_/B VGND VGND VPWR VPWR _4287_/S sky130_fd_sc_hd__nand2_2
X_6021_ _6021_/A _6021_/B VGND VGND VPWR VPWR _6021_/Y sky130_fd_sc_hd__nor2_8
X_3233_ _6845_/Q VGND VGND VPWR VPWR _3233_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_1_1_1_csclk clkbuf_1_1_1_csclk/A VGND VGND VPWR VPWR clkbuf_2_3_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_104_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6923_ _6923_/CLK _6923_/D fanout514/X VGND VGND VPWR VPWR _6923_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_35_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6854_ _6990_/CLK _6854_/D _3873_/A VGND VGND VPWR VPWR _6854_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_22_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5805_ _7023_/Q _5663_/X _5666_/X _6951_/Q VGND VGND VPWR VPWR _5805_/X sky130_fd_sc_hd__a22o_1
X_6785_ _3945_/A1 _6785_/D _6436_/X VGND VGND VPWR VPWR _6785_/Q sky130_fd_sc_hd__dfrtn_1
X_3997_ hold516/X _6397_/A0 _4000_/S VGND VGND VPWR VPWR _3997_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5736_ _6932_/Q _5670_/X _5685_/X _6908_/Q VGND VGND VPWR VPWR _5736_/X sky130_fd_sc_hd__a22o_1
XFILLER_182_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5667_ _5938_/B _5705_/B _5700_/C VGND VGND VPWR VPWR _5667_/X sky130_fd_sc_hd__and3_4
XFILLER_136_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4618_ _5107_/A _4916_/A _4618_/C _4618_/D VGND VGND VPWR VPWR _4642_/A sky130_fd_sc_hd__and4b_1
XFILLER_190_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5598_ _7144_/Q _5604_/D VGND VGND VPWR VPWR _5599_/C sky130_fd_sc_hd__or2_1
XFILLER_190_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold430 _5443_/X VGND VGND VPWR VPWR _7013_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4549_ _4963_/A VGND VGND VPWR VPWR _4549_/Y sky130_fd_sc_hd__inv_2
Xhold441 hold441/A VGND VGND VPWR VPWR hold441/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold452 _5236_/X VGND VGND VPWR VPWR _6829_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 _6600_/Q VGND VGND VPWR VPWR hold463/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold474 _7211_/Q VGND VGND VPWR VPWR hold474/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold485 _4140_/X VGND VGND VPWR VPWR _6605_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold496 _6529_/Q VGND VGND VPWR VPWR hold496/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6219_ _7181_/Q _6218_/X _6318_/S VGND VGND VPWR VPWR _6219_/X sky130_fd_sc_hd__mux2_1
XFILLER_104_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7199_ _7200_/CLK _7199_/D fanout529/X VGND VGND VPWR VPWR hold61/A sky130_fd_sc_hd__dfrtp_1
XFILLER_58_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1130 _4138_/X VGND VGND VPWR VPWR _6603_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1141 _6517_/Q VGND VGND VPWR VPWR _4024_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1152 _4137_/X VGND VGND VPWR VPWR _6602_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1163 _6800_/Q VGND VGND VPWR VPWR _5196_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_161_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1174 _5189_/X VGND VGND VPWR VPWR _6794_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1185 _6475_/Q VGND VGND VPWR VPWR _3970_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1196 _6763_/Q VGND VGND VPWR VPWR _4321_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_721 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3920_ _3197_/Y input92/X _3921_/S VGND VGND VPWR VPWR _3920_/X sky130_fd_sc_hd__mux2_2
XFILLER_17_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3851_ _6455_/Q _6454_/Q _3834_/B VGND VGND VPWR VPWR _3851_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_177_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6570_ _6925_/CLK _6570_/D fanout516/X VGND VGND VPWR VPWR _6570_/Q sky130_fd_sc_hd__dfrtp_1
X_3782_ _6474_/Q _3966_/A _5184_/A _6791_/Q _3735_/X VGND VGND VPWR VPWR _3788_/A
+ sky130_fd_sc_hd__a221o_1
X_5521_ _5521_/A0 _5521_/A1 _5528_/S VGND VGND VPWR VPWR _5521_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5452_ _5584_/A0 hold427/X _5456_/S VGND VGND VPWR VPWR _5452_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4403_ _4404_/B _4415_/A _4546_/A VGND VGND VPWR VPWR _4731_/C sky130_fd_sc_hd__a21o_1
X_5383_ _5587_/A0 hold884/X _5384_/S VGND VGND VPWR VPWR _5383_/X sky130_fd_sc_hd__mux2_1
X_7122_ _7138_/CLK _7122_/D fanout521/X VGND VGND VPWR VPWR _7122_/Q sky130_fd_sc_hd__dfrtp_4
X_4334_ _6396_/A0 hold459/X _4335_/S VGND VGND VPWR VPWR _4334_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7053_ _7053_/CLK _7053_/D fanout520/X VGND VGND VPWR VPWR _7053_/Q sky130_fd_sc_hd__dfrtp_4
X_4265_ _4265_/A0 _5212_/C _4269_/S VGND VGND VPWR VPWR _4265_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6004_ _7018_/Q _6002_/Y _6340_/A2 _6922_/Q VGND VGND VPWR VPWR _6004_/X sky130_fd_sc_hd__a22o_1
XFILLER_101_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3216_ _6989_/Q VGND VGND VPWR VPWR _3216_/Y sky130_fd_sc_hd__inv_2
X_4196_ _4196_/A0 _3410_/X _4197_/S VGND VGND VPWR VPWR _6653_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6906_ _7123_/CLK _6906_/D _6407_/A VGND VGND VPWR VPWR _6906_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_23_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6837_ _6925_/CLK _6837_/D fanout516/X VGND VGND VPWR VPWR _6837_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_10_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6768_ _6825_/CLK _6768_/D fanout490/X VGND VGND VPWR VPWR _6768_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_10_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5719_ _5719_/A _5719_/B _5719_/C _5719_/D VGND VGND VPWR VPWR _5719_/X sky130_fd_sc_hd__or4_1
XFILLER_148_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6699_ _7200_/CLK _6699_/D _6348_/B VGND VGND VPWR VPWR _6699_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_148_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold260 _5540_/X VGND VGND VPWR VPWR _7099_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 _6573_/Q VGND VGND VPWR VPWR hold271/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 _4107_/X VGND VGND VPWR VPWR _6576_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 _6712_/Q VGND VGND VPWR VPWR hold293/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_93_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_100 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_111 _3949_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_122 _3949_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_133 input84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_144 _4951_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_155 _6044_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_166 _6024_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_177 _3927_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_188 _5203_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_199 _3717_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_731 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4050_ _5533_/A1 hold761/X _4051_/S VGND VGND VPWR VPWR _4050_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput6 mask_rev_in[11] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4952_ _4952_/A _5031_/B _5059_/B VGND VGND VPWR VPWR _4954_/C sky130_fd_sc_hd__or3_1
X_3903_ _7153_/Q _7154_/Q VGND VGND VPWR VPWR _6014_/A sky130_fd_sc_hd__and2b_4
X_4883_ _4931_/B _4657_/C _4870_/B _4876_/A VGND VGND VPWR VPWR _4885_/C sky130_fd_sc_hd__o31a_1
XFILLER_177_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3834_ _6541_/Q _3834_/B VGND VGND VPWR VPWR _3835_/S sky130_fd_sc_hd__nand2_1
X_6622_ _6679_/CLK _6622_/D fanout511/X VGND VGND VPWR VPWR _6622_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_177_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6553_ _7136_/CLK _6553_/D fanout520/X VGND VGND VPWR VPWR _6553_/Q sky130_fd_sc_hd__dfrtp_1
X_3765_ _6611_/Q _4147_/A _3760_/X _3764_/X _3472_/Y VGND VGND VPWR VPWR _3790_/C
+ sky130_fd_sc_hd__a2111o_1
XFILLER_158_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5504_ _5573_/A0 hold651/X _5510_/S VGND VGND VPWR VPWR _5504_/X sky130_fd_sc_hd__mux2_1
X_6484_ _6760_/CLK _6484_/D fanout490/X VGND VGND VPWR VPWR _6484_/Q sky130_fd_sc_hd__dfstp_2
X_3696_ input44/X _3308_/Y _4102_/S input72/X _3695_/X VGND VGND VPWR VPWR _3701_/B
+ sky130_fd_sc_hd__a221o_1
X_5435_ _5549_/A0 hold649/X _5438_/S VGND VGND VPWR VPWR _5435_/X sky130_fd_sc_hd__mux2_1
Xoutput310 _3940_/X VGND VGND VPWR VPWR serial_load sky130_fd_sc_hd__buf_12
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput321 hold1327/X VGND VGND VPWR VPWR hold1328/A sky130_fd_sc_hd__buf_12
XFILLER_133_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput332 hold1305/X VGND VGND VPWR VPWR hold1306/A sky130_fd_sc_hd__buf_12
XFILLER_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput343 hold1343/X VGND VGND VPWR VPWR hold1344/A sky130_fd_sc_hd__buf_12
X_5366_ _5579_/A0 hold508/X _5366_/S VGND VGND VPWR VPWR _5366_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4317_ hold488/X _6397_/A0 _4317_/S VGND VGND VPWR VPWR _4317_/X sky130_fd_sc_hd__mux2_1
X_7105_ _7129_/CLK _7105_/D fanout518/X VGND VGND VPWR VPWR _7105_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_59_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5297_ _5555_/A0 hold351/X _5303_/S VGND VGND VPWR VPWR _5297_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7036_ _7137_/CLK _7036_/D fanout501/X VGND VGND VPWR VPWR _7036_/Q sky130_fd_sc_hd__dfrtp_4
X_4248_ _5531_/A1 hold930/X _4251_/S VGND VGND VPWR VPWR _4248_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_48 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4179_ _5534_/A1 hold361/X _4179_/S VGND VGND VPWR VPWR _4179_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_41_csclk _6931_/CLK VGND VGND VPWR VPWR _6992_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_56_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7141_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_186_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3550_ _7069_/Q _5502_/A hold77/A _7045_/Q VGND VGND VPWR VPWR _3550_/X sky130_fd_sc_hd__a22o_2
XFILLER_155_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3481_ _6478_/Q _3966_/A _3992_/A _6494_/Q VGND VGND VPWR VPWR _3481_/X sky130_fd_sc_hd__a22o_2
X_5220_ _5555_/A0 hold355/X _5220_/S VGND VGND VPWR VPWR _5220_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5151_ _5151_/A _5151_/B _5151_/C _5174_/C VGND VGND VPWR VPWR _5151_/X sky130_fd_sc_hd__or4_1
XFILLER_96_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4102_ hold81/X hold40/X _4102_/S VGND VGND VPWR VPWR _4102_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5082_ _4694_/B _5108_/B _5015_/B VGND VGND VPWR VPWR _5083_/D sky130_fd_sc_hd__o21bai_1
XFILLER_96_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4033_ hold721/X _5534_/A1 _4033_/S VGND VGND VPWR VPWR _4033_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5984_ _6019_/A _6021_/B VGND VGND VPWR VPWR _6023_/B sky130_fd_sc_hd__nor2_4
XFILLER_52_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4935_ _4935_/A _4935_/B _4935_/C VGND VGND VPWR VPWR _4947_/B sky130_fd_sc_hd__or3_1
Xclkbuf_3_7_0_csclk clkbuf_3_7_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_7_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_11 _5340_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_22 _3410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4866_ _5126_/A _5162_/A _4866_/C _4866_/D VGND VGND VPWR VPWR _4866_/X sky130_fd_sc_hd__or4_1
XANTENNA_33 _3542_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6605_ _7209_/CLK _6605_/D fanout485/X VGND VGND VPWR VPWR _6605_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA_44 _3721_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_55 _5659_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3817_ hold72/A _3821_/S _6467_/Q VGND VGND VPWR VPWR _3818_/B sky130_fd_sc_hd__o21a_1
XFILLER_165_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_66 _5683_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4797_ _4797_/A _4797_/B VGND VGND VPWR VPWR _4810_/D sky130_fd_sc_hd__nand2_1
XFILLER_165_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_77 _6007_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_88 _7061_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6536_ _6764_/CLK _6536_/D _3946_/B VGND VGND VPWR VPWR _6536_/Q sky130_fd_sc_hd__dfrtp_2
X_3748_ _7111_/Q _5553_/A _4174_/A _6634_/Q _3747_/X VGND VGND VPWR VPWR _3749_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA_99 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3679_ _3679_/A _3679_/B _3679_/C _3679_/D VGND VGND VPWR VPWR _3689_/A sky130_fd_sc_hd__or4_1
X_6467_ _3487_/B2 _6467_/D _6422_/X VGND VGND VPWR VPWR _6467_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5418_ _5550_/A0 hold613/X _5420_/S VGND VGND VPWR VPWR _5418_/X sky130_fd_sc_hd__mux2_1
X_6398_ _6433_/A _6440_/B VGND VGND VPWR VPWR _6398_/X sky130_fd_sc_hd__and2_1
XFILLER_0_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput173 _3960_/X VGND VGND VPWR VPWR irq[1] sky130_fd_sc_hd__buf_12
XFILLER_0_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5349_ _5349_/A _5385_/B VGND VGND VPWR VPWR _5357_/S sky130_fd_sc_hd__nand2_8
Xoutput184 _3216_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[18] sky130_fd_sc_hd__buf_12
Xoutput195 _3206_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[28] sky130_fd_sc_hd__buf_12
XFILLER_102_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7019_ _7136_/CLK _7019_/D fanout519/X VGND VGND VPWR VPWR _7019_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4720_ _5031_/B _4899_/B _4720_/C VGND VGND VPWR VPWR _4722_/C sky130_fd_sc_hd__or3_1
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4651_ _4693_/A _5023_/B VGND VGND VPWR VPWR _4707_/B sky130_fd_sc_hd__or2_4
XFILLER_174_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput20 mask_rev_in[24] VGND VGND VPWR VPWR input20/X sky130_fd_sc_hd__clkbuf_1
X_3602_ _3601_/X _6785_/Q _3791_/A VGND VGND VPWR VPWR _3602_/X sky130_fd_sc_hd__mux2_1
Xinput31 mask_rev_in[5] VGND VGND VPWR VPWR input31/X sky130_fd_sc_hd__clkbuf_1
X_4582_ _5016_/A _4582_/B VGND VGND VPWR VPWR _4984_/A sky130_fd_sc_hd__nor2_1
Xinput42 mgmt_gpio_in[15] VGND VGND VPWR VPWR input42/X sky130_fd_sc_hd__clkbuf_4
XFILLER_174_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput53 mgmt_gpio_in[25] VGND VGND VPWR VPWR input53/X sky130_fd_sc_hd__clkbuf_2
Xinput64 mgmt_gpio_in[35] VGND VGND VPWR VPWR input64/X sky130_fd_sc_hd__clkbuf_2
Xinput75 porb VGND VGND VPWR VPWR input75/X sky130_fd_sc_hd__clkbuf_1
X_6321_ _6775_/Q _6002_/Y _6030_/X _6745_/Q VGND VGND VPWR VPWR _6321_/X sky130_fd_sc_hd__a22o_1
X_3533_ _7006_/Q _5430_/A _5544_/A _7107_/Q _3532_/X VGND VGND VPWR VPWR _3541_/B
+ sky130_fd_sc_hd__a221o_1
Xhold804 _5513_/X VGND VGND VPWR VPWR _7075_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold815 _6964_/Q VGND VGND VPWR VPWR hold815/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput86 spimemio_flash_io0_oeb VGND VGND VPWR VPWR _3947_/B sky130_fd_sc_hd__clkbuf_4
Xhold826 _5302_/X VGND VGND VPWR VPWR _6888_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold837 _5392_/X VGND VGND VPWR VPWR _6968_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput97 usr2_vcc_pwrgood VGND VGND VPWR VPWR input97/X sky130_fd_sc_hd__buf_2
XFILLER_116_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold848 _6971_/Q VGND VGND VPWR VPWR hold848/X sky130_fd_sc_hd__dlygate4sd3_1
X_6252_ _6507_/Q _6049_/B _6006_/Y _6752_/Q _6248_/X VGND VGND VPWR VPWR _6257_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold859 _5578_/X VGND VGND VPWR VPWR _7133_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3464_ _6755_/Q _4306_/A _4294_/A _6745_/Q VGND VGND VPWR VPWR _3464_/X sky130_fd_sc_hd__a22o_1
X_5203_ _5203_/A _5203_/B VGND VGND VPWR VPWR _5204_/S sky130_fd_sc_hd__nand2_1
X_6183_ _7133_/Q _6023_/A _6022_/A _6880_/Q _6182_/X VGND VGND VPWR VPWR _6193_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3395_ _6968_/Q _5385_/A _3393_/X _3394_/X VGND VGND VPWR VPWR _3395_/X sky130_fd_sc_hd__a211o_1
XFILLER_97_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5134_ _5134_/A _5134_/B _5134_/C _5134_/D VGND VGND VPWR VPWR _5148_/D sky130_fd_sc_hd__or4_1
Xhold1504 _7164_/Q VGND VGND VPWR VPWR _5753_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1515 _6824_/Q VGND VGND VPWR VPWR hold1515/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1526 _7198_/Q VGND VGND VPWR VPWR hold7/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1537 _7174_/Q VGND VGND VPWR VPWR _5970_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5065_ _5065_/A _5065_/B _5065_/C _5065_/D VGND VGND VPWR VPWR _5066_/C sky130_fd_sc_hd__or4_1
XFILLER_123_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1548 _7188_/Q VGND VGND VPWR VPWR _6347_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1559 _6454_/Q VGND VGND VPWR VPWR _3855_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4016_ _4016_/A _4330_/B VGND VGND VPWR VPWR _4021_/S sky130_fd_sc_hd__nand2_2
XFILLER_38_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5967_ _5967_/A _5967_/B _5967_/C _5967_/D VGND VGND VPWR VPWR _5967_/X sky130_fd_sc_hd__or4_1
X_4918_ _5023_/A _5016_/A _4719_/A VGND VGND VPWR VPWR _4963_/B sky130_fd_sc_hd__a21oi_2
XFILLER_33_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5898_ _6635_/Q _5655_/X _5688_/X _6607_/Q _5897_/X VGND VGND VPWR VPWR _5901_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4849_ _5002_/A _5035_/B _4708_/A VGND VGND VPWR VPWR _4865_/C sky130_fd_sc_hd__o21ai_1
XFILLER_193_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6519_ _6708_/CLK _6519_/D _6432_/A VGND VGND VPWR VPWR _6519_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_107_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6870_ _7082_/CLK _6870_/D _3873_/A VGND VGND VPWR VPWR _6870_/Q sky130_fd_sc_hd__dfrtp_4
X_5821_ _7008_/Q _5664_/X _5686_/X _7016_/Q VGND VGND VPWR VPWR _5821_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5752_ _5650_/A _7163_/Q _5751_/X VGND VGND VPWR VPWR _5752_/X sky130_fd_sc_hd__a21o_1
X_4703_ _4639_/B _4704_/B _4701_/X _4702_/X VGND VGND VPWR VPWR _4703_/X sky130_fd_sc_hd__o211a_1
XFILLER_175_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5683_ _5938_/B _5706_/B _5703_/B VGND VGND VPWR VPWR _5683_/X sky130_fd_sc_hd__and3_4
XFILLER_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4634_ _4634_/A _4915_/A _4987_/A _4982_/A VGND VGND VPWR VPWR _4642_/B sky130_fd_sc_hd__nor4_1
XFILLER_163_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold601 _6969_/Q VGND VGND VPWR VPWR hold601/X sky130_fd_sc_hd__dlygate4sd3_1
X_4565_ _4621_/B _4666_/B VGND VGND VPWR VPWR _4784_/A sky130_fd_sc_hd__or2_4
Xhold612 _5450_/X VGND VGND VPWR VPWR _7019_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold623 _7030_/Q VGND VGND VPWR VPWR hold623/X sky130_fd_sc_hd__dlygate4sd3_1
X_6304_ _6774_/Q _6002_/Y _6007_/Y _6759_/Q _6303_/X VGND VGND VPWR VPWR _6304_/X
+ sky130_fd_sc_hd__a221o_1
Xhold634 _5327_/X VGND VGND VPWR VPWR _6910_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3516_ _6958_/Q _5376_/A _5385_/A _6966_/Q VGND VGND VPWR VPWR _3516_/X sky130_fd_sc_hd__a22o_1
Xhold645 _6901_/Q VGND VGND VPWR VPWR hold645/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap353 _3333_/Y VGND VGND VPWR VPWR _3751_/A2 sky130_fd_sc_hd__buf_8
Xmax_cap364 _6094_/A VGND VGND VPWR VPWR _6341_/A sky130_fd_sc_hd__clkbuf_2
X_4496_ _4745_/A _5094_/A VGND VGND VPWR VPWR _5050_/A sky130_fd_sc_hd__or2_1
Xhold656 _5567_/X VGND VGND VPWR VPWR _7123_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap375 _4001_/A VGND VGND VPWR VPWR _3778_/A2 sky130_fd_sc_hd__buf_12
Xhold667 _6869_/Q VGND VGND VPWR VPWR hold667/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap386 _3300_/A VGND VGND VPWR VPWR _3534_/A sky130_fd_sc_hd__buf_12
Xhold678 _5436_/X VGND VGND VPWR VPWR _7007_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6235_ _6665_/Q wire412/X _6016_/X _6681_/Q VGND VGND VPWR VPWR _6235_/X sky130_fd_sc_hd__a22o_1
Xmax_cap397 _6002_/Y VGND VGND VPWR VPWR _6204_/A2 sky130_fd_sc_hd__buf_8
XFILLER_89_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold689 _6673_/Q VGND VGND VPWR VPWR hold689/X sky130_fd_sc_hd__dlygate4sd3_1
X_3447_ _3447_/A _3447_/B _3447_/C _3447_/D VGND VGND VPWR VPWR _3447_/X sky130_fd_sc_hd__or4_4
XFILLER_103_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3378_ hold75/X _3378_/B VGND VGND VPWR VPWR _3538_/B sky130_fd_sc_hd__nand2_8
XFILLER_134_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6166_ _6871_/Q _6199_/B1 _6025_/D _6967_/Q _6165_/X VGND VGND VPWR VPWR _6167_/D
+ sky130_fd_sc_hd__a221o_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1301 _6761_/Q VGND VGND VPWR VPWR _4319_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1312 hold1312/A VGND VGND VPWR VPWR wb_dat_o[14] sky130_fd_sc_hd__buf_12
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1323 hold1406/X VGND VGND VPWR VPWR hold1323/X sky130_fd_sc_hd__dlygate4sd3_1
X_5117_ _4971_/A _4783_/Y _4973_/B VGND VGND VPWR VPWR _5117_/X sky130_fd_sc_hd__a21o_1
X_6097_ _6121_/A2 _6096_/X _6319_/S VGND VGND VPWR VPWR _6097_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1334 hold1334/A VGND VGND VPWR VPWR wb_dat_o[9] sky130_fd_sc_hd__buf_12
XFILLER_111_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1345 _4190_/A0 VGND VGND VPWR VPWR hold1345/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1356 hold1356/A VGND VGND VPWR VPWR wb_dat_o[2] sky130_fd_sc_hd__buf_12
Xhold1367 _6349_/A0 VGND VGND VPWR VPWR hold1367/X sky130_fd_sc_hd__dlygate4sd3_1
X_5048_ _5134_/C _5132_/A _5048_/C VGND VGND VPWR VPWR _5048_/X sky130_fd_sc_hd__or3_1
Xhold1378 _6832_/Q VGND VGND VPWR VPWR _5239_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1389 _6875_/Q VGND VGND VPWR VPWR _5288_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6999_ _7110_/CLK _6999_/D fanout507/X VGND VGND VPWR VPWR _6999_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_159_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4350_ _4654_/A _4350_/B _4542_/A VGND VGND VPWR VPWR _4351_/B sky130_fd_sc_hd__nand3_1
XFILLER_125_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3301_ hold48/X hold18/X _3301_/C VGND VGND VPWR VPWR _3547_/B sky130_fd_sc_hd__or3_4
XFILLER_98_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4281_ _5567_/A0 hold629/X _4281_/S VGND VGND VPWR VPWR _4281_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6020_ _6033_/A _6039_/A _6020_/C VGND VGND VPWR VPWR _6020_/X sky130_fd_sc_hd__and3_4
X_3232_ _6853_/Q VGND VGND VPWR VPWR _3232_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6922_ _7012_/CLK _6922_/D fanout505/X VGND VGND VPWR VPWR _6922_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_82_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6853_ _7053_/CLK _6853_/D fanout518/X VGND VGND VPWR VPWR _6853_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_50_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5804_ _6999_/Q _5656_/X _5799_/X _5803_/X VGND VGND VPWR VPWR _5804_/X sky130_fd_sc_hd__a211o_1
X_6784_ _3927_/A1 _6784_/D _6435_/X VGND VGND VPWR VPWR _6784_/Q sky130_fd_sc_hd__dfrtn_1
X_3996_ hold526/X _6396_/A0 _4000_/S VGND VGND VPWR VPWR _3996_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5735_ _6884_/Q _5846_/A2 _5666_/X _6948_/Q _5734_/X VGND VGND VPWR VPWR _5740_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5666_ _5938_/B _5706_/C _5703_/C VGND VGND VPWR VPWR _5666_/X sky130_fd_sc_hd__and3_4
XFILLER_108_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4617_ _4420_/A _4667_/C _4846_/B _4684_/B _5019_/A VGND VGND VPWR VPWR _5107_/A
+ sky130_fd_sc_hd__a41o_1
XFILLER_163_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5597_ _7144_/Q _5604_/D VGND VGND VPWR VPWR _5599_/B sky130_fd_sc_hd__nand2_1
Xhold420 _5526_/X VGND VGND VPWR VPWR _7087_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold431 _6557_/Q VGND VGND VPWR VPWR hold431/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_163_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4548_ _4780_/A _4802_/B _6699_/Q VGND VGND VPWR VPWR _4963_/A sky130_fd_sc_hd__o21ai_2
XFILLER_89_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold442 _5247_/X VGND VGND VPWR VPWR _6839_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold453 _6770_/Q VGND VGND VPWR VPWR hold453/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold464 _4134_/X VGND VGND VPWR VPWR _6600_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 _6397_/X VGND VGND VPWR VPWR _7211_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 _6486_/Q VGND VGND VPWR VPWR hold486/X sky130_fd_sc_hd__dlygate4sd3_1
X_4479_ _5076_/A _4672_/A VGND VGND VPWR VPWR _5148_/A sky130_fd_sc_hd__nor2_4
Xhold497 _4038_/X VGND VGND VPWR VPWR _6529_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6218_ _6201_/X _6207_/X _6217_/X _6046_/B _6849_/Q VGND VGND VPWR VPWR _6218_/X
+ sky130_fd_sc_hd__o32a_1
X_7198_ _7200_/CLK _7198_/D _6348_/B VGND VGND VPWR VPWR _7198_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1120 _5574_/X VGND VGND VPWR VPWR _7129_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6149_ _7087_/Q _5977_/X _6323_/B1 _7124_/Q VGND VGND VPWR VPWR _6149_/X sky130_fd_sc_hd__a22o_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1131 _7004_/Q VGND VGND VPWR VPWR _5433_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1142 _4024_/X VGND VGND VPWR VPWR _6517_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1153 _7052_/Q VGND VGND VPWR VPWR _5487_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1164 _5196_/X VGND VGND VPWR VPWR _6800_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1175 hold1456/X VGND VGND VPWR VPWR _3995_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1186 _3970_/X VGND VGND VPWR VPWR _6475_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1197 _6575_/Q VGND VGND VPWR VPWR _4106_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_733 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3850_ hold72/A _3850_/B _6541_/Q VGND VGND VPWR VPWR _3866_/S sky130_fd_sc_hd__or3_4
X_3781_ _3781_/A _3781_/B _3781_/C _3781_/D VGND VGND VPWR VPWR _3789_/C sky130_fd_sc_hd__or4_1
X_5520_ _5520_/A _5571_/B VGND VGND VPWR VPWR _5528_/S sky130_fd_sc_hd__nand2_8
XFILLER_157_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5451_ _5583_/A0 hold287/X _5456_/S VGND VGND VPWR VPWR _5451_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4402_ _4935_/A _4819_/C _4538_/B VGND VGND VPWR VPWR _4415_/A sky130_fd_sc_hd__and3_1
X_5382_ _5586_/A0 _5382_/A1 _5384_/S VGND VGND VPWR VPWR _5382_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7121_ _7136_/CLK _7121_/D fanout520/X VGND VGND VPWR VPWR _7121_/Q sky130_fd_sc_hd__dfrtp_1
X_4333_ _6395_/A0 _4333_/A1 _4335_/S VGND VGND VPWR VPWR _4333_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4264_ _4264_/A _5535_/B VGND VGND VPWR VPWR _4269_/S sky130_fd_sc_hd__and2_2
XFILLER_101_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7052_ _7053_/CLK _7052_/D fanout526/X VGND VGND VPWR VPWR _7052_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_115_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6003_ _6014_/A _6020_/C _6040_/C VGND VGND VPWR VPWR _6027_/B sky130_fd_sc_hd__and3_4
X_3215_ _6997_/Q VGND VGND VPWR VPWR _3215_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4195_ _4195_/A0 _3447_/X _4197_/S VGND VGND VPWR VPWR _6652_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6905_ _7079_/CLK _6905_/D fanout516/X VGND VGND VPWR VPWR _6905_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6836_ _6925_/CLK _6836_/D fanout516/X VGND VGND VPWR VPWR _6836_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6767_ _7002_/CLK _6767_/D fanout498/X VGND VGND VPWR VPWR _6767_/Q sky130_fd_sc_hd__dfrtp_1
X_3979_ hold1/X hold99/X _3979_/S VGND VGND VPWR VPWR _3979_/X sky130_fd_sc_hd__mux2_2
XFILLER_183_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5718_ _6963_/Q _5675_/X _5677_/X _6915_/Q _5717_/X VGND VGND VPWR VPWR _5719_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6698_ _7200_/CLK _6698_/D _6348_/B VGND VGND VPWR VPWR _6698_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_40_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5649_ _7145_/Q _5648_/X _5647_/S _5649_/B2 VGND VGND VPWR VPWR _7161_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_164_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold250 _5505_/X VGND VGND VPWR VPWR _7068_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold261 _7100_/Q VGND VGND VPWR VPWR hold261/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold272 _4103_/X VGND VGND VPWR VPWR _6573_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 _6815_/Q VGND VGND VPWR VPWR hold283/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 _4260_/X VGND VGND VPWR VPWR _6712_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_101 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_112 _3949_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_123 _3949_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_134 _3960_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_145 input169/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_156 _3684_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_167 _6323_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_178 _3927_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_189 hold565/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_1_1_1_csclk/A sky130_fd_sc_hd__clkbuf_8
XFILLER_167_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput7 mask_rev_in[12] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4951_ _4951_/A _4951_/B _5060_/A VGND VGND VPWR VPWR _5059_/B sky130_fd_sc_hd__and3_1
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3902_ _7157_/Q _7158_/Q VGND VGND VPWR VPWR _6019_/A sky130_fd_sc_hd__nand2b_4
XFILLER_44_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4882_ _4882_/A _4882_/B VGND VGND VPWR VPWR _4896_/B sky130_fd_sc_hd__nand2_1
XFILLER_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6621_ _6679_/CLK _6621_/D fanout511/X VGND VGND VPWR VPWR _6621_/Q sky130_fd_sc_hd__dfrtp_4
X_3833_ _3832_/X _3833_/A1 _3833_/S VGND VGND VPWR VPWR _6463_/D sky130_fd_sc_hd__mux2_1
XFILLER_32_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6552_ _7130_/CLK _6552_/D fanout520/X VGND VGND VPWR VPWR _6552_/Q sky130_fd_sc_hd__dfrtp_1
X_3764_ _6804_/Q _5200_/A _3761_/X _3763_/X VGND VGND VPWR VPWR _3764_/X sky130_fd_sc_hd__a211o_1
X_5503_ _5521_/A0 _5503_/A1 _5510_/S VGND VGND VPWR VPWR _5503_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_530 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6483_ _6760_/CLK _6483_/D fanout490/X VGND VGND VPWR VPWR _6483_/Q sky130_fd_sc_hd__dfstp_1
X_3695_ _6931_/Q _5349_/A _5205_/A _6808_/Q VGND VGND VPWR VPWR _3695_/X sky130_fd_sc_hd__a22o_1
XFILLER_173_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput300 _6483_/Q VGND VGND VPWR VPWR pll_trim[9] sky130_fd_sc_hd__buf_12
X_5434_ _5584_/A0 hold556/X _5438_/S VGND VGND VPWR VPWR _5434_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput311 _3939_/X VGND VGND VPWR VPWR serial_resetn sky130_fd_sc_hd__buf_12
Xoutput322 hold1329/X VGND VGND VPWR VPWR hold1330/A sky130_fd_sc_hd__buf_12
Xoutput333 hold1319/X VGND VGND VPWR VPWR hold1320/A sky130_fd_sc_hd__buf_12
XFILLER_133_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput344 hold1351/X VGND VGND VPWR VPWR hold1352/A sky130_fd_sc_hd__buf_12
X_5365_ _5569_/A0 hold263/X _5366_/S VGND VGND VPWR VPWR _5365_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_3_0_csclk clkbuf_3_3_0_csclk/A VGND VGND VPWR VPWR _6970_/CLK sky130_fd_sc_hd__clkbuf_8
X_7104_ _7135_/CLK _7104_/D fanout519/X VGND VGND VPWR VPWR _7104_/Q sky130_fd_sc_hd__dfstp_1
X_4316_ hold502/X _6396_/A0 _4317_/S VGND VGND VPWR VPWR _4316_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5296_ _5581_/A0 _5296_/A1 _5303_/S VGND VGND VPWR VPWR _5296_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7035_ _7050_/CLK _7035_/D fanout498/X VGND VGND VPWR VPWR _7035_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_59_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4247_ _5476_/A0 _4247_/A1 _4251_/S VGND VGND VPWR VPWR _4247_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4178_ _5533_/A1 hold693/X _4179_/S VGND VGND VPWR VPWR _4178_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_0_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_70_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6819_ _7002_/CLK _6819_/D fanout498/X VGND VGND VPWR VPWR _6819_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_11_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3480_ _6990_/Q _3298_/Y _4010_/A _6510_/Q _3479_/X VGND VGND VPWR VPWR _3484_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_155_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5150_ _4876_/A _5035_/Y _5036_/Y _4744_/X _5039_/X VGND VGND VPWR VPWR _5174_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_170_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4101_ hold349/X _4100_/X _4103_/S VGND VGND VPWR VPWR _4101_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5081_ _4679_/B _5027_/B _5080_/X VGND VGND VPWR VPWR _5109_/C sky130_fd_sc_hd__o21ai_1
XFILLER_2_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4032_ hold743/X _5533_/A1 _4033_/S VGND VGND VPWR VPWR _4032_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_764 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5983_ _6000_/A _6040_/A VGND VGND VPWR VPWR _6021_/B sky130_fd_sc_hd__nand2_4
XFILLER_18_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4934_ _4957_/A _4933_/Y _4842_/Y VGND VGND VPWR VPWR _5065_/D sky130_fd_sc_hd__a21o_1
XFILLER_178_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4865_ _5162_/B _4865_/B _4865_/C _4865_/D VGND VGND VPWR VPWR _4866_/D sky130_fd_sc_hd__or4_1
XFILLER_20_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_12 _5358_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_23 _3410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6604_ _7209_/CLK _6604_/D fanout484/X VGND VGND VPWR VPWR _6604_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA_34 _3527_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3816_ hold72/A _3821_/S VGND VGND VPWR VPWR _3816_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_45 _3755_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_56 _5659_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4796_ _5076_/B _4784_/A _4795_/Y _4971_/A VGND VGND VPWR VPWR _4797_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_20_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_67 _5685_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_78 _6272_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6535_ _6755_/CLK _6535_/D fanout497/X VGND VGND VPWR VPWR _6535_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_89 _7083_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3747_ _6962_/Q _5385_/A _4216_/A _6670_/Q VGND VGND VPWR VPWR _3747_/X sky130_fd_sc_hd__a22o_1
X_6466_ _3487_/B2 _6466_/D _6421_/X VGND VGND VPWR VPWR hold16/A sky130_fd_sc_hd__dfrtp_1
X_3678_ input35/X _3295_/Y _4210_/A _6666_/Q _3677_/X VGND VGND VPWR VPWR _3679_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5417_ _5567_/A0 hold735/X _5420_/S VGND VGND VPWR VPWR _5417_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6397_ _6397_/A0 hold474/X _6397_/S VGND VGND VPWR VPWR _6397_/X sky130_fd_sc_hd__mux2_1
Xoutput174 _3961_/X VGND VGND VPWR VPWR irq[2] sky130_fd_sc_hd__buf_12
X_5348_ _5579_/A0 hold520/X _5348_/S VGND VGND VPWR VPWR _5348_/X sky130_fd_sc_hd__mux2_1
Xoutput185 _3215_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[19] sky130_fd_sc_hd__buf_12
Xoutput196 _3205_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[29] sky130_fd_sc_hd__buf_12
XFILLER_102_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5279_ _5459_/A0 hold325/X _5285_/S VGND VGND VPWR VPWR _5279_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7018_ _7018_/CLK _7018_/D fanout505/X VGND VGND VPWR VPWR _7018_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_102_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4650_ _5031_/A VGND VGND VPWR VPWR _4650_/Y sky130_fd_sc_hd__inv_2
Xinput10 mask_rev_in[15] VGND VGND VPWR VPWR input10/X sky130_fd_sc_hd__clkbuf_1
X_3601_ _3601_/A _3601_/B _3601_/C _3601_/D VGND VGND VPWR VPWR _3601_/X sky130_fd_sc_hd__or4_4
XFILLER_147_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput21 mask_rev_in[25] VGND VGND VPWR VPWR input21/X sky130_fd_sc_hd__clkbuf_1
XFILLER_175_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput32 mask_rev_in[6] VGND VGND VPWR VPWR input32/X sky130_fd_sc_hd__clkbuf_1
X_4581_ _4814_/A _4646_/A VGND VGND VPWR VPWR _4582_/B sky130_fd_sc_hd__or2_4
Xinput43 mgmt_gpio_in[16] VGND VGND VPWR VPWR input43/X sky130_fd_sc_hd__clkbuf_1
Xinput54 mgmt_gpio_in[26] VGND VGND VPWR VPWR input54/X sky130_fd_sc_hd__clkbuf_2
X_6320_ _6730_/Q _6320_/A2 _6320_/B1 _6620_/Q VGND VGND VPWR VPWR _6332_/A sky130_fd_sc_hd__a22o_1
Xhold805 _6757_/Q VGND VGND VPWR VPWR hold805/X sky130_fd_sc_hd__dlygate4sd3_1
X_3532_ _6725_/Q _4270_/A _4204_/A _6664_/Q VGND VGND VPWR VPWR _3532_/X sky130_fd_sc_hd__a22o_1
Xinput65 mgmt_gpio_in[36] VGND VGND VPWR VPWR _7214_/A sky130_fd_sc_hd__clkbuf_4
Xinput76 qspi_enabled VGND VGND VPWR VPWR _3921_/S sky130_fd_sc_hd__buf_6
Xhold816 _5388_/X VGND VGND VPWR VPWR _6964_/D sky130_fd_sc_hd__dlygate4sd3_1
Xinput87 spimemio_flash_io1_do VGND VGND VPWR VPWR _7213_/A sky130_fd_sc_hd__clkbuf_4
Xinput98 usr2_vdd_pwrgood VGND VGND VPWR VPWR input98/X sky130_fd_sc_hd__clkbuf_4
Xhold827 _6657_/Q VGND VGND VPWR VPWR hold827/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold838 _6947_/Q VGND VGND VPWR VPWR hold838/X sky130_fd_sc_hd__dlygate4sd3_1
X_6251_ _6522_/Q _5994_/X _5998_/Y _6762_/Q _6250_/X VGND VGND VPWR VPWR _6257_/A
+ sky130_fd_sc_hd__a221o_1
Xhold849 _5396_/X VGND VGND VPWR VPWR _6971_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3463_ _3507_/B _3538_/B VGND VGND VPWR VPWR _4294_/A sky130_fd_sc_hd__nor2_8
XFILLER_115_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5202_ _5555_/A0 hold321/X _5202_/S VGND VGND VPWR VPWR _5202_/X sky130_fd_sc_hd__mux2_1
X_6182_ _6504_/Q _6323_/A2 _6027_/D _6888_/Q _6181_/X VGND VGND VPWR VPWR _6182_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_170_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3394_ input32/X _3304_/Y _5466_/A _7040_/Q _3382_/X VGND VGND VPWR VPWR _3394_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_97_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5133_ _4999_/B _5060_/A _4670_/Y _4897_/C VGND VGND VPWR VPWR _5134_/D sky130_fd_sc_hd__a211o_1
XFILLER_69_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1505 _5753_/X VGND VGND VPWR VPWR _7164_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1516 _7167_/Q VGND VGND VPWR VPWR _5816_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1527 _7176_/Q VGND VGND VPWR VPWR _6072_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1538 _7206_/Q VGND VGND VPWR VPWR _6391_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5064_ _5064_/A _5064_/B _5064_/C _5064_/D VGND VGND VPWR VPWR _5125_/A sky130_fd_sc_hd__or4_1
Xhold1549 _7173_/Q VGND VGND VPWR VPWR _5948_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4015_ hold369/X _5534_/A1 _4015_/S VGND VGND VPWR VPWR _4015_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5966_ _6625_/Q _5661_/X _5966_/B1 _6520_/Q _5965_/X VGND VGND VPWR VPWR _5967_/D
+ sky130_fd_sc_hd__a221o_1
X_4917_ _4832_/B _5027_/A _5115_/B VGND VGND VPWR VPWR _5109_/A sky130_fd_sc_hd__o21bai_1
X_5897_ _6742_/Q _5656_/X _5670_/X hold87/A VGND VGND VPWR VPWR _5897_/X sky130_fd_sc_hd__a22o_1
XFILLER_32_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4848_ _4832_/B _4677_/B _5049_/A VGND VGND VPWR VPWR _4865_/B sky130_fd_sc_hd__o21bai_1
XFILLER_20_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4779_ _4484_/A _4668_/X _4794_/A VGND VGND VPWR VPWR _5095_/B sky130_fd_sc_hd__a21oi_1
XFILLER_181_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6518_ _6664_/CLK _6518_/D _3946_/B VGND VGND VPWR VPWR _6518_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_134_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6449_ net499_2/A _6449_/D _6404_/X VGND VGND VPWR VPWR _6449_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_40_csclk _6931_/CLK VGND VGND VPWR VPWR _6925_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_164_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_0_0_csclk clkbuf_2_1_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_1_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_87_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_55_csclk _6970_/CLK VGND VGND VPWR VPWR _7133_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_189_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5820_ _6864_/Q _5688_/X _5694_/X _7080_/Q _5819_/X VGND VGND VPWR VPWR _5825_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_34_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5751_ _6844_/Q _5691_/Y _5740_/X _5750_/X _3195_/Y VGND VGND VPWR VPWR _5751_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_15_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4702_ _4814_/C _4683_/B _4692_/B _4639_/B VGND VGND VPWR VPWR _4702_/X sky130_fd_sc_hd__o22a_1
X_5682_ _7152_/Q _5699_/B _5706_/C VGND VGND VPWR VPWR _5682_/X sky130_fd_sc_hd__and3_4
XFILLER_30_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4633_ _4638_/B _4639_/A VGND VGND VPWR VPWR _4982_/A sky130_fd_sc_hd__nor2_1
XFILLER_147_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4564_ _4588_/A _4935_/A _4605_/A VGND VGND VPWR VPWR _4666_/B sky130_fd_sc_hd__nand3b_4
Xhold602 _5393_/X VGND VGND VPWR VPWR _6969_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold613 _6991_/Q VGND VGND VPWR VPWR hold613/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6303_ _6734_/Q _5997_/Y _6015_/X _6663_/Q VGND VGND VPWR VPWR _6303_/X sky130_fd_sc_hd__a22o_1
Xhold624 _5462_/X VGND VGND VPWR VPWR _7030_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3515_ _3515_/A _3515_/B _3515_/C _3515_/D VGND VGND VPWR VPWR _3542_/B sky130_fd_sc_hd__or4_1
Xhold635 _6679_/Q VGND VGND VPWR VPWR hold635/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap354 _3333_/Y VGND VGND VPWR VPWR _4102_/S sky130_fd_sc_hd__buf_8
X_4495_ _4570_/D _4993_/A VGND VGND VPWR VPWR _5094_/A sky130_fd_sc_hd__nand2_4
Xhold646 _5317_/X VGND VGND VPWR VPWR _6901_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 _6950_/Q VGND VGND VPWR VPWR hold657/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap376 hold21/X VGND VGND VPWR VPWR _3528_/A sky130_fd_sc_hd__buf_12
Xhold668 _5281_/X VGND VGND VPWR VPWR _6869_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6234_ _6746_/Q _6322_/B1 _6030_/X _6741_/Q _6233_/X VGND VGND VPWR VPWR _6242_/B
+ sky130_fd_sc_hd__a221o_1
Xmax_cap387 _3495_/A VGND VGND VPWR VPWR _3536_/A sky130_fd_sc_hd__buf_12
Xhold679 _7071_/Q VGND VGND VPWR VPWR hold679/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap398 _6025_/A VGND VGND VPWR VPWR _6326_/A2 sky130_fd_sc_hd__buf_12
X_3446_ _3446_/A _3446_/B _3446_/C _3446_/D VGND VGND VPWR VPWR _3447_/D sky130_fd_sc_hd__or4_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6165_ _7055_/Q _5988_/X _6022_/B _6903_/Q VGND VGND VPWR VPWR _6165_/X sky130_fd_sc_hd__a22o_1
X_3377_ _5212_/A _3526_/A VGND VGND VPWR VPWR _3658_/A sky130_fd_sc_hd__nor2_8
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1302 _4319_/X VGND VGND VPWR VPWR _6761_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1313 hold1402/X VGND VGND VPWR VPWR hold1313/X sky130_fd_sc_hd__dlygate4sd3_1
X_5116_ _4454_/Y _4729_/Y _4988_/D _5092_/D _5115_/X VGND VGND VPWR VPWR _5172_/A
+ sky130_fd_sc_hd__a2111o_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6096_ _5650_/A _7176_/Q _6095_/X VGND VGND VPWR VPWR _6096_/X sky130_fd_sc_hd__a21o_1
Xhold1324 hold1324/A VGND VGND VPWR VPWR wb_dat_o[10] sky130_fd_sc_hd__buf_12
Xhold1335 hold1413/X VGND VGND VPWR VPWR hold1335/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1346 hold1346/A VGND VGND VPWR VPWR wb_dat_o[0] sky130_fd_sc_hd__buf_12
XFILLER_27_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1357 _4168_/A0 VGND VGND VPWR VPWR hold1357/X sky130_fd_sc_hd__dlygate4sd3_1
X_5047_ _5049_/A _5049_/B _5049_/C _5049_/D VGND VGND VPWR VPWR _5048_/C sky130_fd_sc_hd__or4_1
Xhold1368 hold1368/A VGND VGND VPWR VPWR wb_dat_o[24] sky130_fd_sc_hd__buf_12
XFILLER_26_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1379 _6446_/Q VGND VGND VPWR VPWR hold4/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6998_ _7050_/CLK _6998_/D fanout498/X VGND VGND VPWR VPWR _6998_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5949_ _6535_/Q _5678_/X _5686_/X _6765_/Q VGND VGND VPWR VPWR _5949_/X sky130_fd_sc_hd__a22o_1
XFILLER_185_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_558 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3300_ _3300_/A _3340_/B VGND VGND VPWR VPWR _3300_/Y sky130_fd_sc_hd__nor2_8
XFILLER_4_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4280_ hold36/X hold185/X _4281_/S VGND VGND VPWR VPWR _4280_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3231_ _6861_/Q VGND VGND VPWR VPWR _3231_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6921_ _6992_/CLK _6921_/D fanout517/X VGND VGND VPWR VPWR _6921_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6852_ _7129_/CLK _6852_/D fanout518/X VGND VGND VPWR VPWR _6852_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_90_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5803_ _6991_/Q _5697_/X _5800_/X _5802_/X VGND VGND VPWR VPWR _5803_/X sky130_fd_sc_hd__a211o_1
XFILLER_22_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6783_ _3927_/A1 _6783_/D _6434_/X VGND VGND VPWR VPWR _6783_/Q sky130_fd_sc_hd__dfrtn_1
X_3995_ _3995_/A0 _6395_/A0 _4000_/S VGND VGND VPWR VPWR _3995_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5734_ _7060_/Q _5671_/X _5688_/X _6860_/Q VGND VGND VPWR VPWR _5734_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5665_ _7018_/Q _5663_/X _5664_/X _7002_/Q VGND VGND VPWR VPWR _5665_/X sky130_fd_sc_hd__a22o_1
XFILLER_129_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4616_ _5023_/C _4694_/B VGND VGND VPWR VPWR _5019_/A sky130_fd_sc_hd__nor2_1
XFILLER_190_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5596_ _6565_/Q _5596_/B _5651_/B VGND VGND VPWR VPWR _5606_/A sky130_fd_sc_hd__or3_1
XFILLER_135_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold410 _4084_/X VGND VGND VPWR VPWR _6560_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_191_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4547_ _4547_/A _4573_/B VGND VGND VPWR VPWR _4802_/B sky130_fd_sc_hd__or2_2
Xhold421 _6552_/Q VGND VGND VPWR VPWR hold421/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 _4078_/X VGND VGND VPWR VPWR _6557_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold443 _7122_/Q VGND VGND VPWR VPWR hold443/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold454 _4329_/X VGND VGND VPWR VPWR _6770_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold465 _6885_/Q VGND VGND VPWR VPWR hold465/X sky130_fd_sc_hd__dlygate4sd3_1
X_4478_ _4672_/A VGND VGND VPWR VPWR _4478_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold476 _7069_/Q VGND VGND VPWR VPWR hold476/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 _3988_/X VGND VGND VPWR VPWR _6486_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold498 _6599_/Q VGND VGND VPWR VPWR hold498/X sky130_fd_sc_hd__dlygate4sd3_1
X_6217_ _6217_/A _6217_/B _6217_/C _6217_/D VGND VGND VPWR VPWR _6217_/X sky130_fd_sc_hd__or4_1
X_3429_ _7116_/Q _5553_/A _5544_/A _7108_/Q _3424_/X VGND VGND VPWR VPWR _3431_/C
+ sky130_fd_sc_hd__a221o_1
X_7197_ _7200_/CLK _7197_/D _6348_/B VGND VGND VPWR VPWR _7197_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_58_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6148_ _7071_/Q _6272_/B VGND VGND VPWR VPWR _6148_/X sky130_fd_sc_hd__and2_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1110 _5251_/X VGND VGND VPWR VPWR _6842_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1121 _6527_/Q VGND VGND VPWR VPWR _4036_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1132 _5433_/X VGND VGND VPWR VPWR _7004_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1143 _6900_/Q VGND VGND VPWR VPWR _5316_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6079_ _6900_/Q _6022_/B _6025_/B _7105_/Q _6078_/X VGND VGND VPWR VPWR _6084_/B
+ sky130_fd_sc_hd__a221o_1
Xhold1154 _5487_/X VGND VGND VPWR VPWR _7052_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1165 _6597_/Q VGND VGND VPWR VPWR _4131_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1176 hold1588/X VGND VGND VPWR VPWR _4072_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1187 _6799_/Q VGND VGND VPWR VPWR _5195_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1198 _4106_/X VGND VGND VPWR VPWR _6575_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_692 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3780_ input11/X _3268_/Y _4294_/A _6741_/Q _3779_/X VGND VGND VPWR VPWR _3781_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_9_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5450_ _5573_/A0 hold611/X _5456_/S VGND VGND VPWR VPWR _5450_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4401_ _4667_/C _4538_/B VGND VGND VPWR VPWR _4739_/A sky130_fd_sc_hd__nand2_2
X_5381_ _5567_/A0 hold763/X _5384_/S VGND VGND VPWR VPWR _5381_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_3_2_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A VGND VGND VPWR VPWR _7182_/CLK sky130_fd_sc_hd__clkbuf_8
X_7120_ _7135_/CLK _7120_/D fanout519/X VGND VGND VPWR VPWR _7120_/Q sky130_fd_sc_hd__dfstp_1
X_4332_ _5531_/A1 hold872/X _4335_/S VGND VGND VPWR VPWR _4332_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7051_ _7075_/CLK _7051_/D fanout515/X VGND VGND VPWR VPWR _7051_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_87_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4263_ hold615/X _5549_/A0 _4263_/S VGND VGND VPWR VPWR _4263_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6002_ _6018_/A _6038_/A VGND VGND VPWR VPWR _6002_/Y sky130_fd_sc_hd__nor2_8
XFILLER_39_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3214_ _7005_/Q VGND VGND VPWR VPWR _3214_/Y sky130_fd_sc_hd__inv_2
X_4194_ _4194_/A0 _6353_/A1 _4197_/S VGND VGND VPWR VPWR _6651_/D sky130_fd_sc_hd__mux2_1
XFILLER_94_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6904_ _6925_/CLK _6904_/D fanout516/X VGND VGND VPWR VPWR _6904_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6835_ _7049_/CLK hold15/X fanout522/X VGND VGND VPWR VPWR _6835_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_11_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6766_ _6825_/CLK _6766_/D fanout490/X VGND VGND VPWR VPWR _6766_/Q sky130_fd_sc_hd__dfrtp_1
X_3978_ hold144/X hold127/X _3982_/S VGND VGND VPWR VPWR _3978_/X sky130_fd_sc_hd__mux2_1
X_5717_ _6931_/Q _5670_/X _5705_/X _6939_/Q VGND VGND VPWR VPWR _5717_/X sky130_fd_sc_hd__a22o_1
XFILLER_183_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6697_ _7200_/CLK _6697_/D _6348_/B VGND VGND VPWR VPWR _6697_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_1__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR _3945_/A1
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_40_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5648_ _7146_/Q _7147_/Q _5648_/C _7144_/Q VGND VGND VPWR VPWR _5648_/X sky130_fd_sc_hd__or4b_1
XFILLER_156_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5579_ _5579_/A0 hold401/X _5579_/S VGND VGND VPWR VPWR _5579_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold240 _5424_/X VGND VGND VPWR VPWR _6996_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 _6816_/Q VGND VGND VPWR VPWR hold251/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 _5541_/X VGND VGND VPWR VPWR _7100_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 _6623_/Q VGND VGND VPWR VPWR hold273/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold284 _5217_/X VGND VGND VPWR VPWR _6815_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold295 hold295/A VGND VGND VPWR VPWR hold295/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_102 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_113 _3949_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_124 _3949_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_135 _3872_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_146 _3924_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_157 _3684_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_168 _5552_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_179 _3927_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput8 mask_rev_in[13] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4950_ _5064_/C _4950_/B _4950_/C VGND VGND VPWR VPWR _4954_/B sky130_fd_sc_hd__nand3b_1
XFILLER_64_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3901_ _3901_/A _5596_/B VGND VGND VPWR VPWR _6563_/D sky130_fd_sc_hd__or2_1
X_4881_ _4396_/X _4740_/Y _4453_/A VGND VGND VPWR VPWR _4885_/B sky130_fd_sc_hd__a21oi_1
XTAP_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6620_ _6725_/CLK _6620_/D fanout509/X VGND VGND VPWR VPWR _6620_/Q sky130_fd_sc_hd__dfrtp_4
X_3832_ _3830_/A input58/X hold72/A VGND VGND VPWR VPWR _3832_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_550 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6551_ _7130_/CLK _6551_/D fanout519/X VGND VGND VPWR VPWR _6551_/Q sky130_fd_sc_hd__dfrtp_1
X_3763_ input4/X _3304_/Y _5430_/A _7002_/Q _3762_/X VGND VGND VPWR VPWR _3763_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5502_ _5502_/A _5571_/B VGND VGND VPWR VPWR _5510_/S sky130_fd_sc_hd__nand2_8
XFILLER_146_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6482_ _6760_/CLK _6482_/D fanout490/X VGND VGND VPWR VPWR _6482_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_145_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3694_ input53/X _5232_/A _3335_/Y _7128_/Q _3693_/X VGND VGND VPWR VPWR _3701_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5433_ _5574_/A0 _5433_/A1 _5438_/S VGND VGND VPWR VPWR _5433_/X sky130_fd_sc_hd__mux2_1
Xoutput301 _6807_/Q VGND VGND VPWR VPWR pwr_ctrl_out[0] sky130_fd_sc_hd__buf_12
XFILLER_133_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput312 _3958_/X VGND VGND VPWR VPWR spi_sdi sky130_fd_sc_hd__buf_12
XFILLER_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput323 hold1311/X VGND VGND VPWR VPWR hold1312/A sky130_fd_sc_hd__buf_12
XFILLER_160_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput334 hold1367/X VGND VGND VPWR VPWR hold1368/A sky130_fd_sc_hd__buf_12
X_5364_ _5586_/A0 _5364_/A1 _5366_/S VGND VGND VPWR VPWR _5364_/X sky130_fd_sc_hd__mux2_1
Xoutput345 hold1321/X VGND VGND VPWR VPWR hold1322/A sky130_fd_sc_hd__buf_12
XFILLER_126_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7103_ _7130_/CLK _7103_/D fanout521/X VGND VGND VPWR VPWR _7103_/Q sky130_fd_sc_hd__dfstp_2
X_4315_ hold749/X _4327_/A1 _4317_/S VGND VGND VPWR VPWR _4315_/X sky130_fd_sc_hd__mux2_1
X_5295_ _5295_/A _5571_/B VGND VGND VPWR VPWR _5303_/S sky130_fd_sc_hd__nand2_8
X_7034_ _7137_/CLK _7034_/D fanout501/X VGND VGND VPWR VPWR _7034_/Q sky130_fd_sc_hd__dfstp_4
X_4246_ _4246_/A _4330_/B VGND VGND VPWR VPWR _4251_/S sky130_fd_sc_hd__nand2_4
XFILLER_19_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4177_ _4327_/A1 hold787/X _4179_/S VGND VGND VPWR VPWR _4177_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6818_ _7050_/CLK _6818_/D fanout499/X VGND VGND VPWR VPWR _6818_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_50_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6749_ _6963_/CLK _6749_/D fanout509/X VGND VGND VPWR VPWR _6749_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_149_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4100_ hold123/X _5569_/A0 _4102_/S VGND VGND VPWR VPWR _4100_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5080_ _5027_/A _5108_/B _4922_/B VGND VGND VPWR VPWR _5080_/X sky130_fd_sc_hd__o21ba_1
XFILLER_56_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4031_ hold830/X _4327_/A1 _4033_/S VGND VGND VPWR VPWR _4031_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5982_ _6040_/A _6039_/A _6020_/C VGND VGND VPWR VPWR _5982_/X sky130_fd_sc_hd__and3_2
XFILLER_80_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4933_ _4933_/A _4935_/C VGND VGND VPWR VPWR _4933_/Y sky130_fd_sc_hd__nor2_1
XFILLER_33_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4864_ _5064_/A _5124_/B _4864_/C _4864_/D VGND VGND VPWR VPWR _4865_/D sky130_fd_sc_hd__or4_1
XANTENNA_13 hold30/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6603_ _7209_/CLK _6603_/D fanout484/X VGND VGND VPWR VPWR _6603_/Q sky130_fd_sc_hd__dfrtp_1
X_3815_ _3814_/X _3815_/A1 _3833_/S VGND VGND VPWR VPWR _6469_/D sky130_fd_sc_hd__mux2_1
XANTENNA_24 _3410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_35 _4204_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_46 _3760_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4795_ _4802_/D _4795_/B VGND VGND VPWR VPWR _4795_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_57 _5659_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6534_ _6755_/CLK _6534_/D fanout497/X VGND VGND VPWR VPWR _6534_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_68 _5693_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_79 _6045_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3746_ _6938_/Q _5358_/A _4153_/A _6616_/Q _3745_/X VGND VGND VPWR VPWR _3749_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_192_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6465_ _3487_/B2 _6465_/D _6420_/X VGND VGND VPWR VPWR hold64/A sky130_fd_sc_hd__dfrtp_1
X_3677_ _6612_/Q _4147_/A _4135_/A _6602_/Q VGND VGND VPWR VPWR _3677_/X sky130_fd_sc_hd__a22o_1
XFILLER_173_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5416_ _5557_/A0 hold619/X _5420_/S VGND VGND VPWR VPWR _5416_/X sky130_fd_sc_hd__mux2_1
X_6396_ _6396_/A0 hold522/X _6397_/S VGND VGND VPWR VPWR _6396_/X sky130_fd_sc_hd__mux2_1
X_5347_ _5578_/A0 hold813/X _5348_/S VGND VGND VPWR VPWR _5347_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput175 _3935_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[0] sky130_fd_sc_hd__buf_12
Xoutput186 _3934_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[1] sky130_fd_sc_hd__buf_12
Xoutput197 _3231_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[2] sky130_fd_sc_hd__buf_12
XFILLER_102_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5278_ _5521_/A0 _5278_/A1 _5285_/S VGND VGND VPWR VPWR _5278_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7017_ _7126_/CLK _7017_/D fanout524/X VGND VGND VPWR VPWR _7017_/Q sky130_fd_sc_hd__dfrtp_4
X_4229_ _6699_/Q _6698_/Q _6700_/Q VGND VGND VPWR VPWR _4232_/B sky130_fd_sc_hd__or3_2
XFILLER_75_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3600_ _3600_/A _3600_/B _3600_/C _3600_/D VGND VGND VPWR VPWR _3601_/D sky130_fd_sc_hd__or4_1
Xinput11 mask_rev_in[16] VGND VGND VPWR VPWR input11/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput22 mask_rev_in[26] VGND VGND VPWR VPWR input22/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4580_ _4814_/A _4646_/A VGND VGND VPWR VPWR _4684_/B sky130_fd_sc_hd__nor2_2
Xinput33 mask_rev_in[7] VGND VGND VPWR VPWR input33/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput44 mgmt_gpio_in[17] VGND VGND VPWR VPWR input44/X sky130_fd_sc_hd__clkbuf_2
X_3531_ hold20/X _4120_/B VGND VGND VPWR VPWR _4204_/A sky130_fd_sc_hd__nor2_8
Xinput55 mgmt_gpio_in[27] VGND VGND VPWR VPWR input55/X sky130_fd_sc_hd__clkbuf_2
XFILLER_183_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput66 mgmt_gpio_in[37] VGND VGND VPWR VPWR _7215_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput77 ser_tx VGND VGND VPWR VPWR input77/X sky130_fd_sc_hd__clkbuf_1
Xhold806 _4314_/X VGND VGND VPWR VPWR _6757_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold817 _7060_/Q VGND VGND VPWR VPWR hold817/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold828 _4201_/X VGND VGND VPWR VPWR _6657_/D sky130_fd_sc_hd__dlygate4sd3_1
Xinput88 spimemio_flash_io1_oeb VGND VGND VPWR VPWR _3949_/B sky130_fd_sc_hd__clkbuf_4
X_6250_ _6512_/Q _5977_/X _6323_/B1 _6737_/Q VGND VGND VPWR VPWR _6250_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold839 _5369_/X VGND VGND VPWR VPWR _6947_/D sky130_fd_sc_hd__dlygate4sd3_1
Xinput99 wb_adr_i[0] VGND VGND VPWR VPWR _4570_/B sky130_fd_sc_hd__buf_12
X_3462_ hold57/X _3462_/B VGND VGND VPWR VPWR _4306_/A sky130_fd_sc_hd__nor2_8
X_5201_ _5536_/A1 _5201_/A1 _5202_/S VGND VGND VPWR VPWR _5201_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6181_ _7109_/Q _6025_/B _6036_/X _7040_/Q VGND VGND VPWR VPWR _6181_/X sky130_fd_sc_hd__a22o_1
X_3393_ _7072_/Q _5502_/A _5520_/A _7088_/Q _3383_/X VGND VGND VPWR VPWR _3393_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_170_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5132_ _5132_/A _5132_/B VGND VGND VPWR VPWR _5151_/B sky130_fd_sc_hd__or2_1
XFILLER_96_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1506 _7178_/Q VGND VGND VPWR VPWR _6145_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1517 _5816_/X VGND VGND VPWR VPWR _7167_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5063_ _5023_/A _5027_/A _4515_/C VGND VGND VPWR VPWR _5064_/D sky130_fd_sc_hd__o21ai_1
Xhold1528 _7202_/Q VGND VGND VPWR VPWR _6380_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1539 _6391_/X VGND VGND VPWR VPWR _7206_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4014_ hold741/X _5533_/A1 _4015_/S VGND VGND VPWR VPWR _4014_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5965_ _6659_/Q _5693_/X _5700_/X _6510_/Q VGND VGND VPWR VPWR _5965_/X sky130_fd_sc_hd__a22o_1
X_4916_ _4916_/A _4916_/B VGND VGND VPWR VPWR _5153_/A sky130_fd_sc_hd__nand2_1
XFILLER_178_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5896_ _6762_/Q _5686_/X _5694_/X _6522_/Q _5895_/X VGND VGND VPWR VPWR _5901_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4847_ _4847_/A _4882_/B VGND VGND VPWR VPWR _4847_/Y sky130_fd_sc_hd__nand2_1
XFILLER_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4778_ _4993_/A _4778_/B VGND VGND VPWR VPWR _4778_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3729_ _5212_/A _3729_/B VGND VGND VPWR VPWR _5203_/A sky130_fd_sc_hd__nor2_1
X_6517_ _6664_/CLK _6517_/D _6426_/A VGND VGND VPWR VPWR _6517_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_180_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6448_ net499_2/A _6448_/D _6403_/X VGND VGND VPWR VPWR hold34/A sky130_fd_sc_hd__dfrtp_1
XFILLER_134_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6379_ _6700_/Q _6379_/A2 _6379_/B1 _6699_/Q _6378_/X VGND VGND VPWR VPWR _6379_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_88_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5750_ _5750_/A _5750_/B _5750_/C _5750_/D VGND VGND VPWR VPWR _5750_/X sky130_fd_sc_hd__or4_1
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4701_ _4471_/B _4814_/A _4639_/B _4699_/X _4700_/X VGND VGND VPWR VPWR _4701_/X
+ sky130_fd_sc_hd__o311a_1
X_5681_ _5681_/A _5681_/B _5681_/C _5681_/D VGND VGND VPWR VPWR _5681_/X sky130_fd_sc_hd__or4_1
XFILLER_30_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4632_ _5016_/A _5027_/A VGND VGND VPWR VPWR _4987_/A sky130_fd_sc_hd__nor2_1
XFILLER_135_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4563_ _4846_/B _4563_/B VGND VGND VPWR VPWR _4718_/B sky130_fd_sc_hd__nand2_2
Xhold603 _6981_/Q VGND VGND VPWR VPWR hold603/X sky130_fd_sc_hd__dlygate4sd3_1
X_6302_ _6509_/Q _6049_/B _6006_/Y _6754_/Q VGND VGND VPWR VPWR _6302_/X sky130_fd_sc_hd__a22o_1
X_3514_ _6974_/Q _5394_/A _4324_/A _6770_/Q _3513_/X VGND VGND VPWR VPWR _3515_/D
+ sky130_fd_sc_hd__a221o_1
Xhold614 _5418_/X VGND VGND VPWR VPWR _6991_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold625 _7086_/Q VGND VGND VPWR VPWR hold625/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold636 _4227_/X VGND VGND VPWR VPWR _6679_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4494_ _4846_/C _4532_/B VGND VGND VPWR VPWR _4870_/B sky130_fd_sc_hd__nor2_4
Xmax_cap355 _3318_/Y VGND VGND VPWR VPWR _5295_/A sky130_fd_sc_hd__buf_6
Xhold647 _6886_/Q VGND VGND VPWR VPWR hold647/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 _5372_/X VGND VGND VPWR VPWR _6950_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6233_ _6716_/Q _6023_/B _6338_/B1 _6766_/Q _6221_/X VGND VGND VPWR VPWR _6233_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_171_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap377 hold20/X VGND VGND VPWR VPWR hold21/A sky130_fd_sc_hd__buf_12
X_3445_ _3445_/A _3445_/B _3445_/C _3445_/D VGND VGND VPWR VPWR _3446_/D sky130_fd_sc_hd__or4_1
XFILLER_116_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold669 _6625_/Q VGND VGND VPWR VPWR hold669/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_170_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap388 _3525_/A VGND VGND VPWR VPWR _3495_/A sky130_fd_sc_hd__buf_12
Xmax_cap399 _5997_/Y VGND VGND VPWR VPWR _6203_/A2 sky130_fd_sc_hd__buf_8
XFILLER_170_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6164_ _6855_/Q _6027_/A _6329_/B1 _7039_/Q _6163_/X VGND VGND VPWR VPWR _6167_/C
+ sky130_fd_sc_hd__a221o_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3376_ _3375_/X _3376_/A1 _3917_/A VGND VGND VPWR VPWR _6790_/D sky130_fd_sc_hd__mux2_1
XFILLER_97_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5115_ _5115_/A _5115_/B VGND VGND VPWR VPWR _5115_/X sky130_fd_sc_hd__or2_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1303 _6526_/Q VGND VGND VPWR VPWR _4035_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6095_ _6844_/Q _6046_/B _6085_/X _6094_/X _3195_/Y VGND VGND VPWR VPWR _6095_/X
+ sky130_fd_sc_hd__o221a_1
Xhold1314 hold1314/A VGND VGND VPWR VPWR wb_dat_o[17] sky130_fd_sc_hd__buf_12
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1325 hold1408/X VGND VGND VPWR VPWR hold1325/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1336 hold1336/A VGND VGND VPWR VPWR wb_dat_o[8] sky130_fd_sc_hd__buf_12
Xhold1347 _4191_/A0 VGND VGND VPWR VPWR hold1347/X sky130_fd_sc_hd__dlygate4sd3_1
X_5046_ _4516_/B _5001_/B _4746_/Y _4880_/X _5008_/C VGND VGND VPWR VPWR _5132_/A
+ sky130_fd_sc_hd__a2111o_1
XFILLER_27_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1358 hold1358/A VGND VGND VPWR VPWR wb_dat_o[18] sky130_fd_sc_hd__buf_12
XFILLER_84_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1369 _6347_/A1 VGND VGND VPWR VPWR hold1369/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6997_ _7033_/CLK _6997_/D fanout503/X VGND VGND VPWR VPWR _6997_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_25_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5948_ _5948_/A0 _5947_/X _6319_/S VGND VGND VPWR VPWR _7173_/D sky130_fd_sc_hd__mux2_1
XFILLER_178_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5879_ _5879_/A _5879_/B _5879_/C _5879_/D VGND VGND VPWR VPWR _5879_/X sky130_fd_sc_hd__or4_1
XFILLER_139_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3230_ _6877_/Q VGND VGND VPWR VPWR _3230_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6920_ _6977_/CLK _6920_/D fanout507/X VGND VGND VPWR VPWR _6920_/Q sky130_fd_sc_hd__dfrtp_2
X_6851_ _6923_/CLK _6851_/D fanout514/X VGND VGND VPWR VPWR _6851_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_23_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5802_ _6959_/Q _5659_/X _5685_/X _6911_/Q _5801_/X VGND VGND VPWR VPWR _5802_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_90_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3994_ _3994_/A0 _6394_/A0 _4000_/S VGND VGND VPWR VPWR _3994_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6782_ _7200_/CLK _6782_/D fanout529/X VGND VGND VPWR VPWR _6782_/Q sky130_fd_sc_hd__dfrtp_1
X_5733_ _7068_/Q _5678_/X _5700_/X _7028_/Q _5732_/X VGND VGND VPWR VPWR _5740_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_176_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5664_ _7152_/Q _5705_/B _5700_/C VGND VGND VPWR VPWR _5664_/X sky130_fd_sc_hd__and3_4
XFILLER_176_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_54_csclk _6970_/CLK VGND VGND VPWR VPWR _6969_/CLK sky130_fd_sc_hd__clkbuf_16
X_4615_ _4784_/B _4707_/A _5021_/B _4677_/B VGND VGND VPWR VPWR _4618_/D sky130_fd_sc_hd__o22a_1
XFILLER_135_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5595_ _5604_/D VGND VGND VPWR VPWR _5595_/Y sky130_fd_sc_hd__inv_2
XFILLER_163_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold400 _5240_/X VGND VGND VPWR VPWR _6833_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4546_ _4546_/A _4546_/B VGND VGND VPWR VPWR _4573_/B sky130_fd_sc_hd__xnor2_2
Xhold411 _6831_/Q VGND VGND VPWR VPWR hold411/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 _4067_/X VGND VGND VPWR VPWR _6552_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold433 _7118_/Q VGND VGND VPWR VPWR hold433/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 _5566_/X VGND VGND VPWR VPWR _7122_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 _6735_/Q VGND VGND VPWR VPWR hold455/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold466 _5299_/X VGND VGND VPWR VPWR _6885_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4477_ _5018_/A _4664_/A VGND VGND VPWR VPWR _4672_/A sky130_fd_sc_hd__or2_4
Xhold477 _5506_/X VGND VGND VPWR VPWR _7069_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold488 _6760_/Q VGND VGND VPWR VPWR hold488/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold499 _4133_/X VGND VGND VPWR VPWR _6599_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_69_csclk _7018_/CLK VGND VGND VPWR VPWR _7042_/CLK sky130_fd_sc_hd__clkbuf_16
X_6216_ _6216_/A _6216_/B _6216_/C _6216_/D VGND VGND VPWR VPWR _6217_/D sky130_fd_sc_hd__or4_1
X_3428_ _7015_/Q _5439_/A _5511_/A _7079_/Q _3419_/X VGND VGND VPWR VPWR _3431_/B
+ sky130_fd_sc_hd__a221o_1
X_7196_ _7196_/CLK _7196_/D VGND VGND VPWR VPWR _7196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6147_ _7132_/Q _6320_/A2 _6320_/B1 _6879_/Q VGND VGND VPWR VPWR _6147_/X sky130_fd_sc_hd__a22o_1
X_3359_ _7009_/Q _5430_/A _4085_/S _3960_/B _3358_/X VGND VGND VPWR VPWR _3359_/X
+ sky130_fd_sc_hd__a221o_1
Xhold1100 _4297_/X VGND VGND VPWR VPWR _6743_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1111 _6922_/Q VGND VGND VPWR VPWR _5341_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1122 _4036_/X VGND VGND VPWR VPWR _6527_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_161_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1133 _6733_/Q VGND VGND VPWR VPWR _4285_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_6078_ _6964_/Q _6025_/D _6212_/B1 _7044_/Q VGND VGND VPWR VPWR _6078_/X sky130_fd_sc_hd__a22o_1
Xhold1144 _5316_/X VGND VGND VPWR VPWR _6900_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1155 _7050_/Q VGND VGND VPWR VPWR _5485_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1166 _4131_/X VGND VGND VPWR VPWR _6597_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1177 _4072_/X VGND VGND VPWR VPWR _6554_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5029_ _5109_/B _5029_/B _5029_/C _5029_/D VGND VGND VPWR VPWR _5029_/X sky130_fd_sc_hd__and4b_1
Xhold1188 _5195_/X VGND VGND VPWR VPWR _6799_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1199 hold1605/X VGND VGND VPWR VPWR _5556_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4400_ _4570_/B _4400_/B VGND VGND VPWR VPWR _4742_/A sky130_fd_sc_hd__nor2_4
X_5380_ _5557_/A0 hold627/X _5384_/S VGND VGND VPWR VPWR _5380_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4331_ _5212_/C _4331_/A1 _4335_/S VGND VGND VPWR VPWR _4331_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7050_ _7050_/CLK _7050_/D fanout498/X VGND VGND VPWR VPWR _7050_/Q sky130_fd_sc_hd__dfstp_1
X_4262_ hold148/X hold36/X _4263_/S VGND VGND VPWR VPWR _4262_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6001_ _6021_/A _6019_/B VGND VGND VPWR VPWR _6025_/A sky130_fd_sc_hd__nor2_8
X_3213_ _7013_/Q VGND VGND VPWR VPWR _3213_/Y sky130_fd_sc_hd__inv_2
X_4193_ _4193_/A0 _3601_/X _4197_/S VGND VGND VPWR VPWR _6650_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6903_ _7055_/CLK _6903_/D fanout522/X VGND VGND VPWR VPWR _6903_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6834_ _6925_/CLK _6834_/D fanout522/X VGND VGND VPWR VPWR _6834_/Q sky130_fd_sc_hd__dfrtp_1
X_6765_ _7042_/CLK _6765_/D fanout491/X VGND VGND VPWR VPWR _6765_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3977_ hold125/X hold131/X _6680_/Q VGND VGND VPWR VPWR _3977_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5716_ _7003_/Q _5664_/X _5715_/X VGND VGND VPWR VPWR _5719_/C sky130_fd_sc_hd__a21o_1
XFILLER_148_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6696_ _7200_/CLK _6696_/D _6348_/B VGND VGND VPWR VPWR _6696_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_109_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5647_ _5651_/A _5647_/A1 _5647_/S VGND VGND VPWR VPWR _7160_/D sky130_fd_sc_hd__mux2_1
XFILLER_40_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5578_ _5578_/A0 hold858/X _5579_/S VGND VGND VPWR VPWR _5578_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold230 _4069_/X VGND VGND VPWR VPWR _6553_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 _6608_/Q VGND VGND VPWR VPWR hold241/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold252 _5218_/X VGND VGND VPWR VPWR _6816_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4529_ _4838_/B _4475_/A _5148_/A VGND VGND VPWR VPWR _4530_/D sky130_fd_sc_hd__a21oi_1
XFILLER_6_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold263 _6944_/Q VGND VGND VPWR VPWR hold263/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 _4162_/X VGND VGND VPWR VPWR _6623_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold285 _6810_/Q VGND VGND VPWR VPWR hold285/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold296 _4124_/X VGND VGND VPWR VPWR _6591_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7179_ _7181_/CLK _7179_/D fanout506/X VGND VGND VPWR VPWR _7179_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_58_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_103 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_114 _3949_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_125 _3949_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_136 _3872_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_147 _6801_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_158 _3684_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_169 _5558_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput9 mask_rev_in[14] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__clkbuf_1
XFILLER_76_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3900_ _6318_/S _3908_/B VGND VGND VPWR VPWR _5596_/B sky130_fd_sc_hd__nor2_1
XFILLER_32_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4880_ _4516_/B _4657_/C _4985_/B VGND VGND VPWR VPWR _4880_/X sky130_fd_sc_hd__a21o_1
XTAP_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3831_ _3831_/A _3831_/B VGND VGND VPWR VPWR _6464_/D sky130_fd_sc_hd__xnor2_1
XFILLER_32_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3762_ _6994_/Q _3300_/Y _4330_/A _6771_/Q VGND VGND VPWR VPWR _3762_/X sky130_fd_sc_hd__a22o_1
X_6550_ _7130_/CLK _6550_/D fanout519/X VGND VGND VPWR VPWR _6550_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_158_562 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5501_ _5579_/A0 hold562/X _5501_/S VGND VGND VPWR VPWR _5501_/X sky130_fd_sc_hd__mux2_1
X_6481_ _7050_/CLK _6481_/D fanout498/X VGND VGND VPWR VPWR _6481_/Q sky130_fd_sc_hd__dfstp_2
X_3693_ _7067_/Q _5502_/A hold58/A hold89/A VGND VGND VPWR VPWR _3693_/X sky130_fd_sc_hd__a22o_1
XFILLER_145_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5432_ _5555_/A0 hold357/X _5438_/S VGND VGND VPWR VPWR _5432_/X sky130_fd_sc_hd__mux2_1
Xoutput302 _6808_/Q VGND VGND VPWR VPWR pwr_ctrl_out[1] sky130_fd_sc_hd__buf_12
XFILLER_133_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput313 _3952_/X VGND VGND VPWR VPWR spimemio_flash_io0_di sky130_fd_sc_hd__buf_12
Xoutput324 hold1307/X VGND VGND VPWR VPWR hold1308/A sky130_fd_sc_hd__buf_12
X_5363_ _5567_/A0 hold675/X _5366_/S VGND VGND VPWR VPWR _5363_/X sky130_fd_sc_hd__mux2_1
Xoutput335 hold1365/X VGND VGND VPWR VPWR hold1366/A sky130_fd_sc_hd__buf_12
Xoutput346 hold1325/X VGND VGND VPWR VPWR hold1326/A sky130_fd_sc_hd__buf_12
X_7102_ _7102_/CLK _7102_/D fanout503/X VGND VGND VPWR VPWR _7102_/Q sky130_fd_sc_hd__dfrtp_4
X_4314_ hold805/X _5531_/A1 _4317_/S VGND VGND VPWR VPWR _4314_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5294_ _5579_/A0 hold397/X hold32/X VGND VGND VPWR VPWR _5294_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7033_ _7033_/CLK _7033_/D fanout504/X VGND VGND VPWR VPWR _7033_/Q sky130_fd_sc_hd__dfrtp_4
X_4245_ hold697/X _5534_/A1 _4245_/S VGND VGND VPWR VPWR _4245_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4176_ _5531_/A1 hold950/X _4179_/S VGND VGND VPWR VPWR _4176_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6817_ _7050_/CLK _6817_/D fanout499/X VGND VGND VPWR VPWR _6817_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6748_ _6963_/CLK _6748_/D fanout509/X VGND VGND VPWR VPWR _6748_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_167_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6679_ _6679_/CLK _6679_/D fanout511/X VGND VGND VPWR VPWR _6679_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_109_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4030_ hold940/X _5531_/A1 _4033_/S VGND VGND VPWR VPWR _4030_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5981_ _7082_/Q _5977_/X _6027_/A _6850_/Q VGND VGND VPWR VPWR _5981_/X sky130_fd_sc_hd__a22o_1
XFILLER_18_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4932_ _4932_/A _4932_/B VGND VGND VPWR VPWR _4935_/C sky130_fd_sc_hd__or2_1
XFILLER_17_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4863_ _4863_/A _4863_/B VGND VGND VPWR VPWR _4864_/D sky130_fd_sc_hd__nand2_1
XFILLER_33_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_14 _3355_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6602_ _7209_/CLK _6602_/D fanout484/X VGND VGND VPWR VPWR _6602_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_25 _3410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3814_ _3252_/B _3811_/S _3813_/X _3244_/X VGND VGND VPWR VPWR _3814_/X sky130_fd_sc_hd__a31o_1
XFILLER_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_36 _4204_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4794_ _4794_/A _4795_/B _4794_/C VGND VGND VPWR VPWR _5094_/B sky130_fd_sc_hd__or3_1
XANTENNA_47 _3779_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_58 _5661_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6533_ _7042_/CLK _6533_/D fanout491/X VGND VGND VPWR VPWR _6533_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA_69 _5697_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3745_ _6686_/Q _4240_/A _4246_/A _6701_/Q VGND VGND VPWR VPWR _3745_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6464_ _3487_/B2 _6464_/D _6419_/X VGND VGND VPWR VPWR hold53/A sky130_fd_sc_hd__dfrtp_1
X_3676_ _6702_/Q _4246_/A _4300_/A _6747_/Q _3675_/X VGND VGND VPWR VPWR _3679_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_134_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5415_ _5583_/A0 hold317/X _5420_/S VGND VGND VPWR VPWR _5415_/X sky130_fd_sc_hd__mux2_1
X_6395_ _6395_/A0 hold981/X _6397_/S VGND VGND VPWR VPWR _6395_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5346_ _5550_/A0 hold587/X _5348_/S VGND VGND VPWR VPWR _5346_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput176 _3224_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[10] sky130_fd_sc_hd__buf_12
Xoutput187 _3214_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[20] sky130_fd_sc_hd__buf_12
XFILLER_99_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput198 _3204_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[30] sky130_fd_sc_hd__buf_12
XFILLER_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5277_ _5277_/A _5571_/B VGND VGND VPWR VPWR _5285_/S sky130_fd_sc_hd__nand2_8
XFILLER_87_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7016_ _7098_/CLK _7016_/D fanout506/X VGND VGND VPWR VPWR _7016_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_102_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4228_ _6699_/Q _6698_/Q _6700_/Q VGND VGND VPWR VPWR _4228_/Y sky130_fd_sc_hd__nor3_1
XFILLER_28_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4159_ _4159_/A _5580_/B VGND VGND VPWR VPWR _4164_/S sky130_fd_sc_hd__and2_2
XFILLER_83_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput12 mask_rev_in[17] VGND VGND VPWR VPWR input12/X sky130_fd_sc_hd__clkbuf_1
Xinput23 mask_rev_in[27] VGND VGND VPWR VPWR input23/X sky130_fd_sc_hd__clkbuf_2
Xinput34 mask_rev_in[8] VGND VGND VPWR VPWR input34/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput45 mgmt_gpio_in[18] VGND VGND VPWR VPWR input45/X sky130_fd_sc_hd__clkbuf_2
X_3530_ _3726_/B _3530_/B VGND VGND VPWR VPWR _4270_/A sky130_fd_sc_hd__nor2_2
Xinput56 mgmt_gpio_in[28] VGND VGND VPWR VPWR input56/X sky130_fd_sc_hd__buf_2
Xinput67 mgmt_gpio_in[3] VGND VGND VPWR VPWR _3872_/C sky130_fd_sc_hd__buf_6
Xhold807 _6613_/Q VGND VGND VPWR VPWR hold807/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput78 spi_csb VGND VGND VPWR VPWR input78/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold818 _5496_/X VGND VGND VPWR VPWR _7060_/D sky130_fd_sc_hd__dlygate4sd3_1
Xinput89 spimemio_flash_io2_do VGND VGND VPWR VPWR input89/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold829 hold829/A VGND VGND VPWR VPWR hold829/X sky130_fd_sc_hd__dlygate4sd3_1
X_3461_ input48/X _3308_/Y _4288_/A _6740_/Q _3459_/X VGND VGND VPWR VPWR _3468_/C
+ sky130_fd_sc_hd__a221o_1
X_5200_ _5200_/A _6392_/B VGND VGND VPWR VPWR _5202_/S sky130_fd_sc_hd__nand2_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6180_ _6180_/A _6180_/B _6180_/C _6180_/D VGND VGND VPWR VPWR _6193_/A sky130_fd_sc_hd__or4_1
X_3392_ _3392_/A _3392_/B _3392_/C _3392_/D VGND VGND VPWR VPWR _3410_/A sky130_fd_sc_hd__or4_1
X_5131_ _4454_/Y _5001_/B _4815_/A _4878_/X _5008_/A VGND VGND VPWR VPWR _5132_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1507 _7175_/Q VGND VGND VPWR VPWR _6071_/A2 sky130_fd_sc_hd__dlygate4sd3_1
X_5062_ _5163_/B _5123_/B _5159_/A _5062_/D VGND VGND VPWR VPWR _5066_/A sky130_fd_sc_hd__nand4_1
Xhold1518 _7179_/Q VGND VGND VPWR VPWR _6146_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1529 hold99/A VGND VGND VPWR VPWR _6383_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_4013_ _4013_/A0 _6395_/A0 _4015_/S VGND VGND VPWR VPWR _4013_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5964_ _6664_/Q _5685_/X _5694_/X _6525_/Q _5963_/X VGND VGND VPWR VPWR _5967_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_52_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4915_ _4915_/A _4915_/B _4915_/C _4914_/X VGND VGND VPWR VPWR _4924_/A sky130_fd_sc_hd__or4b_1
XFILLER_178_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5895_ _6752_/Q _5664_/X _5689_/X _5894_/X VGND VGND VPWR VPWR _5895_/X sky130_fd_sc_hd__a22o_1
XFILLER_178_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4846_ _4846_/A _4846_/B _4846_/C _4846_/D VGND VGND VPWR VPWR _4868_/C sky130_fd_sc_hd__and4_1
XFILLER_193_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4777_ _5094_/A _5076_/B _4745_/A VGND VGND VPWR VPWR _5158_/B sky130_fd_sc_hd__a21oi_2
XFILLER_165_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6516_ _6664_/CLK _6516_/D _6426_/A VGND VGND VPWR VPWR _6516_/Q sky130_fd_sc_hd__dfrtp_1
X_3728_ _6866_/Q _5277_/A _4141_/A _6606_/Q VGND VGND VPWR VPWR _3728_/X sky130_fd_sc_hd__a22o_1
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6447_ net499_2/A _6447_/D _6402_/X VGND VGND VPWR VPWR hold42/A sky130_fd_sc_hd__dfrtp_1
X_3659_ _3659_/A _3659_/B _3659_/C _3659_/D VGND VGND VPWR VPWR _3660_/C sky130_fd_sc_hd__or4_1
XFILLER_164_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6378_ _6698_/Q _6378_/A2 _6378_/B1 _6390_/A2 VGND VGND VPWR VPWR _6378_/X sky130_fd_sc_hd__a22o_1
XFILLER_87_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5329_ _5329_/A0 hold2/X _5330_/S VGND VGND VPWR VPWR hold3/A sky130_fd_sc_hd__mux2_1
XFILLER_0_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_48 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4700_ _4707_/B _4704_/B _4692_/B _4683_/A VGND VGND VPWR VPWR _4700_/X sky130_fd_sc_hd__a31o_1
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5680_ _6962_/Q _5675_/X _5676_/X _7042_/Q _5679_/X VGND VGND VPWR VPWR _5681_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_187_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4631_ _5083_/A _4631_/B VGND VGND VPWR VPWR _4915_/A sky130_fd_sc_hd__nand2b_1
XFILLER_147_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4562_ _4570_/D _4596_/B VGND VGND VPWR VPWR _4569_/B sky130_fd_sc_hd__or2_2
XFILLER_116_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6301_ _6524_/Q _5994_/X _5998_/Y _6764_/Q _6299_/X VGND VGND VPWR VPWR _6301_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_156_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold604 _5407_/X VGND VGND VPWR VPWR _6981_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3513_ _6710_/Q _4252_/A _4135_/A _6605_/Q VGND VGND VPWR VPWR _3513_/X sky130_fd_sc_hd__a22o_1
Xhold615 _6715_/Q VGND VGND VPWR VPWR hold615/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold626 _5525_/X VGND VGND VPWR VPWR _7086_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4493_ _4745_/A _4832_/B VGND VGND VPWR VPWR _4493_/X sky130_fd_sc_hd__or2_1
Xhold637 _6982_/Q VGND VGND VPWR VPWR hold637/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap356 _3308_/Y VGND VGND VPWR VPWR _4068_/S sky130_fd_sc_hd__buf_8
Xhold648 _5300_/X VGND VGND VPWR VPWR _6886_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6232_ _6232_/A _6232_/B _6232_/C _6232_/D VGND VGND VPWR VPWR _6232_/X sky130_fd_sc_hd__or4_1
Xmax_cap367 _3341_/Y VGND VGND VPWR VPWR _5403_/A sky130_fd_sc_hd__buf_8
XFILLER_131_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold659 _6973_/Q VGND VGND VPWR VPWR hold659/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap378 hold95/X VGND VGND VPWR VPWR _3546_/A sky130_fd_sc_hd__buf_12
XFILLER_131_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3444_ input49/X _4068_/S _5562_/A _7124_/Q _3443_/X VGND VGND VPWR VPWR _3445_/D
+ sky130_fd_sc_hd__a221o_1
Xmax_cap389 _5212_/A VGND VGND VPWR VPWR _3731_/A sky130_fd_sc_hd__buf_12
XFILLER_131_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3375_ _3373_/X _3412_/A1 _3791_/A VGND VGND VPWR VPWR _3375_/X sky130_fd_sc_hd__mux2_1
X_6163_ _6503_/Q _6323_/A2 _6024_/B _6935_/Q VGND VGND VPWR VPWR _6163_/X sky130_fd_sc_hd__a22o_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5114_ _5114_/A _5114_/B _5114_/C _5114_/D VGND VGND VPWR VPWR _5171_/A sky130_fd_sc_hd__or4_1
Xhold1304 _4035_/X VGND VGND VPWR VPWR _6526_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6094_ _6094_/A _6094_/B _6094_/C _6094_/D VGND VGND VPWR VPWR _6094_/X sky130_fd_sc_hd__or4_1
XFILLER_111_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1315 hold1401/X VGND VGND VPWR VPWR hold1315/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1326 hold1326/A VGND VGND VPWR VPWR wb_dat_o[6] sky130_fd_sc_hd__buf_12
Xhold1337 hold1414/X VGND VGND VPWR VPWR hold1337/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1348 hold1348/A VGND VGND VPWR VPWR wb_dat_o[1] sky130_fd_sc_hd__buf_12
X_5045_ _5045_/A _5045_/B VGND VGND VPWR VPWR _5134_/C sky130_fd_sc_hd__or2_1
Xhold1359 _4170_/A0 VGND VGND VPWR VPWR hold1359/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6996_ _7068_/CLK _6996_/D fanout505/X VGND VGND VPWR VPWR _6996_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5947_ _6563_/Q _7172_/Q _5946_/X VGND VGND VPWR VPWR _5947_/X sky130_fd_sc_hd__a21o_1
XFILLER_43_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5878_ _6616_/Q _5667_/X _5694_/X _6521_/Q _5877_/X VGND VGND VPWR VPWR _5879_/D
+ sky130_fd_sc_hd__a221o_1
X_4829_ _4596_/B _4483_/A _4847_/A VGND VGND VPWR VPWR _4829_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_138_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_560 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1 hold1/A VGND VGND VPWR VPWR hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6850_ _6990_/CLK _6850_/D _3873_/A VGND VGND VPWR VPWR _6850_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5801_ _6927_/Q _5672_/X _5705_/X _6943_/Q VGND VGND VPWR VPWR _5801_/X sky130_fd_sc_hd__a22o_1
X_6781_ _3937_/A1 _6781_/D fanout529/X VGND VGND VPWR VPWR _6781_/Q sky130_fd_sc_hd__dfrtp_1
X_3993_ _3993_/A0 _6393_/A0 _4000_/S VGND VGND VPWR VPWR _3993_/X sky130_fd_sc_hd__mux2_1
X_5732_ _7004_/Q _5664_/X _5706_/X _6500_/Q VGND VGND VPWR VPWR _5732_/X sky130_fd_sc_hd__a22o_1
X_5663_ _7152_/Q _5700_/C _5699_/B VGND VGND VPWR VPWR _5663_/X sky130_fd_sc_hd__and3_4
XFILLER_148_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4614_ _4638_/B _4646_/B VGND VGND VPWR VPWR _4916_/A sky130_fd_sc_hd__or2_1
X_5594_ _6565_/Q _5650_/A _6564_/Q _5592_/Y VGND VGND VPWR VPWR _5604_/D sky130_fd_sc_hd__o31a_1
XFILLER_128_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold401 _7134_/Q VGND VGND VPWR VPWR hold401/X sky130_fd_sc_hd__dlygate4sd3_1
X_4545_ _4793_/A _4610_/A _4621_/C VGND VGND VPWR VPWR _4683_/A sky130_fd_sc_hd__or3_4
XFILLER_144_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold412 _5238_/X VGND VGND VPWR VPWR _6831_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 _7108_/Q VGND VGND VPWR VPWR hold423/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold434 _5561_/X VGND VGND VPWR VPWR _7118_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold445 _6909_/Q VGND VGND VPWR VPWR hold445/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold456 _4287_/X VGND VGND VPWR VPWR _6735_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4476_ _4588_/A _4935_/A _4605_/A _4621_/B VGND VGND VPWR VPWR _4664_/A sky130_fd_sc_hd__or4b_1
Xhold467 _6530_/Q VGND VGND VPWR VPWR hold467/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold478 _6797_/Q VGND VGND VPWR VPWR hold478/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold489 _4317_/X VGND VGND VPWR VPWR _6760_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6215_ _6857_/Q _6027_/A _6329_/B1 _7041_/Q _6214_/X VGND VGND VPWR VPWR _6216_/D
+ sky130_fd_sc_hd__a221o_1
X_3427_ _6855_/Q _5259_/A _4104_/A _7215_/A _3426_/X VGND VGND VPWR VPWR _3431_/A
+ sky130_fd_sc_hd__a221o_1
X_7195_ _7196_/CLK _7195_/D VGND VGND VPWR VPWR _7195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6146_ _6146_/A0 _6145_/X _6319_/S VGND VGND VPWR VPWR _7179_/D sky130_fd_sc_hd__mux2_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3358_ input51/X _3308_/Y _5403_/A _6985_/Q VGND VGND VPWR VPWR _3358_/X sky130_fd_sc_hd__a22o_2
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1101 _6598_/Q VGND VGND VPWR VPWR _4132_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1112 _5341_/X VGND VGND VPWR VPWR _6922_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1123 _6956_/Q VGND VGND VPWR VPWR _5379_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1134 _4285_/X VGND VGND VPWR VPWR _6733_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6077_ _6860_/Q _6025_/A wire394/X _6892_/Q _6076_/X VGND VGND VPWR VPWR _6084_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_161_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1145 _6611_/Q VGND VGND VPWR VPWR _4148_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_3289_ _3313_/B _3378_/B VGND VGND VPWR VPWR _3726_/B sky130_fd_sc_hd__nand2_8
Xhold1156 _5485_/X VGND VGND VPWR VPWR _7050_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1167 _6606_/Q VGND VGND VPWR VPWR _4142_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1178 _6731_/Q VGND VGND VPWR VPWR _4283_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5028_ _4596_/X _4781_/Y _4672_/A VGND VGND VPWR VPWR _5029_/B sky130_fd_sc_hd__a21o_1
XTAP_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1189 _6546_/Q VGND VGND VPWR VPWR _4055_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6979_ _7107_/CLK _6979_/D fanout514/X VGND VGND VPWR VPWR _6979_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_110_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold990 _5355_/X VGND VGND VPWR VPWR _6935_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_663 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4330_ _4330_/A _4330_/B VGND VGND VPWR VPWR _4335_/S sky130_fd_sc_hd__nand2_2
XFILLER_5_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4261_ hold233/X hold44/X _4263_/S VGND VGND VPWR VPWR _4261_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6000_ _6000_/A _6033_/A _6040_/B VGND VGND VPWR VPWR _6049_/B sky130_fd_sc_hd__and3_4
XFILLER_140_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3212_ _7021_/Q VGND VGND VPWR VPWR _3212_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4192_ _4192_/A0 _3660_/X _4197_/S VGND VGND VPWR VPWR _6649_/D sky130_fd_sc_hd__mux2_1
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6902_ _7082_/CLK _6902_/D _3873_/A VGND VGND VPWR VPWR _6902_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_54_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6833_ _7134_/CLK _6833_/D fanout524/X VGND VGND VPWR VPWR _6833_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_24_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6764_ _6764_/CLK _6764_/D _6426_/A VGND VGND VPWR VPWR _6764_/Q sky130_fd_sc_hd__dfrtp_4
X_3976_ hold482/X _6397_/A0 _3982_/S VGND VGND VPWR VPWR _3976_/X sky130_fd_sc_hd__mux2_1
X_5715_ _7059_/Q _5671_/X _5694_/X _7075_/Q VGND VGND VPWR VPWR _5715_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6695_ _7200_/CLK _6695_/D _6348_/B VGND VGND VPWR VPWR _6695_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_136_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5646_ _5593_/Y _5609_/Y _5645_/X _6565_/Q VGND VGND VPWR VPWR _5647_/S sky130_fd_sc_hd__a22o_1
XFILLER_163_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5577_ _5586_/A0 _5577_/A1 _5579_/S VGND VGND VPWR VPWR _5577_/X sky130_fd_sc_hd__mux2_1
Xhold220 _4156_/X VGND VGND VPWR VPWR _6618_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold231 _6814_/Q VGND VGND VPWR VPWR hold231/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4528_ _5126_/A _4847_/A _4882_/A _4528_/D VGND VGND VPWR VPWR _4530_/C sky130_fd_sc_hd__and4b_1
XFILLER_191_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold242 _4144_/X VGND VGND VPWR VPWR _6608_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 _6738_/Q VGND VGND VPWR VPWR hold253/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 _5365_/X VGND VGND VPWR VPWR _6944_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold275 _7029_/Q VGND VGND VPWR VPWR hold275/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 _5209_/X VGND VGND VPWR VPWR _6810_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4459_ _4570_/D _4459_/B VGND VGND VPWR VPWR _5035_/B sky130_fd_sc_hd__nand2_8
XFILLER_131_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold297 _6722_/Q VGND VGND VPWR VPWR hold297/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7178_ _7181_/CLK _7178_/D fanout505/X VGND VGND VPWR VPWR _7178_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_105_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6129_ _6990_/Q _5997_/Y _6024_/C _6910_/Q VGND VGND VPWR VPWR _6129_/X sky130_fd_sc_hd__a22o_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_104 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_115 _3949_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_126 _7213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_137 _3958_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_148 _6803_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_159 _3778_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_53_csclk _6970_/CLK VGND VGND VPWR VPWR _6977_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_189_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3830_ _3830_/A _3833_/S VGND VGND VPWR VPWR _3831_/B sky130_fd_sc_hd__nor2_1
XFILLER_32_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3761_ _6751_/Q _4306_/A _5229_/A _6824_/Q VGND VGND VPWR VPWR _3761_/X sky130_fd_sc_hd__a22o_1
XFILLER_158_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5500_ _5569_/A0 _5500_/A1 _5501_/S VGND VGND VPWR VPWR _5500_/X sky130_fd_sc_hd__mux2_1
XFILLER_158_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6480_ _7050_/CLK _6480_/D fanout498/X VGND VGND VPWR VPWR _6480_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3692_ _6607_/Q _4141_/A _3691_/X _3658_/A VGND VGND VPWR VPWR _3722_/A sky130_fd_sc_hd__a211o_1
XFILLER_185_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5431_ _5536_/A1 _5431_/A1 _5438_/S VGND VGND VPWR VPWR _5431_/X sky130_fd_sc_hd__mux2_1
Xoutput303 _6809_/Q VGND VGND VPWR VPWR pwr_ctrl_out[2] sky130_fd_sc_hd__buf_12
XFILLER_145_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput314 _3953_/X VGND VGND VPWR VPWR spimemio_flash_io1_di sky130_fd_sc_hd__buf_12
XFILLER_114_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5362_ _5584_/A0 hold449/X _5366_/S VGND VGND VPWR VPWR _5362_/X sky130_fd_sc_hd__mux2_1
Xoutput325 hold1363/X VGND VGND VPWR VPWR hold1364/A sky130_fd_sc_hd__buf_12
XFILLER_160_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput336 hold1353/X VGND VGND VPWR VPWR hold1354/A sky130_fd_sc_hd__buf_12
X_7101_ _7141_/CLK _7101_/D fanout504/X VGND VGND VPWR VPWR _7101_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput347 hold1331/X VGND VGND VPWR VPWR hold1332/A sky130_fd_sc_hd__buf_12
X_4313_ _4313_/A0 _5212_/C _4317_/S VGND VGND VPWR VPWR _4313_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5293_ _5569_/A0 hold117/X hold32/X VGND VGND VPWR VPWR _5293_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7032_ _7141_/CLK _7032_/D fanout504/X VGND VGND VPWR VPWR _7032_/Q sky130_fd_sc_hd__dfrtp_4
X_4244_ hold703/X _5533_/A1 _4245_/S VGND VGND VPWR VPWR _4244_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4175_ _5476_/A0 _4175_/A1 _4179_/S VGND VGND VPWR VPWR _4175_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6816_ _7050_/CLK _6816_/D fanout499/X VGND VGND VPWR VPWR _6816_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6747_ _6963_/CLK _6747_/D fanout509/X VGND VGND VPWR VPWR _6747_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_149_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3959_ _3959_/A input1/X VGND VGND VPWR VPWR _3959_/X sky130_fd_sc_hd__and2_1
XFILLER_109_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6678_ _6683_/CLK hold37/X fanout511/X VGND VGND VPWR VPWR _6678_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_137_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5629_ _7154_/Q _7153_/Q VGND VGND VPWR VPWR _6040_/A sky130_fd_sc_hd__and2b_4
XFILLER_137_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout530 _4951_/A VGND VGND VPWR VPWR _4570_/D sky130_fd_sc_hd__buf_12
XFILLER_116_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5980_ _6021_/A _6038_/B VGND VGND VPWR VPWR _5980_/Y sky130_fd_sc_hd__nor2_8
XFILLER_18_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4931_ _4931_/A _4931_/B VGND VGND VPWR VPWR _4932_/B sky130_fd_sc_hd__nor2_1
XFILLER_32_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4862_ _4862_/A _4862_/B _4862_/C _4862_/D VGND VGND VPWR VPWR _4864_/C sky130_fd_sc_hd__or4_1
XFILLER_177_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6601_ _7209_/CLK _6601_/D fanout484/X VGND VGND VPWR VPWR _6601_/Q sky130_fd_sc_hd__dfrtp_4
X_3813_ _6468_/Q _6467_/Q _3821_/S hold46/A VGND VGND VPWR VPWR _3813_/X sky130_fd_sc_hd__a31o_1
XANTENNA_15 _3355_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_26 _3410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4793_ _4793_/A _4793_/B VGND VGND VPWR VPWR _4794_/C sky130_fd_sc_hd__or2_1
XFILLER_193_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_37 _4204_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_48 _3789_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6532_ _7042_/CLK _6532_/D fanout497/X VGND VGND VPWR VPWR _6532_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_59 _5663_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3744_ _6954_/Q _5376_/A _4258_/A _6711_/Q _3743_/X VGND VGND VPWR VPWR _3749_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_186_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6463_ _3487_/B2 _6463_/D _6418_/X VGND VGND VPWR VPWR hold25/A sky130_fd_sc_hd__dfrtp_1
X_3675_ _6799_/Q _5193_/A _5184_/A _6792_/Q VGND VGND VPWR VPWR _3675_/X sky130_fd_sc_hd__a22o_1
X_5414_ _5573_/A0 hold864/X _5420_/S VGND VGND VPWR VPWR _5414_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6394_ _6394_/A0 hold983/X _6397_/S VGND VGND VPWR VPWR _6394_/X sky130_fd_sc_hd__mux2_1
X_5345_ _5549_/A0 hold751/X _5348_/S VGND VGND VPWR VPWR _5345_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput177 _3223_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[11] sky130_fd_sc_hd__buf_12
Xoutput188 _3213_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[21] sky130_fd_sc_hd__buf_12
XFILLER_102_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5276_ _5552_/A0 hold567/X _5276_/S VGND VGND VPWR VPWR _5276_/X sky130_fd_sc_hd__mux2_1
Xoutput199 _3203_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[31] sky130_fd_sc_hd__buf_12
XFILLER_101_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7015_ _7126_/CLK _7015_/D fanout524/X VGND VGND VPWR VPWR _7015_/Q sky130_fd_sc_hd__dfrtp_2
X_4227_ _5549_/A0 hold635/X hold51/X VGND VGND VPWR VPWR _4227_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4158_ _5549_/A0 hold558/X _4158_/S VGND VGND VPWR VPWR _4158_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4089_ _4089_/A0 _4088_/X _4103_/S VGND VGND VPWR VPWR _4089_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput13 mask_rev_in[18] VGND VGND VPWR VPWR input13/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput24 mask_rev_in[28] VGND VGND VPWR VPWR input24/X sky130_fd_sc_hd__clkbuf_2
XFILLER_168_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput35 mask_rev_in[9] VGND VGND VPWR VPWR input35/X sky130_fd_sc_hd__clkbuf_2
XFILLER_155_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput46 mgmt_gpio_in[19] VGND VGND VPWR VPWR input46/X sky130_fd_sc_hd__clkbuf_2
Xinput57 mgmt_gpio_in[29] VGND VGND VPWR VPWR input57/X sky130_fd_sc_hd__clkbuf_1
Xinput68 mgmt_gpio_in[5] VGND VGND VPWR VPWR _3957_/A sky130_fd_sc_hd__buf_4
XFILLER_143_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold808 _4150_/X VGND VGND VPWR VPWR _6613_/D sky130_fd_sc_hd__dlygate4sd3_1
Xinput79 spi_enabled VGND VGND VPWR VPWR _3958_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_6_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold819 _6972_/Q VGND VGND VPWR VPWR hold819/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3460_ hold96/X _3538_/B VGND VGND VPWR VPWR _4288_/A sky130_fd_sc_hd__nor2_4
XFILLER_143_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3391_ input9/X _3295_/Y _5448_/A _7024_/Q _3385_/X VGND VGND VPWR VPWR _3392_/D
+ sky130_fd_sc_hd__a221o_2
XFILLER_170_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5130_ _5130_/A _5130_/B _5130_/C _5050_/X VGND VGND VPWR VPWR _5148_/C sky130_fd_sc_hd__or4b_1
XFILLER_35_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1508 _7186_/Q VGND VGND VPWR VPWR _6319_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5061_ _5158_/C _5127_/C VGND VGND VPWR VPWR _5062_/D sky130_fd_sc_hd__nor2_1
XFILLER_38_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1519 _7197_/Q VGND VGND VPWR VPWR _6365_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_4012_ hold934/X _5531_/A1 _4015_/S VGND VGND VPWR VPWR _4012_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5963_ _6745_/Q _5656_/X _5682_/X _6515_/Q VGND VGND VPWR VPWR _5963_/X sky130_fd_sc_hd__a22o_1
X_4914_ _4675_/A _4692_/B _4912_/X _4913_/X _4713_/A VGND VGND VPWR VPWR _4914_/X
+ sky130_fd_sc_hd__o2111a_1
X_5894_ _6712_/Q _5938_/B VGND VGND VPWR VPWR _5894_/X sky130_fd_sc_hd__or2_1
XFILLER_80_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4845_ _4871_/A _4832_/B _4745_/A VGND VGND VPWR VPWR _4930_/C sky130_fd_sc_hd__a21oi_1
XFILLER_178_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4776_ _4536_/Y _4723_/X _4775_/X _4232_/X _4776_/B2 VGND VGND VPWR VPWR _6776_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_165_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6515_ _7094_/CLK _6515_/D fanout494/X VGND VGND VPWR VPWR _6515_/Q sky130_fd_sc_hd__dfrtp_2
X_3727_ _5212_/A _5212_/B VGND VGND VPWR VPWR _3727_/Y sky130_fd_sc_hd__nor2_1
XFILLER_174_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6446_ net499_2/A _6446_/D _6401_/X VGND VGND VPWR VPWR _6446_/Q sky130_fd_sc_hd__dfrtp_1
X_3658_ _3658_/A _3658_/B _3658_/C _3658_/D VGND VGND VPWR VPWR _3659_/D sky130_fd_sc_hd__or4_1
XFILLER_161_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6377_ _6376_/X _6377_/A1 _6386_/S VGND VGND VPWR VPWR _7201_/D sky130_fd_sc_hd__mux2_1
X_3589_ _6485_/Q _3983_/A _4306_/A _6754_/Q _3551_/X VGND VGND VPWR VPWR _3593_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_88_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5328_ hold995/X _5586_/A0 _5330_/S VGND VGND VPWR VPWR _5328_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5259_ _5259_/A _5571_/B VGND VGND VPWR VPWR _5267_/S sky130_fd_sc_hd__nand2_8
XFILLER_87_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4630_ _5021_/B _5017_/A VGND VGND VPWR VPWR _4631_/B sky130_fd_sc_hd__or2_2
XFILLER_147_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4561_ _4570_/D _4596_/B VGND VGND VPWR VPWR _4563_/B sky130_fd_sc_hd__nor2_2
XFILLER_190_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6300_ _6539_/Q _5988_/X _6022_/B _6658_/Q _6297_/X VGND VGND VPWR VPWR _6315_/A
+ sky130_fd_sc_hd__a221o_1
X_3512_ _3726_/B _3714_/B VGND VGND VPWR VPWR _4135_/A sky130_fd_sc_hd__nor2_4
XFILLER_116_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold605 _6917_/Q VGND VGND VPWR VPWR hold605/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold616 _4263_/X VGND VGND VPWR VPWR _6715_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4492_ _5023_/A _5018_/A _5021_/A VGND VGND VPWR VPWR _4926_/A sky130_fd_sc_hd__or3_1
Xhold627 _6957_/Q VGND VGND VPWR VPWR hold627/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold638 _5408_/X VGND VGND VPWR VPWR _6982_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6231_ _6711_/Q _6009_/X _6038_/Y _6721_/Q _6230_/X VGND VGND VPWR VPWR _6232_/D
+ sky130_fd_sc_hd__a221o_1
Xhold649 _7006_/Q VGND VGND VPWR VPWR hold649/X sky130_fd_sc_hd__dlygate4sd3_1
X_3443_ _7039_/Q _5466_/A hold31/A _6879_/Q VGND VGND VPWR VPWR _3443_/X sky130_fd_sc_hd__a22o_1
XFILLER_170_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap368 _3334_/Y VGND VGND VPWR VPWR _5331_/A sky130_fd_sc_hd__buf_8
Xmax_cap379 hold95/X VGND VGND VPWR VPWR hold96/A sky130_fd_sc_hd__buf_12
XFILLER_131_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6162_ _6863_/Q _6025_/A _6027_/D _6887_/Q _6161_/X VGND VGND VPWR VPWR _6167_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ _6456_/Q _6543_/Q VGND VGND VPWR VPWR _3917_/A sky130_fd_sc_hd__nand2_4
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5113_ _4995_/A _5094_/A _4646_/X VGND VGND VPWR VPWR _5114_/D sky130_fd_sc_hd__o21ai_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6093_ _7028_/Q _6049_/B _6090_/X _6092_/X VGND VGND VPWR VPWR _6094_/D sky130_fd_sc_hd__a211o_1
XFILLER_112_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1305 hold1396/X VGND VGND VPWR VPWR hold1305/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1316 hold1316/A VGND VGND VPWR VPWR wb_dat_o[19] sky130_fd_sc_hd__buf_12
Xhold1327 hold1410/X VGND VGND VPWR VPWR hold1327/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _5136_/A _5044_/B _5130_/C _5174_/B VGND VGND VPWR VPWR _5044_/X sky130_fd_sc_hd__or4_1
Xhold1338 hold1338/A VGND VGND VPWR VPWR wb_dat_o[27] sky130_fd_sc_hd__buf_12
Xhold1349 _6353_/A0 VGND VGND VPWR VPWR hold1349/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6995_ _7115_/CLK _6995_/D fanout498/X VGND VGND VPWR VPWR _6995_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_25_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5946_ _6599_/Q _5691_/Y _5935_/X _5945_/X _6318_/S VGND VGND VPWR VPWR _5946_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_40_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5877_ _6761_/Q _5686_/X _5699_/X _6536_/Q VGND VGND VPWR VPWR _5877_/X sky130_fd_sc_hd__a22o_1
XFILLER_139_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4828_ _4570_/D _4459_/B _4485_/A _4675_/Y VGND VGND VPWR VPWR _4828_/X sky130_fd_sc_hd__a31o_1
XFILLER_193_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4759_ _4759_/A _4759_/B VGND VGND VPWR VPWR _4759_/Y sky130_fd_sc_hd__nand2_1
XFILLER_107_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6429_ _6432_/A _6441_/B VGND VGND VPWR VPWR _6429_/X sky130_fd_sc_hd__and2_1
XFILLER_134_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2 hold2/A VGND VGND VPWR VPWR hold2/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_67_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5800_ _7039_/Q _5696_/X _5700_/X _7031_/Q _5796_/X VGND VGND VPWR VPWR _5800_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_23_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6780_ _3937_/A1 _6780_/D fanout529/X VGND VGND VPWR VPWR _6780_/Q sky130_fd_sc_hd__dfrtp_1
X_3992_ _3992_/A _6392_/B VGND VGND VPWR VPWR _4000_/S sky130_fd_sc_hd__and2_2
X_5731_ _5731_/A0 _5730_/X _6319_/S VGND VGND VPWR VPWR _5731_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5662_ _6954_/Q _5659_/X _5846_/A2 _6882_/Q _5657_/X VGND VGND VPWR VPWR _5681_/A
+ sky130_fd_sc_hd__a221o_2
XFILLER_175_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4613_ _4814_/A _5021_/B VGND VGND VPWR VPWR _4646_/B sky130_fd_sc_hd__or2_2
XFILLER_148_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5593_ _6565_/Q _5650_/A VGND VGND VPWR VPWR _5593_/Y sky130_fd_sc_hd__nor2_1
XFILLER_129_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4544_ _4935_/A _4819_/C VGND VGND VPWR VPWR _4595_/B sky130_fd_sc_hd__and2b_4
Xhold402 _5579_/X VGND VGND VPWR VPWR _7134_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold413 _6569_/Q VGND VGND VPWR VPWR hold413/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold424 _5550_/X VGND VGND VPWR VPWR _7108_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 _7061_/Q VGND VGND VPWR VPWR hold435/X sky130_fd_sc_hd__dlygate4sd3_1
X_4475_ _4475_/A _5060_/A VGND VGND VPWR VPWR _4530_/A sky130_fd_sc_hd__nand2_1
Xhold446 _5326_/X VGND VGND VPWR VPWR _6909_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold457 _6877_/Q VGND VGND VPWR VPWR hold457/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 _4039_/X VGND VGND VPWR VPWR _6530_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6214_ _6505_/Q _6323_/A2 _6024_/B _6937_/Q VGND VGND VPWR VPWR _6214_/X sky130_fd_sc_hd__a22o_1
Xhold479 _5192_/X VGND VGND VPWR VPWR _6797_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3426_ _6847_/Q _5250_/A _3684_/B1 _7055_/Q VGND VGND VPWR VPWR _3426_/X sky130_fd_sc_hd__a22o_1
X_7194_ _3937_/A1 _7194_/D VGND VGND VPWR VPWR _7194_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6145_ _6145_/A0 _6144_/X _6318_/S VGND VGND VPWR VPWR _6145_/X sky130_fd_sc_hd__mux2_1
X_3357_ _6961_/Q _3320_/Y _5385_/A _6969_/Q _3356_/X VGND VGND VPWR VPWR _3357_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1102 _4132_/X VGND VGND VPWR VPWR _6598_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1113 _6508_/Q VGND VGND VPWR VPWR _4013_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6076_ _7084_/Q _5977_/X _6329_/B1 _7036_/Q VGND VGND VPWR VPWR _6076_/X sky130_fd_sc_hd__a22o_1
Xhold1124 _5379_/X VGND VGND VPWR VPWR _6956_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3288_ hold55/X hold27/X VGND VGND VPWR VPWR _3378_/B sky130_fd_sc_hd__and2_4
Xhold1135 _6931_/Q VGND VGND VPWR VPWR _5351_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1146 _4148_/X VGND VGND VPWR VPWR _6611_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5027_ _5027_/A _5027_/B VGND VGND VPWR VPWR _5109_/B sky130_fd_sc_hd__nor2_1
Xhold1157 _6736_/Q VGND VGND VPWR VPWR _4289_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1168 _4142_/X VGND VGND VPWR VPWR _6606_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1179 _4283_/X VGND VGND VPWR VPWR _6731_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6978_ _6990_/CLK _6978_/D _3873_/A VGND VGND VPWR VPWR _6978_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_186_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5929_ _6764_/Q _5686_/X _5688_/X _6609_/Q VGND VGND VPWR VPWR _5929_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold980 _5228_/X VGND VGND VPWR VPWR _6823_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold991 _6879_/Q VGND VGND VPWR VPWR hold991/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_675 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4260_ hold293/X _5459_/A0 _4263_/S VGND VGND VPWR VPWR _4260_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3211_ _7029_/Q VGND VGND VPWR VPWR _3211_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4191_ _4191_/A0 _3723_/X _4197_/S VGND VGND VPWR VPWR _6648_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6901_ _7108_/CLK _6901_/D fanout523/X VGND VGND VPWR VPWR _6901_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_47_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6832_ _7134_/CLK _6832_/D fanout524/X VGND VGND VPWR VPWR _6832_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6763_ _6764_/CLK _6763_/D _3946_/B VGND VGND VPWR VPWR _6763_/Q sky130_fd_sc_hd__dfstp_4
X_3975_ hold83/X _3975_/A1 _3981_/S VGND VGND VPWR VPWR hold84/A sky130_fd_sc_hd__mux2_4
X_5714_ _7083_/Q _5682_/X _5683_/X _6867_/Q _5713_/X VGND VGND VPWR VPWR _5719_/B
+ sky130_fd_sc_hd__a221o_1
X_6694_ _7200_/CLK _6694_/D _6348_/B VGND VGND VPWR VPWR _6694_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_148_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5645_ _7146_/Q _7147_/Q _5600_/Y VGND VGND VPWR VPWR _5645_/X sky130_fd_sc_hd__or3b_1
XFILLER_148_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5576_ hold85/X hold171/X _5579_/S VGND VGND VPWR VPWR _5576_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold210 _4125_/X VGND VGND VPWR VPWR _6592_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold221 _6723_/Q VGND VGND VPWR VPWR hold221/X sky130_fd_sc_hd__dlygate4sd3_1
X_4527_ _4738_/A _4872_/A _4832_/B _4940_/A _4525_/X VGND VGND VPWR VPWR _4528_/D
+ sky130_fd_sc_hd__o221a_1
Xhold232 _5216_/X VGND VGND VPWR VPWR _6814_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold243 _6496_/Q VGND VGND VPWR VPWR hold243/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold254 _4291_/X VGND VGND VPWR VPWR _6738_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 hold265/A VGND VGND VPWR VPWR hold265/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold276 _5461_/X VGND VGND VPWR VPWR _7029_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4458_ _4846_/C _4738_/A VGND VGND VPWR VPWR _5001_/B sky130_fd_sc_hd__nor2_4
Xhold287 _7020_/Q VGND VGND VPWR VPWR hold287/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold298 _4272_/X VGND VGND VPWR VPWR _6722_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3409_ _3658_/A _3409_/B _3409_/C _3409_/D VGND VGND VPWR VPWR _3410_/B sky130_fd_sc_hd__or4_1
XFILLER_131_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7177_ _7181_/CLK _7177_/D fanout505/X VGND VGND VPWR VPWR _7177_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_58_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4389_ _4654_/A _4547_/A VGND VGND VPWR VPWR _4674_/A sky130_fd_sc_hd__nor2_8
XFILLER_131_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6128_ _7030_/Q _6049_/B _6202_/B1 _7006_/Q VGND VGND VPWR VPWR _6128_/X sky130_fd_sc_hd__a22o_1
XFILLER_100_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6059_ _7128_/Q _6320_/A2 _6320_/B1 _6875_/Q _6050_/X VGND VGND VPWR VPWR _6059_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_100_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_105 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_116 _3949_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_127 _7213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_138 input45/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_149 _6796_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3760_ _3760_/A _3760_/B _3760_/C _3760_/D VGND VGND VPWR VPWR _3760_/X sky130_fd_sc_hd__or4_4
XFILLER_158_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3691_ _6899_/Q hold22/A hold31/A _6875_/Q _3690_/X VGND VGND VPWR VPWR _3691_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_185_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5430_ _5430_/A _5535_/B VGND VGND VPWR VPWR _5438_/S sky130_fd_sc_hd__nand2_8
XFILLER_145_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput304 _6810_/Q VGND VGND VPWR VPWR pwr_ctrl_out[3] sky130_fd_sc_hd__buf_12
XFILLER_161_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5361_ _5574_/A0 _5361_/A1 _5366_/S VGND VGND VPWR VPWR _5361_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput315 _7214_/X VGND VGND VPWR VPWR spimemio_flash_io2_di sky130_fd_sc_hd__buf_12
XFILLER_99_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput326 hold1313/X VGND VGND VPWR VPWR hold1314/A sky130_fd_sc_hd__buf_12
XFILLER_114_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput337 hold1337/X VGND VGND VPWR VPWR hold1338/A sky130_fd_sc_hd__buf_12
X_4312_ _4312_/A _4330_/B VGND VGND VPWR VPWR _4317_/S sky130_fd_sc_hd__and2_2
X_7100_ _7102_/CLK _7100_/D fanout503/X VGND VGND VPWR VPWR _7100_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_160_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput348 hold1335/X VGND VGND VPWR VPWR hold1336/A sky130_fd_sc_hd__buf_12
XFILLER_113_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5292_ _5586_/A0 hold991/X hold32/X VGND VGND VPWR VPWR _5292_/X sky130_fd_sc_hd__mux2_1
X_7031_ _7031_/CLK _7031_/D fanout526/X VGND VGND VPWR VPWR _7031_/Q sky130_fd_sc_hd__dfrtp_1
X_4243_ hold789/X _4327_/A1 _4245_/S VGND VGND VPWR VPWR _4243_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4174_ _4174_/A _4330_/B VGND VGND VPWR VPWR _4179_/S sky130_fd_sc_hd__nand2_2
XFILLER_28_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6815_ _7050_/CLK _6815_/D fanout499/X VGND VGND VPWR VPWR _6815_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_51_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6746_ _7070_/CLK _6746_/D fanout510/X VGND VGND VPWR VPWR _6746_/Q sky130_fd_sc_hd__dfrtp_4
X_3958_ _3958_/A _3958_/B VGND VGND VPWR VPWR _3958_/X sky130_fd_sc_hd__and2_1
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6677_ _6683_/CLK hold52/X fanout511/X VGND VGND VPWR VPWR _6677_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_137_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3889_ _6696_/Q _3876_/X _3888_/B _3888_/A VGND VGND VPWR VPWR _6696_/D sky130_fd_sc_hd__a22o_1
XFILLER_149_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5628_ _6564_/Q _7154_/Q _7153_/Q VGND VGND VPWR VPWR _5637_/B sky130_fd_sc_hd__and3_1
XFILLER_164_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5559_ _5586_/A0 hold993/X _5561_/S VGND VGND VPWR VPWR _5559_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout520 fanout521/X VGND VGND VPWR VPWR fanout520/X sky130_fd_sc_hd__buf_8
XFILLER_59_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_1_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A VGND VGND VPWR VPWR _7187_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_27_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4930_ _4930_/A _4964_/A _4930_/C VGND VGND VPWR VPWR _5068_/B sky130_fd_sc_hd__or3_1
XFILLER_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4861_ _4639_/B _4707_/B _4510_/A VGND VGND VPWR VPWR _4862_/D sky130_fd_sc_hd__o21ai_1
XTAP_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6600_ _6759_/CLK _6600_/D fanout489/X VGND VGND VPWR VPWR _6600_/Q sky130_fd_sc_hd__dfstp_2
X_3812_ _3833_/S _3811_/X _3810_/Y VGND VGND VPWR VPWR _6470_/D sky130_fd_sc_hd__o21ai_1
XANTENNA_16 _3355_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4792_ _4792_/A _4792_/B _4792_/C VGND VGND VPWR VPWR _4795_/B sky130_fd_sc_hd__or3_1
XFILLER_193_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_27 _3447_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_38 _3539_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6531_ _7042_/CLK _6531_/D fanout497/X VGND VGND VPWR VPWR _6531_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_49 _4128_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3743_ _6681_/Q hold58/A hold50/A _6675_/Q VGND VGND VPWR VPWR _3743_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3674_ _3731_/A hold68/X VGND VGND VPWR VPWR _5184_/A sky130_fd_sc_hd__nor2_2
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6462_ _3927_/A1 _6462_/D _6417_/X VGND VGND VPWR VPWR _6462_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_146_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5413_ _5212_/C _5413_/A1 _5420_/S VGND VGND VPWR VPWR _5413_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6393_ _6393_/A0 hold969/X _6397_/S VGND VGND VPWR VPWR _6393_/X sky130_fd_sc_hd__mux2_1
X_5344_ hold36/X hold195/X _5348_/S VGND VGND VPWR VPWR _5344_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput178 _3222_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[12] sky130_fd_sc_hd__buf_12
Xoutput189 _3212_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[22] sky130_fd_sc_hd__buf_12
X_5275_ _5587_/A0 hold842/X _5276_/S VGND VGND VPWR VPWR _5275_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4226_ hold36/X _4226_/A1 hold51/X VGND VGND VPWR VPWR hold37/A sky130_fd_sc_hd__mux2_1
X_7014_ _7130_/CLK _7014_/D fanout519/X VGND VGND VPWR VPWR _7014_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4157_ hold36/X hold169/X _4158_/S VGND VGND VPWR VPWR _4157_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4088_ hold918/X _5581_/A0 _4102_/S VGND VGND VPWR VPWR _4088_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6729_ _6740_/CLK _6729_/D _3873_/A VGND VGND VPWR VPWR _6729_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_177_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_52_csclk _6970_/CLK VGND VGND VPWR VPWR _7088_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_124_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_67_csclk _6970_/CLK VGND VGND VPWR VPWR _7012_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_132_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput14 mask_rev_in[19] VGND VGND VPWR VPWR input14/X sky130_fd_sc_hd__clkbuf_1
Xinput25 mask_rev_in[29] VGND VGND VPWR VPWR input25/X sky130_fd_sc_hd__clkbuf_1
Xinput36 mgmt_gpio_in[0] VGND VGND VPWR VPWR _3959_/A sky130_fd_sc_hd__clkbuf_4
Xinput47 mgmt_gpio_in[1] VGND VGND VPWR VPWR input47/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput58 mgmt_gpio_in[2] VGND VGND VPWR VPWR input58/X sky130_fd_sc_hd__buf_12
Xinput69 mgmt_gpio_in[6] VGND VGND VPWR VPWR input69/X sky130_fd_sc_hd__clkbuf_1
XFILLER_182_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold809 _6920_/Q VGND VGND VPWR VPWR hold809/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3390_ _6904_/Q hold22/A _4102_/S input41/X _3389_/X VGND VGND VPWR VPWR _3392_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_123_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5060_ _5060_/A _5060_/B VGND VGND VPWR VPWR _5127_/C sky130_fd_sc_hd__and2_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1509 _7180_/Q VGND VGND VPWR VPWR _6195_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4011_ _4011_/A0 _5212_/C _4015_/S VGND VGND VPWR VPWR _4011_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5962_ _6690_/Q _5666_/X _5675_/X _6710_/Q _5961_/X VGND VGND VPWR VPWR _5967_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_18_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4913_ _4400_/B _5013_/A _5108_/A _5023_/B VGND VGND VPWR VPWR _4913_/X sky130_fd_sc_hd__o22a_1
X_5893_ _6666_/Q _5677_/X _5703_/X _6602_/Q _5892_/X VGND VGND VPWR VPWR _5901_/A
+ sky130_fd_sc_hd__a221o_1
X_4844_ _4926_/A _5050_/B VGND VGND VPWR VPWR _5068_/A sky130_fd_sc_hd__nand2_1
XFILLER_178_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4775_ _4899_/B _4875_/B _4773_/X _4774_/Y _4992_/C VGND VGND VPWR VPWR _4775_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_193_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6514_ _7094_/CLK _6514_/D fanout494/X VGND VGND VPWR VPWR _6514_/Q sky130_fd_sc_hd__dfrtp_2
X_3726_ hold96/X _3726_/B VGND VGND VPWR VPWR _5223_/A sky130_fd_sc_hd__nor2_1
XFILLER_119_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6445_ _3945_/A1 _6445_/D _6400_/X VGND VGND VPWR VPWR _6445_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_161_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3657_ _3731_/A _3525_/B _4135_/A _6603_/Q VGND VGND VPWR VPWR _3658_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_174_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3588_ _3588_/A _3588_/B _3588_/C _3588_/D VGND VGND VPWR VPWR _3601_/B sky130_fd_sc_hd__or4_1
X_6376_ _6700_/Q _6376_/A2 _6376_/B1 _6699_/Q _6375_/X VGND VGND VPWR VPWR _6376_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_88_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5327_ hold633/X _5549_/A0 _5330_/S VGND VGND VPWR VPWR _5327_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5258_ hold595/X _5552_/A0 _5258_/S VGND VGND VPWR VPWR _5258_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4209_ hold461/X _6397_/A0 _4209_/S VGND VGND VPWR VPWR _4209_/X sky130_fd_sc_hd__mux2_1
X_5189_ _6394_/A0 _5189_/A1 _5192_/S VGND VGND VPWR VPWR _5189_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4560_ _4560_/A _4573_/B VGND VGND VPWR VPWR _4794_/A sky130_fd_sc_hd__nand2_2
XFILLER_128_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3511_ _4111_/B _3530_/B VGND VGND VPWR VPWR _4252_/A sky130_fd_sc_hd__nor2_8
X_4491_ _4739_/A _4871_/A VGND VGND VPWR VPWR _4993_/B sky130_fd_sc_hd__nand2_1
Xhold606 _5335_/X VGND VGND VPWR VPWR _6917_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold617 _6514_/Q VGND VGND VPWR VPWR hold617/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold628 _5380_/X VGND VGND VPWR VPWR _6957_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6230_ _6701_/Q _6336_/A2 _6033_/X _7207_/Q VGND VGND VPWR VPWR _6230_/X sky130_fd_sc_hd__a22o_1
X_3442_ _6919_/Q _5331_/A _5193_/A _6803_/Q _3441_/X VGND VGND VPWR VPWR _3445_/C
+ sky130_fd_sc_hd__a221o_1
Xhold639 _7046_/Q VGND VGND VPWR VPWR hold639/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap358 _3278_/Y VGND VGND VPWR VPWR _5553_/A sky130_fd_sc_hd__buf_6
XFILLER_171_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap369 hold77/X VGND VGND VPWR VPWR hold78/A sky130_fd_sc_hd__buf_12
XFILLER_170_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3373_ _3373_/A _3373_/B _3373_/C VGND VGND VPWR VPWR _3373_/X sky130_fd_sc_hd__or3_4
XFILLER_69_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6161_ _6951_/Q _6024_/A _6212_/B1 _7047_/Q VGND VGND VPWR VPWR _6161_/X sky130_fd_sc_hd__a22o_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5112_ _5112_/A _5112_/B _5112_/C _5112_/D VGND VGND VPWR VPWR _5140_/B sky130_fd_sc_hd__or4_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6092_ _7137_/Q _6308_/A2 _6338_/B1 _7097_/Q _6091_/X VGND VGND VPWR VPWR _6092_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1306 hold1306/A VGND VGND VPWR VPWR wb_dat_o[22] sky130_fd_sc_hd__buf_12
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1317 hold1404/X VGND VGND VPWR VPWR hold1317/X sky130_fd_sc_hd__dlygate4sd3_1
X_5043_ _4999_/B _4448_/B _4506_/Y _4984_/B _5007_/B VGND VGND VPWR VPWR _5174_/B
+ sky130_fd_sc_hd__a2111o_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1328 hold1328/A VGND VGND VPWR VPWR wb_dat_o[12] sky130_fd_sc_hd__buf_12
XFILLER_84_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1339 _6356_/A0 VGND VGND VPWR VPWR hold1339/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_0_wbbd_sck _7205_/Q VGND VGND VPWR VPWR clkbuf_0_wbbd_sck/X sky130_fd_sc_hd__clkbuf_16
X_6994_ _7115_/CLK _6994_/D fanout498/X VGND VGND VPWR VPWR _6994_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_80_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5945_ _5945_/A _5945_/B _5945_/C _5945_/D VGND VGND VPWR VPWR _5945_/X sky130_fd_sc_hd__or4_1
XFILLER_43_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5876_ _6621_/Q _5661_/X _5678_/X _6531_/Q _5875_/X VGND VGND VPWR VPWR _5879_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4827_ _4832_/B _4679_/B _4510_/C VGND VGND VPWR VPWR _5064_/B sky130_fd_sc_hd__o21ai_1
XFILLER_178_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4758_ _4758_/A _4758_/B _4758_/C _4971_/B VGND VGND VPWR VPWR _4758_/Y sky130_fd_sc_hd__nand4_2
XFILLER_193_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3709_ _6915_/Q _5331_/A _4085_/S input47/X _3708_/X VGND VGND VPWR VPWR _3710_/D
+ sky130_fd_sc_hd__a221o_1
X_4689_ _5023_/A _4689_/B VGND VGND VPWR VPWR _4689_/X sky130_fd_sc_hd__or2_1
XFILLER_162_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6428_ _6433_/A _6441_/B VGND VGND VPWR VPWR _6428_/X sky130_fd_sc_hd__and2_1
XFILLER_162_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6359_ _6700_/Q _6357_/Y _6358_/Y _6698_/Q VGND VGND VPWR VPWR _6362_/C sky130_fd_sc_hd__a22o_1
XFILLER_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold3 hold3/A VGND VGND VPWR VPWR hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_35_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3991_ _3991_/A0 _5552_/A0 _3991_/S VGND VGND VPWR VPWR _3991_/X sky130_fd_sc_hd__mux2_1
X_5730_ _5650_/A _7162_/Q _5729_/X VGND VGND VPWR VPWR _5730_/X sky130_fd_sc_hd__a21o_1
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5661_ _5938_/B _5700_/C _5703_/C VGND VGND VPWR VPWR _5661_/X sky130_fd_sc_hd__and3_4
XFILLER_176_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4612_ _4784_/B _5018_/C VGND VGND VPWR VPWR _4618_/C sky130_fd_sc_hd__or2_1
XFILLER_176_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5592_ _5650_/A _5592_/B VGND VGND VPWR VPWR _5592_/Y sky130_fd_sc_hd__nand2_2
XFILLER_191_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4543_ _4935_/A _4588_/A VGND VGND VPWR VPWR _4621_/C sky130_fd_sc_hd__nand2b_1
XFILLER_7_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold403 _6559_/Q VGND VGND VPWR VPWR hold403/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold414 _4095_/X VGND VGND VPWR VPWR _6569_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold425 _6547_/Q VGND VGND VPWR VPWR hold425/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold436 _5497_/X VGND VGND VPWR VPWR _7061_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4474_ _4474_/A _4839_/B VGND VGND VPWR VPWR _5060_/A sky130_fd_sc_hd__nor2_4
Xhold447 _7138_/Q VGND VGND VPWR VPWR hold447/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold458 _5290_/X VGND VGND VPWR VPWR _6877_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6213_ _6865_/Q _6025_/A _6027_/D _6889_/Q _6212_/X VGND VGND VPWR VPWR _6216_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold469 _7204_/Q VGND VGND VPWR VPWR hold469/X sky130_fd_sc_hd__dlygate4sd3_1
X_3425_ input17/X _3268_/Y _3992_/A _6495_/Q VGND VGND VPWR VPWR _3425_/X sky130_fd_sc_hd__a22o_2
X_7193_ _7193_/CLK _7193_/D VGND VGND VPWR VPWR _7193_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_131_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3356_ _7033_/Q _5457_/A _3340_/Y input28/X VGND VGND VPWR VPWR _3356_/X sky130_fd_sc_hd__a22o_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6144_ _6127_/X _6133_/X _6143_/X _6046_/B _6846_/Q VGND VGND VPWR VPWR _6144_/X
+ sky130_fd_sc_hd__o32a_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1103 _6518_/Q VGND VGND VPWR VPWR _4025_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1114 _4013_/X VGND VGND VPWR VPWR _6508_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3287_ _3536_/A _5241_/B VGND VGND VPWR VPWR _4001_/A sky130_fd_sc_hd__nor2_4
X_6075_ _7129_/Q _6320_/A2 _6320_/B1 _6876_/Q _6074_/X VGND VGND VPWR VPWR _6085_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1125 _6876_/Q VGND VGND VPWR VPWR _5289_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1136 _5351_/X VGND VGND VPWR VPWR _6931_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1147 _7105_/Q VGND VGND VPWR VPWR _5547_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5026_ _4677_/B _4659_/B _4679_/B _5027_/B VGND VGND VPWR VPWR _5029_/D sky130_fd_sc_hd__a31o_1
Xhold1158 _4289_/X VGND VGND VPWR VPWR _6736_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1169 _6773_/Q VGND VGND VPWR VPWR _4333_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6977_ _6977_/CLK _6977_/D fanout507/X VGND VGND VPWR VPWR _6977_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_53_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5928_ _6744_/Q _5656_/X _5678_/X _6534_/Q _5927_/X VGND VGND VPWR VPWR _5935_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_22_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5859_ _5650_/A _7168_/Q _5858_/X VGND VGND VPWR VPWR _5859_/X sky130_fd_sc_hd__a21o_1
XFILLER_186_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_76 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold970 _6393_/X VGND VGND VPWR VPWR _7207_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold981 _7209_/Q VGND VGND VPWR VPWR hold981/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_134_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold992 _5292_/X VGND VGND VPWR VPWR _6879_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3210_ _7037_/Q VGND VGND VPWR VPWR _3210_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4190_ _4190_/A0 _3790_/X _4197_/S VGND VGND VPWR VPWR _6647_/D sky130_fd_sc_hd__mux2_1
XFILLER_140_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_671 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6900_ _7129_/CLK _6900_/D fanout518/X VGND VGND VPWR VPWR _6900_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_63_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6831_ _7134_/CLK _6831_/D fanout524/X VGND VGND VPWR VPWR _6831_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6762_ _6764_/CLK _6762_/D _6426_/A VGND VGND VPWR VPWR _6762_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3974_ hold528/X _6396_/A0 _3982_/S VGND VGND VPWR VPWR _3974_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5713_ _6987_/Q _5697_/X _5702_/X _6979_/Q VGND VGND VPWR VPWR _5713_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6693_ _7200_/CLK _6693_/D _6348_/B VGND VGND VPWR VPWR _6693_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_148_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5644_ _6564_/Q _5642_/X _5643_/Y _7158_/Q VGND VGND VPWR VPWR _7158_/D sky130_fd_sc_hd__a22o_1
XFILLER_164_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5575_ _5584_/A0 hold691/X _5579_/S VGND VGND VPWR VPWR _5575_/X sky130_fd_sc_hd__mux2_1
Xhold200 _5308_/X VGND VGND VPWR VPWR _6893_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_191_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold211 _6718_/Q VGND VGND VPWR VPWR hold211/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4526_ _4872_/A _5035_/B VGND VGND VPWR VPWR _4843_/A sky130_fd_sc_hd__nor2_1
XFILLER_191_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold222 _4273_/X VGND VGND VPWR VPWR _6723_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold233 _6713_/Q VGND VGND VPWR VPWR hold233/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 _3999_/X VGND VGND VPWR VPWR _6496_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 _7115_/Q VGND VGND VPWR VPWR hold255/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 _5538_/X VGND VGND VPWR VPWR _7097_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4457_ _4759_/B _4657_/C VGND VGND VPWR VPWR _4504_/B sky130_fd_sc_hd__nand2_1
XFILLER_171_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold277 _7037_/Q VGND VGND VPWR VPWR hold277/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 _5451_/X VGND VGND VPWR VPWR _7020_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold299 _6747_/Q VGND VGND VPWR VPWR hold299/X sky130_fd_sc_hd__dlygate4sd3_1
X_3408_ _3408_/A _3408_/B _3408_/C _3408_/D VGND VGND VPWR VPWR _3409_/D sky130_fd_sc_hd__or4_1
X_7176_ _7181_/CLK _7176_/D fanout505/X VGND VGND VPWR VPWR _7176_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_172_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4388_ _4390_/A _4654_/A VGND VGND VPWR VPWR _4467_/C sky130_fd_sc_hd__nor2_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6127_ _7078_/Q _5994_/X _5998_/Y _7014_/Q _6125_/X VGND VGND VPWR VPWR _6127_/X
+ sky130_fd_sc_hd__a221o_2
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3339_ _3528_/A hold29/X VGND VGND VPWR VPWR hold30/A sky130_fd_sc_hd__nor2_4
XFILLER_85_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6058_ _6058_/A _6058_/B _6058_/C _6058_/D VGND VGND VPWR VPWR _6069_/B sky130_fd_sc_hd__or4_1
XFILLER_39_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5009_ _5009_/A _5045_/B _5049_/D _5009_/D VGND VGND VPWR VPWR _5010_/D sky130_fd_sc_hd__or4_1
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_106 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_117 _3949_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_128 _7213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_139 _3961_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3690_ _7104_/Q _5544_/A _4276_/A _6727_/Q VGND VGND VPWR VPWR _3690_/X sky130_fd_sc_hd__a22o_1
XFILLER_187_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput305 _3730_/X VGND VGND VPWR VPWR reset sky130_fd_sc_hd__buf_12
X_5360_ _5573_/A0 hold904/X _5366_/S VGND VGND VPWR VPWR _5360_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput316 _7215_/X VGND VGND VPWR VPWR spimemio_flash_io3_di sky130_fd_sc_hd__buf_12
Xoutput327 hold1357/X VGND VGND VPWR VPWR hold1358/A sky130_fd_sc_hd__buf_12
X_4311_ _5534_/A1 hold767/X _4311_/S VGND VGND VPWR VPWR _4311_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput338 hold1349/X VGND VGND VPWR VPWR hold1350/A sky130_fd_sc_hd__buf_12
Xoutput349 hold1333/X VGND VGND VPWR VPWR hold1334/A sky130_fd_sc_hd__buf_12
XFILLER_126_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5291_ hold85/X hold189/X hold32/X VGND VGND VPWR VPWR _5291_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7030_ _7043_/CLK _7030_/D fanout514/X VGND VGND VPWR VPWR _7030_/Q sky130_fd_sc_hd__dfrtp_2
X_4242_ hold908/X _5531_/A1 _4245_/S VGND VGND VPWR VPWR _4242_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4173_ _4173_/A0 _3373_/X _4173_/S VGND VGND VPWR VPWR _6633_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6814_ _7050_/CLK _6814_/D fanout499/X VGND VGND VPWR VPWR _6814_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_51_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6745_ _7211_/CLK _6745_/D fanout485/X VGND VGND VPWR VPWR _6745_/Q sky130_fd_sc_hd__dfrtp_4
X_3957_ _3957_/A _3957_/B VGND VGND VPWR VPWR _3957_/X sky130_fd_sc_hd__and2_1
XFILLER_176_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6676_ _6683_/CLK hold88/X fanout511/X VGND VGND VPWR VPWR hold87/A sky130_fd_sc_hd__dfrtp_4
X_3888_ _3888_/A _3888_/B VGND VGND VPWR VPWR _3888_/Y sky130_fd_sc_hd__nand2_1
XFILLER_176_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5627_ _7154_/Q _7153_/Q VGND VGND VPWR VPWR _6033_/A sky130_fd_sc_hd__and2_2
XFILLER_136_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5558_ _5558_/A0 hold255/X _5561_/S VGND VGND VPWR VPWR _5558_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4509_ _4512_/B _5001_/B VGND VGND VPWR VPWR _4510_/C sky130_fd_sc_hd__nand2_1
XFILLER_132_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5489_ _5549_/A0 hold701/X _5492_/S VGND VGND VPWR VPWR _5489_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout510 fanout511/X VGND VGND VPWR VPWR fanout510/X sky130_fd_sc_hd__buf_6
XFILLER_104_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout521 fanout526/X VGND VGND VPWR VPWR fanout521/X sky130_fd_sc_hd__buf_6
X_7159_ _7182_/CLK _7159_/D fanout499/X VGND VGND VPWR VPWR _7159_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_58_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4860_ _4860_/A _4860_/B _4860_/C _4860_/D VGND VGND VPWR VPWR _4862_/C sky130_fd_sc_hd__nand4_1
XTAP_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3811_ hold92/A hold93/A _3811_/S VGND VGND VPWR VPWR _3811_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4791_ _4994_/A _4802_/A _5076_/B _5027_/A VGND VGND VPWR VPWR _4987_/C sky130_fd_sc_hd__o22ai_1
XANTENNA_17 _3373_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_28 _4294_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6530_ _7207_/CLK _6530_/D fanout488/X VGND VGND VPWR VPWR _6530_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_39 _3550_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3742_ _6882_/Q _5295_/A _5259_/A _6850_/Q _3741_/X VGND VGND VPWR VPWR _3749_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_158_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6461_ _3945_/A1 _6461_/D _6416_/X VGND VGND VPWR VPWR _6461_/Q sky130_fd_sc_hd__dfrtp_4
X_3673_ _6955_/Q _5376_/A _4270_/A _6722_/Q _3672_/X VGND VGND VPWR VPWR _3679_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5412_ _5412_/A _5535_/B VGND VGND VPWR VPWR _5420_/S sky130_fd_sc_hd__nand2_8
XFILLER_161_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6392_ _6392_/A _6392_/B VGND VGND VPWR VPWR _6397_/S sky130_fd_sc_hd__nand2_2
XFILLER_173_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5343_ _5574_/A0 _5343_/A1 _5348_/S VGND VGND VPWR VPWR _5343_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput179 _3221_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[13] sky130_fd_sc_hd__buf_12
X_5274_ _5550_/A0 hold589/X _5276_/S VGND VGND VPWR VPWR _5274_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7013_ _7136_/CLK _7013_/D fanout521/X VGND VGND VPWR VPWR _7013_/Q sky130_fd_sc_hd__dfrtp_4
X_4225_ hold44/X _4225_/A1 hold51/X VGND VGND VPWR VPWR hold52/A sky130_fd_sc_hd__mux2_1
X_4156_ hold44/X hold219/X _4158_/S VGND VGND VPWR VPWR _4156_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4087_ _5241_/B _6407_/B _4052_/X _3333_/Y _5580_/B VGND VGND VPWR VPWR _4103_/S
+ sky130_fd_sc_hd__o221a_4
XFILLER_24_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4989_ _4980_/X _5119_/B _4989_/C _4989_/D VGND VGND VPWR VPWR _4990_/B sky130_fd_sc_hd__and4bb_1
X_6728_ _6990_/CLK _6728_/D _3873_/A VGND VGND VPWR VPWR _6728_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_137_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6659_ _6709_/CLK _6659_/D fanout494/X VGND VGND VPWR VPWR _6659_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_109_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput15 mask_rev_in[1] VGND VGND VPWR VPWR input15/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput26 mask_rev_in[2] VGND VGND VPWR VPWR input26/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_167_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput37 mgmt_gpio_in[10] VGND VGND VPWR VPWR input37/X sky130_fd_sc_hd__clkbuf_2
Xinput48 mgmt_gpio_in[20] VGND VGND VPWR VPWR input48/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput59 mgmt_gpio_in[30] VGND VGND VPWR VPWR input59/X sky130_fd_sc_hd__buf_2
XFILLER_128_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4010_ _4010_/A _4330_/B VGND VGND VPWR VPWR _4015_/S sky130_fd_sc_hd__and2_2
XFILLER_37_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5961_ _6540_/Q _5699_/X _5960_/X _5689_/X VGND VGND VPWR VPWR _5961_/X sky130_fd_sc_hd__a22o_1
X_4912_ _4666_/B _4692_/B _4910_/X _4911_/X _4646_/X VGND VGND VPWR VPWR _4912_/X
+ sky130_fd_sc_hd__o2111a_1
X_5892_ _6671_/Q _5955_/A2 _5693_/X _6656_/Q VGND VGND VPWR VPWR _5892_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4843_ _4843_/A _4843_/B VGND VGND VPWR VPWR _4866_/C sky130_fd_sc_hd__or2_1
X_4774_ _5050_/B _4992_/B VGND VGND VPWR VPWR _4774_/Y sky130_fd_sc_hd__nand2_1
XFILLER_193_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6513_ _7093_/CLK _6513_/D _6432_/A VGND VGND VPWR VPWR _6513_/Q sky130_fd_sc_hd__dfstp_1
X_3725_ _3724_/X _3725_/A1 _3917_/A VGND VGND VPWR VPWR _3725_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6444_ _3945_/A1 _6444_/D _6399_/X VGND VGND VPWR VPWR _6444_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3656_ _6508_/Q _4010_/A _4022_/A _6518_/Q _3655_/X VGND VGND VPWR VPWR _3658_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6375_ _6698_/Q _6375_/A2 _6375_/B1 _6390_/A2 VGND VGND VPWR VPWR _6375_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3587_ _6514_/Q _4016_/A _5187_/A _6796_/Q _3550_/X VGND VGND VPWR VPWR _3588_/D
+ sky130_fd_sc_hd__a221o_1
X_5326_ hold445/X _5584_/A0 _5330_/S VGND VGND VPWR VPWR _5326_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5257_ hold801/X _5587_/A0 _5258_/S VGND VGND VPWR VPWR _5257_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4208_ hold494/X _6396_/A0 _4209_/S VGND VGND VPWR VPWR _4208_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5188_ _6393_/A0 _5188_/A1 _5192_/S VGND VGND VPWR VPWR _5188_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4139_ hold546/X _6396_/A0 _4140_/S VGND VGND VPWR VPWR _4139_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3510_ _3536_/A _4120_/B VGND VGND VPWR VPWR _4324_/A sky130_fd_sc_hd__nor2_4
XFILLER_128_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4490_ _4872_/A _4942_/A VGND VGND VPWR VPWR _4490_/X sky130_fd_sc_hd__or2_2
Xhold607 _6965_/Q VGND VGND VPWR VPWR hold607/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold618 _4020_/X VGND VGND VPWR VPWR _6514_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold629 _6730_/Q VGND VGND VPWR VPWR hold629/X sky130_fd_sc_hd__dlygate4sd3_1
X_3441_ _6967_/Q _5385_/A _5430_/A _7007_/Q VGND VGND VPWR VPWR _3441_/X sky130_fd_sc_hd__a22o_1
XFILLER_143_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6160_ _6927_/Q _6027_/B wire394/X _6895_/Q _6159_/X VGND VGND VPWR VPWR _6167_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3372_ _3372_/A _3372_/B VGND VGND VPWR VPWR _3373_/C sky130_fd_sc_hd__or2_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5111_ _6780_/Q _6362_/A _5070_/Y _5110_/X VGND VGND VPWR VPWR _5139_/A sky130_fd_sc_hd__a22o_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ _7076_/Q _5994_/X wire412/X _6916_/Q VGND VGND VPWR VPWR _6091_/X sky130_fd_sc_hd__a22o_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1307 hold1397/X VGND VGND VPWR VPWR hold1307/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1318 hold1318/A VGND VGND VPWR VPWR wb_dat_o[30] sky130_fd_sc_hd__buf_12
X_5042_ _5042_/A _5042_/B _5042_/C VGND VGND VPWR VPWR _5130_/C sky130_fd_sc_hd__or3_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1329 hold1409/X VGND VGND VPWR VPWR hold1329/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6993_ _7080_/CLK _6993_/D fanout502/X VGND VGND VPWR VPWR _6993_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_51_csclk _6970_/CLK VGND VGND VPWR VPWR _7098_/CLK sky130_fd_sc_hd__clkbuf_16
X_5944_ _6774_/Q _5663_/X _5670_/X _6678_/Q _5943_/X VGND VGND VPWR VPWR _5945_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_80_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5875_ _6506_/Q _5700_/X _5705_/X _6681_/Q VGND VGND VPWR VPWR _5875_/X sky130_fd_sc_hd__a22o_1
XFILLER_61_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4826_ _4814_/C _4707_/B _4515_/B VGND VGND VPWR VPWR _5064_/A sky130_fd_sc_hd__o21ai_1
XFILLER_21_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4757_ _4981_/B _5094_/A _4424_/Y VGND VGND VPWR VPWR _4761_/C sky130_fd_sc_hd__a21oi_1
XFILLER_181_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3708_ _7112_/Q _3278_/Y _4216_/A _6671_/Q VGND VGND VPWR VPWR _3708_/X sky130_fd_sc_hd__a22o_1
XFILLER_107_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4688_ _5021_/A _5016_/A _5021_/C VGND VGND VPWR VPWR _4713_/B sky130_fd_sc_hd__or3_1
XFILLER_107_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6427_ _6433_/A _6441_/B VGND VGND VPWR VPWR _6427_/X sky130_fd_sc_hd__and2_1
XFILLER_146_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3639_ _7044_/Q hold77/A _5221_/B _6815_/Q _3638_/X VGND VGND VPWR VPWR _3642_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_161_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6358_ _6358_/A _6358_/B VGND VGND VPWR VPWR _6358_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5309_ _5567_/A0 hold663/X _5312_/S VGND VGND VPWR VPWR _5309_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6289_ _6538_/Q _5988_/X _6022_/B _6657_/Q VGND VGND VPWR VPWR _6289_/X sky130_fd_sc_hd__a22o_1
XFILLER_102_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_19_csclk _6820_/CLK VGND VGND VPWR VPWR _7070_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_140_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__1134_ clkbuf_0__1134_/X VGND VGND VPWR VPWR _4185_/A1 sky130_fd_sc_hd__clkbuf_16
XFILLER_138_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold4 hold4/A VGND VGND VPWR VPWR hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_81_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3990_ hold257/X _5569_/A0 _3991_/S VGND VGND VPWR VPWR _3990_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5660_ _7149_/Q _7148_/Q VGND VGND VPWR VPWR _5703_/C sky130_fd_sc_hd__and2b_2
XFILLER_31_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4611_ _4814_/A _4653_/C VGND VGND VPWR VPWR _5024_/A sky130_fd_sc_hd__or2_2
X_5591_ _5650_/A _6564_/Q VGND VGND VPWR VPWR _5651_/B sky130_fd_sc_hd__nor2_1
XFILLER_129_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4542_ _4542_/A _4792_/A VGND VGND VPWR VPWR _4546_/B sky130_fd_sc_hd__nand2_1
Xhold404 _4082_/X VGND VGND VPWR VPWR _6559_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire390 _3255_/X VGND VGND VPWR VPWR _5212_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_128_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold415 _7089_/Q VGND VGND VPWR VPWR hold415/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold426 _4057_/X VGND VGND VPWR VPWR _6547_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4473_ _4944_/A _4947_/A VGND VGND VPWR VPWR _4839_/B sky130_fd_sc_hd__or2_2
Xhold437 _7106_/Q VGND VGND VPWR VPWR hold437/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 _5584_/X VGND VGND VPWR VPWR _7138_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold459 _6774_/Q VGND VGND VPWR VPWR hold459/X sky130_fd_sc_hd__dlygate4sd3_1
X_6212_ _6953_/Q _6024_/A _6212_/B1 _7049_/Q VGND VGND VPWR VPWR _6212_/X sky130_fd_sc_hd__a22o_1
X_3424_ input40/X _4102_/S _5322_/A _6911_/Q VGND VGND VPWR VPWR _3424_/X sky130_fd_sc_hd__a22o_1
X_7192_ _7196_/CLK _7192_/D VGND VGND VPWR VPWR _7192_/Q sky130_fd_sc_hd__dfxtp_1
X_6143_ _6292_/A _6143_/B _6143_/C VGND VGND VPWR VPWR _6143_/X sky130_fd_sc_hd__or3_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3355_ _3355_/A _3355_/B _3355_/C _3355_/D VGND VGND VPWR VPWR _3373_/A sky130_fd_sc_hd__or4_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1104 _4025_/X VGND VGND VPWR VPWR _6518_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6074_ _7020_/Q _6204_/A2 _6027_/B _6924_/Q _6073_/X VGND VGND VPWR VPWR _6074_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3286_ _5241_/B VGND VGND VPWR VPWR _3286_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1115 _6746_/Q VGND VGND VPWR VPWR _4301_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1126 _5289_/X VGND VGND VPWR VPWR _6876_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1137 _7092_/Q VGND VGND VPWR VPWR _5532_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5025_ _4582_/B _5108_/A _5024_/A _5027_/B VGND VGND VPWR VPWR _5029_/C sky130_fd_sc_hd__a31o_1
Xhold1148 _5547_/X VGND VGND VPWR VPWR _7105_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1159 _6484_/Q VGND VGND VPWR VPWR _3986_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6976_ _7065_/CLK _6976_/D fanout517/X VGND VGND VPWR VPWR _6976_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_41_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5927_ _6619_/Q _5667_/X _5675_/X _6709_/Q VGND VGND VPWR VPWR _5927_/X sky130_fd_sc_hd__a22o_1
XFILLER_139_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5858_ _6849_/Q _5691_/Y _5847_/X _5857_/X _6318_/S VGND VGND VPWR VPWR _5858_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_179_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4809_ _5095_/B _4809_/B _4809_/C VGND VGND VPWR VPWR _4810_/B sky130_fd_sc_hd__and3b_1
XFILLER_166_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5789_ _7070_/Q _5678_/X _5682_/X _7086_/Q _5788_/X VGND VGND VPWR VPWR _5792_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_166_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold960 _6751_/Q VGND VGND VPWR VPWR hold960/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold971 _6826_/Q VGND VGND VPWR VPWR hold971/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold982 _6395_/X VGND VGND VPWR VPWR _7209_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold993 _7116_/Q VGND VGND VPWR VPWR hold993/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6830_ _7138_/CLK hold86/X fanout524/X VGND VGND VPWR VPWR _6830_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6761_ _6764_/CLK _6761_/D _6426_/A VGND VGND VPWR VPWR _6761_/Q sky130_fd_sc_hd__dfrtp_2
X_3973_ hold34/X hold158/X _3981_/S VGND VGND VPWR VPWR _3973_/X sky130_fd_sc_hd__mux2_4
X_5712_ _6955_/Q _5659_/X _5700_/X _7027_/Q _5711_/X VGND VGND VPWR VPWR _5719_/A
+ sky130_fd_sc_hd__a221o_1
X_6692_ _7200_/CLK _6692_/D _6348_/B VGND VGND VPWR VPWR _6692_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5643_ _5643_/A _5643_/B VGND VGND VPWR VPWR _5643_/Y sky130_fd_sc_hd__nor2_1
XFILLER_129_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5574_ _5574_/A0 _5574_/A1 _5579_/S VGND VGND VPWR VPWR _5574_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold201 _7038_/Q VGND VGND VPWR VPWR hold201/X sky130_fd_sc_hd__dlygate4sd3_1
X_4525_ _4738_/A _4997_/A _4490_/X _4522_/X _4524_/Y VGND VGND VPWR VPWR _4525_/X
+ sky130_fd_sc_hd__o2111a_1
Xhold212 _4267_/X VGND VGND VPWR VPWR _6718_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 _6872_/Q VGND VGND VPWR VPWR hold223/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 _4261_/X VGND VGND VPWR VPWR _6713_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 _7012_/Q VGND VGND VPWR VPWR hold245/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold256 _5558_/X VGND VGND VPWR VPWR _7115_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4456_ _4456_/A _4724_/B VGND VGND VPWR VPWR _4997_/A sky130_fd_sc_hd__or2_4
XFILLER_131_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold267 _6908_/Q VGND VGND VPWR VPWR hold267/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold278 _5470_/X VGND VGND VPWR VPWR _7037_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3407_ input18/X _3268_/Y _5232_/A input59/X _3406_/X VGND VGND VPWR VPWR _3408_/D
+ sky130_fd_sc_hd__a221o_1
Xhold289 _6607_/Q VGND VGND VPWR VPWR hold289/X sky130_fd_sc_hd__dlygate4sd3_1
X_7175_ _7183_/CLK _7175_/D fanout505/X VGND VGND VPWR VPWR _7175_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_132_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4387_ _4570_/B _4999_/B VGND VGND VPWR VPWR _4981_/B sky130_fd_sc_hd__nand2_8
XFILLER_86_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6126_ _6902_/Q _6022_/B _6025_/D _6966_/Q _6124_/X VGND VGND VPWR VPWR _6142_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3338_ _3528_/A hold76/X VGND VGND VPWR VPWR _5259_/A sky130_fd_sc_hd__nor2_8
XFILLER_85_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6057_ _6971_/Q _6009_/X _6206_/B1 _6979_/Q _6056_/X VGND VGND VPWR VPWR _6058_/D
+ sky130_fd_sc_hd__a221o_1
X_3269_ _3971_/S hold93/X hold47/X VGND VGND VPWR VPWR hold94/A sky130_fd_sc_hd__o21ai_1
XFILLER_45_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5008_ _5008_/A _5008_/B _5008_/C _5008_/D VGND VGND VPWR VPWR _5009_/D sky130_fd_sc_hd__or4_1
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_107 input93/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_118 _3949_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_129 _7213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6959_ _7049_/CLK _6959_/D fanout522/X VGND VGND VPWR VPWR _6959_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold790 _4243_/X VGND VGND VPWR VPWR _6688_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1490 _7195_/Q VGND VGND VPWR VPWR _6355_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_2_0__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR _3927_/A1
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput306 _3957_/X VGND VGND VPWR VPWR ser_rx sky130_fd_sc_hd__buf_12
Xoutput317 hold1369/X VGND VGND VPWR VPWR wb_ack_o sky130_fd_sc_hd__buf_12
X_4310_ _6396_/A0 hold719/X _4311_/S VGND VGND VPWR VPWR _4310_/X sky130_fd_sc_hd__mux2_1
Xoutput328 hold1315/X VGND VGND VPWR VPWR hold1316/A sky130_fd_sc_hd__buf_12
Xoutput339 hold1361/X VGND VGND VPWR VPWR hold1362/A sky130_fd_sc_hd__buf_12
X_5290_ _5584_/A0 hold457/X hold32/X VGND VGND VPWR VPWR _5290_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4241_ _4241_/A0 _5476_/A0 _4245_/S VGND VGND VPWR VPWR _4241_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4172_ _4172_/A0 _3410_/X _4173_/S VGND VGND VPWR VPWR _6632_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6813_ _7050_/CLK _6813_/D fanout499/X VGND VGND VPWR VPWR _6813_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6744_ _7211_/CLK _6744_/D fanout488/X VGND VGND VPWR VPWR _6744_/Q sky130_fd_sc_hd__dfrtp_4
X_3956_ _6699_/Q _3962_/B VGND VGND VPWR VPWR _6693_/D sky130_fd_sc_hd__and2_1
X_6675_ _6683_/CLK _6675_/D fanout511/X VGND VGND VPWR VPWR _6675_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_167_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3887_ _3887_/A _3887_/B _3887_/C _3887_/D VGND VGND VPWR VPWR _3887_/Y sky130_fd_sc_hd__nor4_1
X_5626_ _5610_/X _5650_/B _7153_/Q VGND VGND VPWR VPWR _7153_/D sky130_fd_sc_hd__mux2_1
XFILLER_137_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5557_ _5557_/A0 hold575/X _5561_/S VGND VGND VPWR VPWR _5557_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4508_ _4871_/A _4995_/A _4447_/Y _4505_/X _4507_/X VGND VGND VPWR VPWR _4508_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_132_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5488_ _5584_/A0 hold542/X _5492_/S VGND VGND VPWR VPWR _5488_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4439_ _4453_/C _4456_/A VGND VGND VPWR VPWR _4996_/A sky130_fd_sc_hd__or2_4
Xfanout500 fanout508/X VGND VGND VPWR VPWR fanout500/X sky130_fd_sc_hd__buf_4
XFILLER_116_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout511 fanout527/X VGND VGND VPWR VPWR fanout511/X sky130_fd_sc_hd__buf_8
XFILLER_132_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout522 fanout523/X VGND VGND VPWR VPWR fanout522/X sky130_fd_sc_hd__buf_8
X_7158_ _7182_/CLK _7158_/D fanout502/X VGND VGND VPWR VPWR _7158_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6109_ _6109_/A _6109_/B _6109_/C _6109_/D VGND VGND VPWR VPWR _6110_/B sky130_fd_sc_hd__or4_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7089_ _7108_/CLK _7089_/D fanout523/X VGND VGND VPWR VPWR _7089_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_86_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3810_ _3810_/A _3833_/S VGND VGND VPWR VPWR _3810_/Y sky130_fd_sc_hd__nand2_1
X_4790_ _4784_/B _4675_/A _4759_/Y VGND VGND VPWR VPWR _5114_/A sky130_fd_sc_hd__o21ai_1
XFILLER_32_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_18 _3658_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_29 _3484_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3741_ _6930_/Q _5349_/A _4270_/A _6721_/Q VGND VGND VPWR VPWR _3741_/X sky130_fd_sc_hd__a22o_1
XFILLER_158_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6460_ _3945_/A1 _6460_/D _6415_/X VGND VGND VPWR VPWR _6460_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3672_ _6963_/Q _5385_/A _4240_/A _6687_/Q VGND VGND VPWR VPWR _3672_/X sky130_fd_sc_hd__a22o_1
XFILLER_173_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5411_ _5579_/A0 hold512/X _5411_/S VGND VGND VPWR VPWR _5411_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6391_ _6391_/A1 _6697_/Q _4232_/X _6390_/X VGND VGND VPWR VPWR _6391_/X sky130_fd_sc_hd__o31a_1
XFILLER_127_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5342_ _5573_/A0 hold924/X _5348_/S VGND VGND VPWR VPWR _5342_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_720 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5273_ _5567_/A0 hold661/X _5276_/S VGND VGND VPWR VPWR _5273_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7012_ _7012_/CLK _7012_/D fanout505/X VGND VGND VPWR VPWR _7012_/Q sky130_fd_sc_hd__dfrtp_2
X_4224_ _5459_/A0 hold87/X hold51/X VGND VGND VPWR VPWR hold88/A sky130_fd_sc_hd__mux2_1
X_4155_ _5459_/A0 hold367/X _4158_/S VGND VGND VPWR VPWR _4155_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4086_ hold973/X _4085_/X _4086_/S VGND VGND VPWR VPWR _4086_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4988_ _5090_/B _4988_/B _5170_/A _4988_/D VGND VGND VPWR VPWR _4989_/D sky130_fd_sc_hd__nor4_1
X_6727_ _6990_/CLK _6727_/D _3873_/A VGND VGND VPWR VPWR _6727_/Q sky130_fd_sc_hd__dfrtp_1
X_3939_ _7159_/Q _6815_/Q _6818_/Q VGND VGND VPWR VPWR _3939_/X sky130_fd_sc_hd__mux2_2
XFILLER_176_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6658_ _6709_/CLK _6658_/D _6441_/A VGND VGND VPWR VPWR _6658_/Q sky130_fd_sc_hd__dfrtp_1
X_5609_ _6562_/Q _6564_/Q VGND VGND VPWR VPWR _5609_/Y sky130_fd_sc_hd__nor2_1
XFILLER_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6589_ _6707_/CLK _6589_/D _6433_/A VGND VGND VPWR VPWR _6589_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput16 mask_rev_in[20] VGND VGND VPWR VPWR input16/X sky130_fd_sc_hd__clkbuf_2
Xinput27 mask_rev_in[30] VGND VGND VPWR VPWR input27/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput38 mgmt_gpio_in[11] VGND VGND VPWR VPWR input38/X sky130_fd_sc_hd__clkbuf_4
XFILLER_167_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput49 mgmt_gpio_in[21] VGND VGND VPWR VPWR input49/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_182_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5960_ _6715_/Q _5960_/B VGND VGND VPWR VPWR _5960_/X sky130_fd_sc_hd__or2_1
X_4911_ _5076_/B _5016_/A _4672_/A VGND VGND VPWR VPWR _4911_/X sky130_fd_sc_hd__a21o_1
X_5891_ _5891_/A _5891_/B _5891_/C _5891_/D VGND VGND VPWR VPWR _5891_/X sky130_fd_sc_hd__or4_1
XFILLER_61_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4842_ _4646_/A _4692_/B _4860_/A VGND VGND VPWR VPWR _4842_/Y sky130_fd_sc_hd__o21ai_1
X_4773_ _4570_/D _5042_/A _5042_/B _4772_/X _5158_/A VGND VGND VPWR VPWR _4773_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_20_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6512_ _7093_/CLK _6512_/D _6432_/A VGND VGND VPWR VPWR _6512_/Q sky130_fd_sc_hd__dfrtp_1
X_3724_ _3723_/X _6783_/Q _3791_/A VGND VGND VPWR VPWR _3724_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3655_ _6753_/Q _4306_/A _4034_/A _6528_/Q VGND VGND VPWR VPWR _3655_/X sky130_fd_sc_hd__a22o_1
X_6443_ _6443_/CLK _6443_/D _3873_/X VGND VGND VPWR VPWR _6443_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_106_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6374_ _6373_/X _6374_/A1 _6386_/S VGND VGND VPWR VPWR _7200_/D sky130_fd_sc_hd__mux2_1
X_3586_ _6534_/Q _4040_/A _6392_/A _7210_/Q _3553_/X VGND VGND VPWR VPWR _3588_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_161_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5325_ hold267/X hold44/X _5330_/S VGND VGND VPWR VPWR _5325_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5256_ hold621/X _5550_/A0 _5258_/S VGND VGND VPWR VPWR _5256_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4207_ _4207_/A0 _6395_/A0 _4209_/S VGND VGND VPWR VPWR _4207_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5187_ _5187_/A _6392_/B VGND VGND VPWR VPWR _5192_/S sky130_fd_sc_hd__nand2_2
XFILLER_96_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4138_ _4138_/A0 _6395_/A0 _4140_/S VGND VGND VPWR VPWR _4138_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4069_ hold229/X _4068_/X _4069_/S VGND VGND VPWR VPWR _4069_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_523 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold608 _5389_/X VGND VGND VPWR VPWR _6965_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3440_ _6999_/Q _3300_/Y hold22/A _6903_/Q _3439_/X VGND VGND VPWR VPWR _3446_/C
+ sky130_fd_sc_hd__a221o_1
Xhold619 _6989_/Q VGND VGND VPWR VPWR hold619/X sky130_fd_sc_hd__dlygate4sd3_1
X_3371_ _3371_/A _3371_/B _3371_/C _3371_/D VGND VGND VPWR VPWR _3372_/B sky130_fd_sc_hd__or4_1
XFILLER_112_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5110_ _5156_/C _5178_/B _5110_/C VGND VGND VPWR VPWR _5110_/X sky130_fd_sc_hd__or3_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6090_ _6908_/Q _6024_/C _6272_/B _7068_/Q VGND VGND VPWR VPWR _6090_/X sky130_fd_sc_hd__a22o_1
XFILLER_112_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _4999_/B _4838_/B _5158_/A _5039_/X _5040_/X VGND VGND VPWR VPWR _5044_/B
+ sky130_fd_sc_hd__a2111o_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1308 hold1308/A VGND VGND VPWR VPWR wb_dat_o[15] sky130_fd_sc_hd__buf_12
XFILLER_84_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1319 hold1405/X VGND VGND VPWR VPWR hold1319/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_wb_clk_i wb_clk_i VGND VGND VPWR VPWR clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_92_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6992_ _6992_/CLK _6992_/D fanout516/X VGND VGND VPWR VPWR _6992_/Q sky130_fd_sc_hd__dfrtp_4
X_5943_ _7210_/Q _5671_/X _5706_/X _7093_/Q VGND VGND VPWR VPWR _5943_/X sky130_fd_sc_hd__a22o_1
XFILLER_179_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5874_ _6611_/Q _5683_/X _5706_/X _7090_/Q _5873_/X VGND VGND VPWR VPWR _5879_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_178_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4825_ _5158_/B _4823_/X _4824_/Y _4549_/Y VGND VGND VPWR VPWR _4825_/X sky130_fd_sc_hd__o31a_1
XFILLER_166_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4756_ _4876_/A _4744_/X _4755_/X _4971_/B VGND VGND VPWR VPWR _4761_/B sky130_fd_sc_hd__o22a_1
XFILLER_119_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3707_ _6907_/Q _5322_/A _4306_/A _6752_/Q _3706_/X VGND VGND VPWR VPWR _3710_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4687_ _4739_/A _5013_/A VGND VGND VPWR VPWR _4822_/A sky130_fd_sc_hd__nor2_1
XFILLER_174_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6426_ _6426_/A _6441_/B VGND VGND VPWR VPWR _6426_/X sky130_fd_sc_hd__and2_1
X_3638_ _6768_/Q _4324_/A _4312_/A _6758_/Q VGND VGND VPWR VPWR _3638_/X sky130_fd_sc_hd__a22o_1
XFILLER_162_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3569_ _7138_/Q hold69/A _5544_/A _7106_/Q VGND VGND VPWR VPWR _3569_/X sky130_fd_sc_hd__a22o_1
X_6357_ _6357_/A _6358_/A VGND VGND VPWR VPWR _6357_/Y sky130_fd_sc_hd__nand2_1
X_5308_ hold36/X hold199/X _5312_/S VGND VGND VPWR VPWR _5308_/X sky130_fd_sc_hd__mux2_1
X_6288_ _6603_/Q _5980_/Y _6036_/X _6518_/Q _6287_/X VGND VGND VPWR VPWR _6291_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_48_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5239_ _5569_/A0 _5239_/A1 _5240_/S VGND VGND VPWR VPWR _5239_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold5 hold8/X VGND VGND VPWR VPWR hold9/A sky130_fd_sc_hd__buf_6
XFILLER_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4610_ _4610_/A _4666_/B VGND VGND VPWR VPWR _4653_/C sky130_fd_sc_hd__or2_2
XFILLER_175_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5590_ _5615_/A _6819_/Q _6565_/Q _3896_/X _5589_/X VGND VGND VPWR VPWR _7143_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_128_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4541_ _4935_/A _4553_/B VGND VGND VPWR VPWR _4780_/A sky130_fd_sc_hd__nand2_2
XFILLER_144_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold405 _6717_/Q VGND VGND VPWR VPWR hold405/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire380 _4846_/D VGND VGND VPWR VPWR _4838_/B sky130_fd_sc_hd__buf_2
XFILLER_190_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold416 _5528_/X VGND VGND VPWR VPWR _7089_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4472_ _4846_/A _4570_/D _4846_/B _4570_/B VGND VGND VPWR VPWR _5023_/B sky130_fd_sc_hd__or4bb_4
Xhold427 _7021_/Q VGND VGND VPWR VPWR hold427/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold438 _5548_/X VGND VGND VPWR VPWR _7106_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3423_ _6991_/Q _3298_/Y _3326_/Y _7031_/Q _3422_/X VGND VGND VPWR VPWR _3445_/B
+ sky130_fd_sc_hd__a221o_1
X_6211_ _6929_/Q _6027_/B wire394/X _6897_/Q _6210_/X VGND VGND VPWR VPWR _6217_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_116_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold449 _6941_/Q VGND VGND VPWR VPWR hold449/X sky130_fd_sc_hd__dlygate4sd3_1
X_7191_ _7193_/CLK _7191_/D VGND VGND VPWR VPWR _7191_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_144_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6142_ _6142_/A _6142_/B _6142_/C _6142_/D VGND VGND VPWR VPWR _6143_/C sky130_fd_sc_hd__or4_4
X_3354_ _7142_/Q hold69/A hold78/A _7049_/Q _3353_/X VGND VGND VPWR VPWR _3355_/D
+ sky130_fd_sc_hd__a221o_4
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6073_ _7004_/Q _6202_/B1 _6323_/B1 _7121_/Q VGND VGND VPWR VPWR _6073_/X sky130_fd_sc_hd__a22o_1
Xhold1105 _6528_/Q VGND VGND VPWR VPWR _4037_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3285_ _3313_/B _3299_/B VGND VGND VPWR VPWR _5241_/B sky130_fd_sc_hd__nand2_8
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1116 _4301_/X VGND VGND VPWR VPWR _6746_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _5024_/A _5027_/B VGND VGND VPWR VPWR _5155_/A sky130_fd_sc_hd__nor2_1
Xhold1127 _6852_/Q VGND VGND VPWR VPWR _5262_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1138 _5532_/X VGND VGND VPWR VPWR _7092_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1149 _6795_/Q VGND VGND VPWR VPWR _5190_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_81_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6975_ _7108_/CLK _6975_/D fanout523/X VGND VGND VPWR VPWR _6975_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5926_ _5926_/A0 _5925_/X _6319_/S VGND VGND VPWR VPWR _7172_/D sky130_fd_sc_hd__mux2_1
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5857_ _5857_/A _5857_/B _5857_/C _5857_/D VGND VGND VPWR VPWR _5857_/X sky130_fd_sc_hd__or4_1
XFILLER_139_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4808_ _4814_/A _4784_/A _4814_/B _4424_/Y _4981_/B VGND VGND VPWR VPWR _4809_/C
+ sky130_fd_sc_hd__o32a_1
XFILLER_186_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5788_ _7006_/Q _5664_/X _5688_/X _6862_/Q VGND VGND VPWR VPWR _5788_/X sky130_fd_sc_hd__a22o_1
X_4739_ _4739_/A _4739_/B VGND VGND VPWR VPWR _5042_/B sky130_fd_sc_hd__nor2_1
XFILLER_181_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6409_ _6433_/A _6440_/B VGND VGND VPWR VPWR _6409_/X sky130_fd_sc_hd__and2_1
XFILLER_135_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold950 _6635_/Q VGND VGND VPWR VPWR hold950/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold961 _4307_/X VGND VGND VPWR VPWR _6751_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold972 _5233_/X VGND VGND VPWR VPWR _6826_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold983 _7208_/Q VGND VGND VPWR VPWR hold983/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold994 _5559_/X VGND VGND VPWR VPWR _7116_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_50_csclk _6970_/CLK VGND VGND VPWR VPWR _7110_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_99_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_65_csclk _6970_/CLK VGND VGND VPWR VPWR _7068_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_47_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6760_ _6760_/CLK _6760_/D fanout490/X VGND VGND VPWR VPWR _6760_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3972_ _3972_/A0 _6395_/A0 _3982_/S VGND VGND VPWR VPWR _3972_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5711_ _7051_/Q _5699_/X _5706_/X _6499_/Q VGND VGND VPWR VPWR _5711_/X sky130_fd_sc_hd__a22o_1
XFILLER_149_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6691_ _7200_/CLK _6691_/D _6348_/B VGND VGND VPWR VPWR _6691_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_149_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5642_ _6033_/A _6039_/A _6040_/B VGND VGND VPWR VPWR _5642_/X sky130_fd_sc_hd__and3_4
XFILLER_176_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5573_ _5573_/A0 hold896/X _5579_/S VGND VGND VPWR VPWR _5573_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold202 _5471_/X VGND VGND VPWR VPWR _7038_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4524_ _4742_/A _4524_/B VGND VGND VPWR VPWR _4524_/Y sky130_fd_sc_hd__nand2_1
Xhold213 _7084_/Q VGND VGND VPWR VPWR hold213/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 _5284_/X VGND VGND VPWR VPWR _6872_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_18_csclk _6820_/CLK VGND VGND VPWR VPWR _6740_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold235 _6769_/Q VGND VGND VPWR VPWR hold235/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold246 _5442_/X VGND VGND VPWR VPWR _7012_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4455_ _4456_/A _4724_/B VGND VGND VPWR VPWR _4524_/B sky130_fd_sc_hd__nor2_2
Xhold257 _6488_/Q VGND VGND VPWR VPWR hold257/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold268 _5325_/X VGND VGND VPWR VPWR _6908_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold279 _6997_/Q VGND VGND VPWR VPWR hold279/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3406_ input27/X _3340_/Y _5544_/A _7109_/Q VGND VGND VPWR VPWR _3406_/X sky130_fd_sc_hd__a22o_1
X_7174_ _7182_/CLK _7174_/D fanout499/X VGND VGND VPWR VPWR _7174_/Q sky130_fd_sc_hd__dfrtp_1
X_4386_ _4667_/C _5035_/A VGND VGND VPWR VPWR _4759_/A sky130_fd_sc_hd__nor2_8
XFILLER_131_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3337_ hold95/X _4120_/B VGND VGND VPWR VPWR _4083_/S sky130_fd_sc_hd__nor2_8
X_6125_ _7086_/Q _5977_/X _6323_/B1 _7123_/Q VGND VGND VPWR VPWR _6125_/X sky130_fd_sc_hd__a22o_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3268_ _5212_/A hold57/A VGND VGND VPWR VPWR _3268_/Y sky130_fd_sc_hd__nor2_8
XFILLER_86_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6056_ _6955_/Q _6336_/A2 _6205_/B1 _7059_/Q VGND VGND VPWR VPWR _6056_/X sky130_fd_sc_hd__a22o_1
XFILLER_65_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5007_ _5039_/A _5007_/B _5039_/B _5007_/D VGND VGND VPWR VPWR _5008_/D sky130_fd_sc_hd__or4_1
XFILLER_54_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3199_ _7122_/Q VGND VGND VPWR VPWR _3199_/Y sky130_fd_sc_hd__clkinv_2
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_108 _3949_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_119 _3949_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6958_ _7082_/CLK _6958_/D _3873_/A VGND VGND VPWR VPWR _6958_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_53_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5909_ _6613_/Q _5683_/X _5693_/X _6657_/Q VGND VGND VPWR VPWR _5909_/X sky130_fd_sc_hd__a22o_1
X_6889_ _6992_/CLK _6889_/D fanout517/X VGND VGND VPWR VPWR _6889_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_139_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold780 _5438_/X VGND VGND VPWR VPWR _7009_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold791 _7093_/Q VGND VGND VPWR VPWR hold791/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1480 _6645_/Q VGND VGND VPWR VPWR _4187_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1491 _6644_/Q VGND VGND VPWR VPWR _4186_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput307 _5592_/B VGND VGND VPWR VPWR serial_clock sky130_fd_sc_hd__buf_12
Xoutput318 hold1345/X VGND VGND VPWR VPWR hold1346/A sky130_fd_sc_hd__buf_12
Xoutput329 hold1347/X VGND VGND VPWR VPWR hold1348/A sky130_fd_sc_hd__buf_12
XFILLER_141_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4240_ _4240_/A _4330_/B VGND VGND VPWR VPWR _4245_/S sky130_fd_sc_hd__and2_2
XFILLER_113_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4171_ _4171_/A0 _3447_/X _4173_/S VGND VGND VPWR VPWR _6631_/D sky130_fd_sc_hd__mux2_1
XFILLER_122_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6812_ _6986_/CLK _6812_/D fanout491/X VGND VGND VPWR VPWR _6812_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_51_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6743_ _7207_/CLK _6743_/D fanout484/X VGND VGND VPWR VPWR _6743_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_189_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3955_ _6696_/Q _3962_/B VGND VGND VPWR VPWR _6694_/D sky130_fd_sc_hd__and2_1
XFILLER_188_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6674_ _7094_/CLK _6674_/D fanout496/X VGND VGND VPWR VPWR _6674_/Q sky130_fd_sc_hd__dfrtp_2
X_3886_ _4467_/A _4654_/B _3886_/C _3886_/D VGND VGND VPWR VPWR _3887_/D sky130_fd_sc_hd__or4_1
X_5625_ _5624_/Y _5960_/B _5625_/S VGND VGND VPWR VPWR _7152_/D sky130_fd_sc_hd__mux2_1
XFILLER_137_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5556_ _5574_/A0 _5556_/A1 _5561_/S VGND VGND VPWR VPWR _5556_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4507_ _4738_/A _4942_/A _4996_/A VGND VGND VPWR VPWR _4507_/X sky130_fd_sc_hd__a21o_1
X_5487_ _5574_/A0 _5487_/A1 _5492_/S VGND VGND VPWR VPWR _5487_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4438_ _4453_/C _4456_/A VGND VGND VPWR VPWR _4448_/B sky130_fd_sc_hd__nor2_1
Xfanout501 fanout508/X VGND VGND VPWR VPWR fanout501/X sky130_fd_sc_hd__buf_8
Xfanout512 fanout527/X VGND VGND VPWR VPWR _3873_/A sky130_fd_sc_hd__buf_8
XFILLER_132_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout523 fanout526/X VGND VGND VPWR VPWR fanout523/X sky130_fd_sc_hd__buf_6
X_7157_ _7181_/CLK _7157_/D fanout502/X VGND VGND VPWR VPWR _7157_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_116_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4369_ _4596_/A _4369_/B VGND VGND VPWR VPWR _5076_/A sky130_fd_sc_hd__or2_4
XFILLER_112_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6108_ _7013_/Q _5998_/Y _6049_/B _7029_/Q _6107_/X VGND VGND VPWR VPWR _6109_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_59_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7088_ _7088_/CLK _7088_/D fanout507/X VGND VGND VPWR VPWR _7088_/Q sky130_fd_sc_hd__dfrtp_2
X_6039_ _6039_/A _6040_/B _6039_/C VGND VGND VPWR VPWR _6272_/B sky130_fd_sc_hd__and3_4
XFILLER_27_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_19 _3410_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3740_ _6898_/Q hold22/A _4276_/A _6726_/Q VGND VGND VPWR VPWR _3740_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3671_ _7096_/Q _5535_/A _4046_/A _6537_/Q _3670_/X VGND VGND VPWR VPWR _3679_/A
+ sky130_fd_sc_hd__a221o_1
X_5410_ _5587_/A0 hold900/X _5411_/S VGND VGND VPWR VPWR _5410_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6390_ _3191_/Y _6390_/A2 _6360_/X _6389_/X _6358_/A VGND VGND VPWR VPWR _6390_/X
+ sky130_fd_sc_hd__a32o_1
X_5341_ _5536_/A1 _5341_/A1 _5348_/S VGND VGND VPWR VPWR _5341_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5272_ _5539_/A1 hold161/X _5276_/S VGND VGND VPWR VPWR _5272_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7011_ _7075_/CLK _7011_/D fanout514/X VGND VGND VPWR VPWR _7011_/Q sky130_fd_sc_hd__dfstp_1
X_4223_ _5521_/A0 hold944/X hold51/X VGND VGND VPWR VPWR _4223_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4154_ _5521_/A0 _4154_/A1 _4158_/S VGND VGND VPWR VPWR _4154_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4085_ hold755/X _5552_/A0 _4085_/S VGND VGND VPWR VPWR _4085_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4987_ _4987_/A _4987_/B _4987_/C VGND VGND VPWR VPWR _4988_/D sky130_fd_sc_hd__or3_1
X_6726_ _6990_/CLK _6726_/D _3873_/A VGND VGND VPWR VPWR _6726_/Q sky130_fd_sc_hd__dfrtp_1
X_3938_ _6571_/Q input93/X _6823_/Q VGND VGND VPWR VPWR _3938_/X sky130_fd_sc_hd__mux2_2
XFILLER_177_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6657_ _6708_/CLK _6657_/D _6432_/A VGND VGND VPWR VPWR _6657_/Q sky130_fd_sc_hd__dfstp_1
X_3869_ _3184_/Y input58/X _3868_/B _3868_/Y VGND VGND VPWR VPWR _6445_/D sky130_fd_sc_hd__a31o_1
XFILLER_164_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5608_ _5608_/A1 _5605_/A _5607_/Y VGND VGND VPWR VPWR _7147_/D sky130_fd_sc_hd__o21a_1
XFILLER_137_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6588_ _6664_/CLK _6588_/D _6426_/A VGND VGND VPWR VPWR _6588_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_117_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5539_ hold207/X _5539_/A1 _5543_/S VGND VGND VPWR VPWR _5539_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7209_ _7209_/CLK _7209_/D fanout485/X VGND VGND VPWR VPWR _7209_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_160_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput17 mask_rev_in[21] VGND VGND VPWR VPWR input17/X sky130_fd_sc_hd__clkbuf_1
XFILLER_168_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput28 mask_rev_in[31] VGND VGND VPWR VPWR input28/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput39 mgmt_gpio_in[12] VGND VGND VPWR VPWR _3961_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_182_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4910_ _4683_/A _4646_/A _4707_/B VGND VGND VPWR VPWR _4910_/X sky130_fd_sc_hd__a21o_1
XFILLER_45_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5890_ _6687_/Q _5666_/X _5699_/X _6537_/Q _5889_/X VGND VGND VPWR VPWR _5891_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_61_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4841_ _5023_/B _4677_/B _4520_/X VGND VGND VPWR VPWR _5162_/B sky130_fd_sc_hd__o21ai_1
XFILLER_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4772_ _4657_/C _5060_/A _4770_/X _4771_/X VGND VGND VPWR VPWR _4772_/X sky130_fd_sc_hd__a211o_1
XFILLER_159_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6511_ _7093_/CLK _6511_/D _6432_/A VGND VGND VPWR VPWR _6511_/Q sky130_fd_sc_hd__dfrtp_2
X_3723_ _3723_/A _3723_/B _3723_/C VGND VGND VPWR VPWR _3723_/X sky130_fd_sc_hd__or3_4
XFILLER_119_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6442_ _3945_/A1 _6442_/D _6398_/X VGND VGND VPWR VPWR hold11/A sky130_fd_sc_hd__dfrtn_1
XFILLER_146_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3654_ _7084_/Q _5520_/A _3684_/B1 _7052_/Q _3605_/X VGND VGND VPWR VPWR _3659_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6373_ _6700_/Q _6373_/A2 _6373_/B1 _6390_/A2 _6372_/X VGND VGND VPWR VPWR _6373_/X
+ sky130_fd_sc_hd__a221o_1
Xclkbuf_3_0_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A VGND VGND VPWR VPWR _7183_/CLK sky130_fd_sc_hd__clkbuf_8
X_3585_ _6801_/Q _5193_/A _3547_/Y input95/X _3552_/X VGND VGND VPWR VPWR _3588_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_161_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5324_ hold339/X _5459_/A0 _5330_/S VGND VGND VPWR VPWR _5324_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5255_ hold156/X _5558_/A0 _5258_/S VGND VGND VPWR VPWR _5255_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4206_ _4206_/A0 _6394_/A0 _4209_/S VGND VGND VPWR VPWR _4206_/X sky130_fd_sc_hd__mux2_1
X_5186_ _6394_/A0 _5186_/A1 _5186_/S VGND VGND VPWR VPWR _5186_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4137_ _4137_/A0 _6394_/A0 _4140_/S VGND VGND VPWR VPWR _4137_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4068_ _4119_/A1 hold40/X _4068_/S VGND VGND VPWR VPWR _4068_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6709_ _6709_/CLK _6709_/D fanout496/X VGND VGND VPWR VPWR _6709_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_177_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold609 _7039_/Q VGND VGND VPWR VPWR hold609/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3370_ _6977_/Q _5394_/A _5277_/A _6873_/Q _3369_/X VGND VGND VPWR VPWR _3371_/D
+ sky130_fd_sc_hd__a221o_1
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _4999_/B _5060_/A _5130_/A VGND VGND VPWR VPWR _5040_/X sky130_fd_sc_hd__a21o_1
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1309 hold1398/X VGND VGND VPWR VPWR hold1309/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6991_ _7065_/CLK _6991_/D fanout517/X VGND VGND VPWR VPWR _6991_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5942_ _6689_/Q _5666_/X _5682_/X _6514_/Q _5941_/X VGND VGND VPWR VPWR _5945_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_18_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5873_ _6741_/Q _5656_/X _5689_/X _5872_/X VGND VGND VPWR VPWR _5873_/X sky130_fd_sc_hd__a22o_1
XFILLER_61_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4824_ _4824_/A _4992_/B VGND VGND VPWR VPWR _4824_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4755_ _4759_/A _4758_/A _5001_/A _4758_/B _4993_/A VGND VGND VPWR VPWR _4755_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_159_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3706_ _6818_/Q _5221_/B _4016_/A _6512_/Q VGND VGND VPWR VPWR _3706_/X sky130_fd_sc_hd__a22o_1
XFILLER_119_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4686_ _5013_/A _5021_/B VGND VGND VPWR VPWR _4882_/B sky130_fd_sc_hd__or2_1
XFILLER_174_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6425_ _6441_/A _6440_/B VGND VGND VPWR VPWR _6425_/X sky130_fd_sc_hd__and2_1
XFILLER_119_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3637_ input5/X _3295_/Y _3992_/A _6492_/Q _3636_/X VGND VGND VPWR VPWR _3642_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6356_ _6356_/A0 _3373_/X _6356_/S VGND VGND VPWR VPWR _7196_/D sky130_fd_sc_hd__mux2_1
X_3568_ _6949_/Q _5367_/A _5205_/A _6810_/Q _3567_/X VGND VGND VPWR VPWR _3573_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_88_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5307_ _5496_/A0 hold854/X _5312_/S VGND VGND VPWR VPWR _5307_/X sky130_fd_sc_hd__mux2_1
X_6287_ _7092_/Q _5642_/X _5992_/X _6677_/Q VGND VGND VPWR VPWR _6287_/X sky130_fd_sc_hd__a22o_1
XFILLER_88_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3499_ _3499_/A _3499_/B _3499_/C _3499_/D VGND VGND VPWR VPWR _3542_/A sky130_fd_sc_hd__or4_2
X_5238_ _5550_/A0 hold411/X _5240_/S VGND VGND VPWR VPWR _5238_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5169_ _4683_/A _4784_/B _4728_/Y _5003_/A _4626_/Y VGND VGND VPWR VPWR _5169_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_56_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold6 hold6/A VGND VGND VPWR VPWR hold6/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_59_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4540_ _4935_/A _4819_/C _4971_/B VGND VGND VPWR VPWR _4792_/A sky130_fd_sc_hd__and3_1
XFILLER_129_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold406 _4266_/X VGND VGND VPWR VPWR _6717_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4471_ _4570_/D _4471_/B VGND VGND VPWR VPWR _4475_/A sky130_fd_sc_hd__nor2_1
XFILLER_183_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold417 _6558_/Q VGND VGND VPWR VPWR hold417/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold428 _5452_/X VGND VGND VPWR VPWR _7021_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6210_ _6921_/Q wire412/X _6024_/D _6945_/Q VGND VGND VPWR VPWR _6210_/X sky130_fd_sc_hd__a22o_1
XFILLER_116_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold439 _7085_/Q VGND VGND VPWR VPWR hold439/X sky130_fd_sc_hd__dlygate4sd3_1
X_3422_ input31/X _3304_/Y _3983_/A _6487_/Q VGND VGND VPWR VPWR _3422_/X sky130_fd_sc_hd__a22o_2
X_7190_ _7193_/CLK _7190_/D VGND VGND VPWR VPWR _7190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6141_ _6854_/Q _6027_/A _6329_/B1 _7038_/Q _6140_/X VGND VGND VPWR VPWR _6142_/D
+ sky130_fd_sc_hd__a221o_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ _7073_/Q _5502_/A _5562_/A _7126_/Q VGND VGND VPWR VPWR _3353_/X sky130_fd_sc_hd__a22o_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6072_ _6072_/A0 _6071_/X _6319_/S VGND VGND VPWR VPWR _7176_/D sky130_fd_sc_hd__mux2_1
XFILLER_112_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3284_ hold55/X hold27/X VGND VGND VPWR VPWR _3330_/B sky130_fd_sc_hd__nor2_8
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1106 _4037_/X VGND VGND VPWR VPWR _6528_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1117 _6742_/Q VGND VGND VPWR VPWR _4296_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5023_ _5023_/A _5023_/B _5023_/C VGND VGND VPWR VPWR _5027_/B sky130_fd_sc_hd__and3_2
Xhold1128 _5262_/X VGND VGND VPWR VPWR _6852_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1139 _6612_/Q VGND VGND VPWR VPWR _4149_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6974_ _7139_/CLK _6974_/D fanout518/X VGND VGND VPWR VPWR _6974_/Q sky130_fd_sc_hd__dfrtp_4
X_5925_ _6563_/Q _7171_/Q _5924_/X VGND VGND VPWR VPWR _5925_/X sky130_fd_sc_hd__a21o_1
XFILLER_61_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5856_ _6921_/Q _5677_/X _5699_/X _7057_/Q _5855_/X VGND VGND VPWR VPWR _5857_/D
+ sky130_fd_sc_hd__a221o_1
X_4807_ _4794_/A _4569_/B _4653_/C _5094_/B _4802_/A VGND VGND VPWR VPWR _4809_/B
+ sky130_fd_sc_hd__o32a_1
X_5787_ _6894_/Q _5655_/X _5775_/X _5786_/X VGND VGND VPWR VPWR _5792_/A sky130_fd_sc_hd__a211o_1
XFILLER_166_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4738_ _4738_/A _4739_/B VGND VGND VPWR VPWR _5042_/A sky130_fd_sc_hd__nor2_1
XFILLER_119_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4669_ _4663_/Y _4666_/Y _4667_/X _4665_/Y _4674_/A VGND VGND VPWR VPWR _4669_/X
+ sky130_fd_sc_hd__o32a_1
X_6408_ _6433_/A _6440_/B VGND VGND VPWR VPWR _6408_/X sky130_fd_sc_hd__and2_1
Xhold940 _6522_/Q VGND VGND VPWR VPWR hold940/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold951 _4176_/X VGND VGND VPWR VPWR _6635_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold962 _6812_/Q VGND VGND VPWR VPWR hold962/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold973 _6561_/Q VGND VGND VPWR VPWR hold973/X sky130_fd_sc_hd__dlygate4sd3_1
X_6339_ _6760_/Q _6007_/Y _6040_/X _6530_/Q _6338_/X VGND VGND VPWR VPWR _6339_/X
+ sky130_fd_sc_hd__a221o_2
Xhold984 _6394_/X VGND VGND VPWR VPWR _7208_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold995 _6911_/Q VGND VGND VPWR VPWR hold995/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3971_ hold42/X hold61/X _3971_/S VGND VGND VPWR VPWR hold62/A sky130_fd_sc_hd__mux2_4
X_5710_ _5710_/A1 _5652_/Y _5709_/X VGND VGND VPWR VPWR _7162_/D sky130_fd_sc_hd__a21o_1
XFILLER_43_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6690_ _7094_/CLK _6690_/D fanout496/X VGND VGND VPWR VPWR _6690_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5641_ _7158_/Q _7157_/Q VGND VGND VPWR VPWR _6038_/A sky130_fd_sc_hd__nand2b_4
XFILLER_148_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5572_ _5581_/A0 _5572_/A1 _5579_/S VGND VGND VPWR VPWR _5572_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_1_csclk clkbuf_1_0_1_csclk/A VGND VGND VPWR VPWR clkbuf_2_1_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_163_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4523_ _4997_/A _5035_/B VGND VGND VPWR VPWR _5049_/A sky130_fd_sc_hd__nor2_2
XFILLER_129_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold203 _6827_/Q VGND VGND VPWR VPWR hold203/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 _5523_/X VGND VGND VPWR VPWR _7084_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold225 _6748_/Q VGND VGND VPWR VPWR hold225/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 _4328_/X VGND VGND VPWR VPWR _6769_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4454_ _5002_/A VGND VGND VPWR VPWR _4454_/Y sky130_fd_sc_hd__inv_2
Xhold247 _6980_/Q VGND VGND VPWR VPWR hold247/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 _3990_/X VGND VGND VPWR VPWR _6488_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold269 _6992_/Q VGND VGND VPWR VPWR hold269/X sky130_fd_sc_hd__dlygate4sd3_1
X_3405_ _7133_/Q _5571_/A _4085_/S input69/X _3384_/X VGND VGND VPWR VPWR _3408_/C
+ sky130_fd_sc_hd__a221o_1
X_7173_ _7187_/CLK _7173_/D fanout488/X VGND VGND VPWR VPWR _7173_/Q sky130_fd_sc_hd__dfrtp_1
X_4385_ _4570_/D _4385_/B VGND VGND VPWR VPWR _5035_/A sky130_fd_sc_hd__or2_4
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6124_ _7054_/Q _5988_/X _6199_/B1 _6870_/Q VGND VGND VPWR VPWR _6124_/X sky130_fd_sc_hd__a22o_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3336_ hold95/X _3340_/B VGND VGND VPWR VPWR _5562_/A sky130_fd_sc_hd__nor2_8
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0__1134_ _3543_/X VGND VGND VPWR VPWR clkbuf_0__1134_/X sky130_fd_sc_hd__clkbuf_16
X_6055_ _7019_/Q _6204_/A2 _6025_/B _7104_/Q _6054_/X VGND VGND VPWR VPWR _6058_/C
+ sky130_fd_sc_hd__a221o_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3267_ _3299_/A hold56/X VGND VGND VPWR VPWR hold57/A sky130_fd_sc_hd__nand2_8
XFILLER_100_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5006_ _4876_/A _4485_/A _4744_/X _4993_/B _4993_/A VGND VGND VPWR VPWR _5007_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_38_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3198_ _7130_/Q VGND VGND VPWR VPWR _3198_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_54_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_109 _3949_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6957_ _7140_/CLK _6957_/D fanout522/X VGND VGND VPWR VPWR _6957_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_81_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5908_ _6513_/Q _5682_/X _5685_/X _6662_/Q _5907_/X VGND VGND VPWR VPWR _5913_/B
+ sky130_fd_sc_hd__a221o_1
X_6888_ _6977_/CLK _6888_/D fanout507/X VGND VGND VPWR VPWR _6888_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_139_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5839_ _7073_/Q _5678_/X _5686_/X _7017_/Q VGND VGND VPWR VPWR _5839_/X sky130_fd_sc_hd__a22o_1
XFILLER_10_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold770 _5318_/X VGND VGND VPWR VPWR _6902_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold781 _6993_/Q VGND VGND VPWR VPWR hold781/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold792 _5533_/X VGND VGND VPWR VPWR _7093_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3234__1 net499_2/A VGND VGND VPWR VPWR _6443_/CLK sky130_fd_sc_hd__inv_2
XFILLER_162_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1470 _6692_/Q VGND VGND VPWR VPWR _6697_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1481 _6629_/Q VGND VGND VPWR VPWR _4169_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1492 _6695_/Q VGND VGND VPWR VPWR _3894_/B1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_644 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput308 _3413_/X VGND VGND VPWR VPWR serial_data_1 sky130_fd_sc_hd__buf_12
Xoutput319 hold1323/X VGND VGND VPWR VPWR hold1324/A sky130_fd_sc_hd__buf_12
XFILLER_4_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4170_ _4170_/A0 _4185_/A1 _4173_/S VGND VGND VPWR VPWR _6630_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6811_ _7209_/CLK _6811_/D _3946_/B VGND VGND VPWR VPWR _6811_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_36_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6742_ _7207_/CLK _6742_/D fanout484/X VGND VGND VPWR VPWR _6742_/Q sky130_fd_sc_hd__dfrtp_4
X_3954_ _6698_/Q _3962_/B VGND VGND VPWR VPWR _6695_/D sky130_fd_sc_hd__and2_1
XFILLER_149_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6673_ _7094_/CLK _6673_/D fanout496/X VGND VGND VPWR VPWR _6673_/Q sky130_fd_sc_hd__dfrtp_1
X_3885_ _3885_/A _3885_/B input120/X input117/X VGND VGND VPWR VPWR _3886_/D sky130_fd_sc_hd__or4bb_1
XFILLER_176_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5624_ _5960_/B _5624_/B VGND VGND VPWR VPWR _5624_/Y sky130_fd_sc_hd__nand2_1
XFILLER_176_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5555_ _5555_/A0 hold373/X _5561_/S VGND VGND VPWR VPWR _5555_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4506_ _4996_/A _5035_/B VGND VGND VPWR VPWR _4506_/Y sky130_fd_sc_hd__nor2_2
X_5486_ _5573_/A0 hold795/X _5492_/S VGND VGND VPWR VPWR _5486_/X sky130_fd_sc_hd__mux2_1
XFILLER_104_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4437_ _4758_/A _4744_/C VGND VGND VPWR VPWR _4456_/A sky130_fd_sc_hd__nand2_1
XFILLER_104_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout502 fanout504/X VGND VGND VPWR VPWR fanout502/X sky130_fd_sc_hd__buf_8
XFILLER_132_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout513 fanout527/X VGND VGND VPWR VPWR _6407_/A sky130_fd_sc_hd__buf_6
X_7156_ _7182_/CLK _7156_/D fanout502/X VGND VGND VPWR VPWR _7156_/Q sky130_fd_sc_hd__dfrtp_1
Xfanout524 fanout525/X VGND VGND VPWR VPWR fanout524/X sky130_fd_sc_hd__buf_8
X_4368_ _4596_/A _4369_/B VGND VGND VPWR VPWR _4931_/A sky130_fd_sc_hd__nor2_2
XFILLER_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6107_ _7077_/Q _5994_/X _6204_/A2 _7021_/Q VGND VGND VPWR VPWR _6107_/X sky130_fd_sc_hd__a22o_1
XFILLER_59_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3319_ _3528_/A _3340_/B VGND VGND VPWR VPWR _5277_/A sky130_fd_sc_hd__nor2_8
X_7087_ _7126_/CLK _7087_/D fanout524/X VGND VGND VPWR VPWR _7087_/Q sky130_fd_sc_hd__dfrtp_2
X_4299_ _6397_/A0 hold480/X _4299_/S VGND VGND VPWR VPWR _4299_/X sky130_fd_sc_hd__mux2_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6038_ _6038_/A _6038_/B VGND VGND VPWR VPWR _6038_/Y sky130_fd_sc_hd__nor2_8
XFILLER_100_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_64_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7137_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_41_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_17_csclk _6882_/CLK VGND VGND VPWR VPWR _6990_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3670_ _6597_/Q _4129_/A _4312_/A _6757_/Q VGND VGND VPWR VPWR _3670_/X sky130_fd_sc_hd__a22o_1
XFILLER_185_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5340_ _5340_/A _5535_/B VGND VGND VPWR VPWR _5348_/S sky130_fd_sc_hd__nand2_8
XFILLER_127_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5271_ _5574_/A0 _5271_/A1 _5276_/S VGND VGND VPWR VPWR _5271_/X sky130_fd_sc_hd__mux2_1
XFILLER_181_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7010_ _7043_/CLK _7010_/D fanout514/X VGND VGND VPWR VPWR _7010_/Q sky130_fd_sc_hd__dfstp_2
X_4222_ hold50/X _5580_/B VGND VGND VPWR VPWR hold51/A sky130_fd_sc_hd__nand2_2
XFILLER_68_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4153_ _4153_/A _5580_/B VGND VGND VPWR VPWR _4158_/S sky130_fd_sc_hd__nand2_2
XFILLER_55_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4084_ hold409/X _4083_/X _4086_/S VGND VGND VPWR VPWR _4084_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4986_ _4986_/A _4986_/B _4799_/X VGND VGND VPWR VPWR _5170_/A sky130_fd_sc_hd__or3b_1
X_6725_ _6725_/CLK _6725_/D fanout510/X VGND VGND VPWR VPWR _6725_/Q sky130_fd_sc_hd__dfrtp_2
X_3937_ _6572_/Q _3937_/A1 _6821_/Q VGND VGND VPWR VPWR _3937_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6656_ _6707_/CLK _6656_/D _6432_/A VGND VGND VPWR VPWR _6656_/Q sky130_fd_sc_hd__dfrtp_4
X_3868_ _3868_/A _3868_/B VGND VGND VPWR VPWR _3868_/Y sky130_fd_sc_hd__nor2_1
XFILLER_137_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5607_ _7147_/Q _5605_/A _5606_/A VGND VGND VPWR VPWR _5607_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_191_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6587_ _7136_/CLK hold41/X fanout520/X VGND VGND VPWR VPWR _6587_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_191_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3799_ _6471_/Q _3801_/B _6472_/Q VGND VGND VPWR VPWR _3800_/B sky130_fd_sc_hd__a21oi_1
XFILLER_152_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5538_ hold265/X _5583_/A0 _5543_/S VGND VGND VPWR VPWR _5538_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5469_ hold313/X _5583_/A0 _5474_/S VGND VGND VPWR VPWR _5469_/X sky130_fd_sc_hd__mux2_1
X_7208_ _7211_/CLK _7208_/D fanout485/X VGND VGND VPWR VPWR _7208_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_132_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7139_ _7139_/CLK _7139_/D fanout518/X VGND VGND VPWR VPWR _7139_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_86_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput18 mask_rev_in[22] VGND VGND VPWR VPWR input18/X sky130_fd_sc_hd__clkbuf_2
XFILLER_183_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput29 mask_rev_in[3] VGND VGND VPWR VPWR input29/X sky130_fd_sc_hd__clkbuf_1
XFILLER_109_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4840_ _5023_/B _4659_/B _4447_/Y VGND VGND VPWR VPWR _5065_/C sky130_fd_sc_hd__o21ai_1
XTAP_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4771_ _4657_/C _4838_/B _4670_/Y VGND VGND VPWR VPWR _4771_/X sky130_fd_sc_hd__a21o_1
XFILLER_14_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6510_ _6709_/CLK _6510_/D _6441_/A VGND VGND VPWR VPWR _6510_/Q sky130_fd_sc_hd__dfrtp_2
X_3722_ _3722_/A _3722_/B _3722_/C _3722_/D VGND VGND VPWR VPWR _3723_/C sky130_fd_sc_hd__or4_1
XFILLER_119_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6441_ _6441_/A _6441_/B VGND VGND VPWR VPWR _6441_/X sky130_fd_sc_hd__and2_1
XFILLER_158_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3653_ _6996_/Q _3300_/Y _5430_/A _7004_/Q _3652_/X VGND VGND VPWR VPWR _3659_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6372_ _6698_/Q _6372_/A2 _6372_/B1 _6699_/Q VGND VGND VPWR VPWR _6372_/X sky130_fd_sc_hd__a22o_1
X_3584_ _7021_/Q _5448_/A _3340_/Y input23/X _3559_/X VGND VGND VPWR VPWR _3588_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5323_ _5323_/A0 _5521_/A0 _5330_/S VGND VGND VPWR VPWR _5323_/X sky130_fd_sc_hd__mux2_1
X_5254_ hold205/X _5539_/A1 _5258_/S VGND VGND VPWR VPWR _5254_/X sky130_fd_sc_hd__mux2_1
X_4205_ _4205_/A0 _6393_/A0 _4209_/S VGND VGND VPWR VPWR _4205_/X sky130_fd_sc_hd__mux2_1
X_5185_ _6393_/A0 _5185_/A1 _5186_/S VGND VGND VPWR VPWR _5185_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_3_6_0_csclk clkbuf_3_7_0_csclk/A VGND VGND VPWR VPWR _6931_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4136_ _4136_/A0 _6393_/A0 _4140_/S VGND VGND VPWR VPWR _4136_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4067_ hold421/X _4066_/X _4069_/S VGND VGND VPWR VPWR _4067_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4969_ _4969_/A _4969_/B VGND VGND VPWR VPWR _5114_/B sky130_fd_sc_hd__nand2_1
XFILLER_149_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6708_ _6708_/CLK _6708_/D fanout494/X VGND VGND VPWR VPWR _6708_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_20_661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6639_ _7193_/CLK _6639_/D VGND VGND VPWR VPWR _6639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6990_ _6990_/CLK _6990_/D _3873_/A VGND VGND VPWR VPWR _6990_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_53_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5941_ _6673_/Q _5955_/A2 _5705_/X _6684_/Q VGND VGND VPWR VPWR _5941_/X sky130_fd_sc_hd__a22o_1
XFILLER_18_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5872_ _6711_/Q _5938_/B VGND VGND VPWR VPWR _5872_/X sky130_fd_sc_hd__or2_1
XFILLER_34_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4823_ _5148_/A _5158_/A _4823_/C _4778_/Y VGND VGND VPWR VPWR _4823_/X sky130_fd_sc_hd__or4b_1
XFILLER_166_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4754_ _4995_/A _5036_/A VGND VGND VPWR VPWR _4984_/B sky130_fd_sc_hd__nor2_1
XFILLER_193_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3705_ _7091_/Q _5529_/A _4288_/A _6737_/Q _3704_/X VGND VGND VPWR VPWR _3710_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_119_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4685_ _5013_/A _4814_/B _5128_/B VGND VGND VPWR VPWR _4714_/A sky130_fd_sc_hd__o21ai_1
XFILLER_134_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3636_ input22/X _3340_/Y _4294_/A _6743_/Q VGND VGND VPWR VPWR _3636_/X sky130_fd_sc_hd__a22o_1
X_6424_ _6441_/A _6441_/B VGND VGND VPWR VPWR _6424_/X sky130_fd_sc_hd__and2_1
XFILLER_146_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6355_ _6355_/A0 _3410_/X _6356_/S VGND VGND VPWR VPWR _7195_/D sky130_fd_sc_hd__mux2_1
X_3567_ _6689_/Q _4240_/A _4216_/A _6673_/Q VGND VGND VPWR VPWR _3567_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5306_ _5555_/A0 hold345/X _5312_/S VGND VGND VPWR VPWR _5306_/X sky130_fd_sc_hd__mux2_1
X_6286_ _6608_/Q _6326_/A2 _6021_/Y _6623_/Q _6285_/X VGND VGND VPWR VPWR _6291_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3498_ _7046_/Q hold77/A _4028_/A _6525_/Q _3497_/X VGND VGND VPWR VPWR _3499_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_88_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5237_ hold85/X _5237_/A1 _5240_/S VGND VGND VPWR VPWR _5237_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5168_ _5168_/A1 _6362_/A _5157_/X _5167_/X VGND VGND VPWR VPWR _6781_/D sky130_fd_sc_hd__a211o_1
XFILLER_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4119_ hold40/X _4119_/A1 hold97/X VGND VGND VPWR VPWR hold41/A sky130_fd_sc_hd__mux2_1
XFILLER_83_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5099_ _4657_/A _4732_/A _4759_/A _4607_/X _4829_/Y VGND VGND VPWR VPWR _5100_/D
+ sky130_fd_sc_hd__a311o_1
XFILLER_56_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold7 hold7/A VGND VGND VPWR VPWR hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_87_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire360 _6217_/A VGND VGND VPWR VPWR _6044_/A sky130_fd_sc_hd__clkbuf_2
X_4470_ _4512_/B _4657_/C VGND VGND VPWR VPWR _4510_/B sky130_fd_sc_hd__nand2_1
Xhold407 _6995_/Q VGND VGND VPWR VPWR hold407/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold418 _4080_/X VGND VGND VPWR VPWR _6558_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3421_ _7100_/Q _5535_/A hold78/A _7047_/Q _3420_/X VGND VGND VPWR VPWR _3445_/A
+ sky130_fd_sc_hd__a221o_2
Xhold429 _7013_/Q VGND VGND VPWR VPWR hold429/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6140_ _6502_/Q _6323_/A2 _6024_/B _6934_/Q VGND VGND VPWR VPWR _6140_/X sky130_fd_sc_hd__a22o_1
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3352_ input60/X _5232_/A _5571_/A _7134_/Q _3351_/X VGND VGND VPWR VPWR _3355_/C
+ sky130_fd_sc_hd__a221o_4
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6071_ _5650_/A _6071_/A2 _6070_/X VGND VGND VPWR VPWR _6071_/X sky130_fd_sc_hd__a21o_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3283_ _3283_/A VGND VGND VPWR VPWR _3313_/B sky130_fd_sc_hd__inv_6
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1107 _6476_/Q VGND VGND VPWR VPWR _3972_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5022_ _4689_/B _5017_/B _5021_/X VGND VGND VPWR VPWR _5079_/B sky130_fd_sc_hd__o21ai_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1118 _4296_/X VGND VGND VPWR VPWR _6742_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1129 _6603_/Q VGND VGND VPWR VPWR _4138_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6973_ _7049_/CLK _6973_/D fanout522/X VGND VGND VPWR VPWR _6973_/Q sky130_fd_sc_hd__dfrtp_4
X_5924_ _6598_/Q _5691_/Y _5913_/X _5923_/X _6318_/S VGND VGND VPWR VPWR _5924_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_22_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5855_ _6897_/Q _5655_/X _5706_/X _6505_/Q VGND VGND VPWR VPWR _5855_/X sky130_fd_sc_hd__a22o_1
XFILLER_167_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4806_ _4971_/A _4797_/A _4607_/D _4574_/Y VGND VGND VPWR VPWR _4806_/X sky130_fd_sc_hd__a31o_1
XFILLER_167_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5786_ _6902_/Q _5693_/X _5703_/X _6854_/Q _5776_/X VGND VGND VPWR VPWR _5786_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_166_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4737_ _4758_/C _5001_/C VGND VGND VPWR VPWR _4739_/B sky130_fd_sc_hd__nand2_1
XFILLER_119_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4668_ _5021_/A _4739_/A VGND VGND VPWR VPWR _4668_/X sky130_fd_sc_hd__or2_2
XFILLER_107_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3619_ input45/X _3308_/Y hold22/A _6900_/Q _3618_/X VGND VGND VPWR VPWR _3633_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_162_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6407_ _6407_/A _6407_/B VGND VGND VPWR VPWR _6407_/X sky130_fd_sc_hd__and2_1
Xhold930 _6702_/Q VGND VGND VPWR VPWR hold930/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold941 _4030_/X VGND VGND VPWR VPWR _6522_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4599_ _5115_/A _4599_/B _4984_/A _4584_/X VGND VGND VPWR VPWR _4599_/X sky130_fd_sc_hd__or4b_1
XFILLER_190_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold952 _6549_/Q VGND VGND VPWR VPWR hold952/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold963 _5213_/X VGND VGND VPWR VPWR _6812_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6338_ _6720_/Q _6023_/B _6338_/B1 _6770_/Q VGND VGND VPWR VPWR _6338_/X sky130_fd_sc_hd__a22o_1
Xhold974 _4086_/X VGND VGND VPWR VPWR _6561_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold985 _7015_/Q VGND VGND VPWR VPWR hold985/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold996 _5328_/X VGND VGND VPWR VPWR _6911_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6269_ _7183_/Q _5592_/Y _5650_/Y VGND VGND VPWR VPWR _6269_/X sky130_fd_sc_hd__o21ba_1
XFILLER_135_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_2_3_0_csclk clkbuf_2_3_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_7_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3970_ _3970_/A0 _6394_/A0 _3982_/S VGND VGND VPWR VPWR _3970_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5640_ _7158_/Q _7157_/Q VGND VGND VPWR VPWR _6040_/B sky130_fd_sc_hd__and2b_4
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5571_ _5571_/A _5571_/B VGND VGND VPWR VPWR _5579_/S sky130_fd_sc_hd__nand2_8
X_4522_ _4738_/A _5002_/A _4519_/X _4520_/X _5054_/A VGND VGND VPWR VPWR _4522_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_172_731 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold204 _5234_/X VGND VGND VPWR VPWR _6827_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 _6904_/Q VGND VGND VPWR VPWR hold215/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold226 _4303_/X VGND VGND VPWR VPWR _6748_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4453_ _4453_/A _4724_/A _4453_/C VGND VGND VPWR VPWR _5002_/A sky130_fd_sc_hd__or3_4
XFILLER_172_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold237 hold237/A VGND VGND VPWR VPWR hold237/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold248 _5406_/X VGND VGND VPWR VPWR _6980_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold259 _7099_/Q VGND VGND VPWR VPWR hold259/X sky130_fd_sc_hd__dlygate4sd3_1
X_3404_ _6960_/Q _3320_/Y _5331_/A _6920_/Q _3403_/X VGND VGND VPWR VPWR _3408_/B
+ sky130_fd_sc_hd__a221o_1
X_7172_ _7187_/CLK _7172_/D fanout488/X VGND VGND VPWR VPWR _7172_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_144_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4384_ _4570_/D _4385_/B VGND VGND VPWR VPWR _4999_/B sky130_fd_sc_hd__nor2_8
XFILLER_98_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6123_ _7131_/Q _6320_/A2 _6320_/B1 _6878_/Q VGND VGND VPWR VPWR _6123_/X sky130_fd_sc_hd__a22o_1
X_3335_ _3546_/A hold29/X VGND VGND VPWR VPWR _3335_/Y sky130_fd_sc_hd__nor2_2
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6054_ _6987_/Q _6203_/A2 _6024_/C _6907_/Q VGND VGND VPWR VPWR _6054_/X sky130_fd_sc_hd__a22o_1
XFILLER_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3266_ hold55/X hold27/X VGND VGND VPWR VPWR hold56/A sky130_fd_sc_hd__and2b_4
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5005_ _4931_/B _4744_/C _5001_/C _4896_/B _4822_/A VGND VGND VPWR VPWR _5134_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3197_ _7138_/Q VGND VGND VPWR VPWR _3197_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6956_ _7129_/CLK _6956_/D fanout526/X VGND VGND VPWR VPWR _6956_/Q sky130_fd_sc_hd__dfrtp_4
X_5907_ _6518_/Q _5966_/B1 _5699_/X _6538_/Q VGND VGND VPWR VPWR _5907_/X sky130_fd_sc_hd__a22o_1
X_6887_ _6925_/CLK _6887_/D fanout516/X VGND VGND VPWR VPWR _6887_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5838_ _5838_/A0 _5837_/X _6171_/S VGND VGND VPWR VPWR _5838_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5769_ _6877_/Q _5667_/X _5675_/X _6965_/Q _5768_/X VGND VGND VPWR VPWR _5770_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_6_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold760 _4151_/X VGND VGND VPWR VPWR _6614_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 _7022_/Q VGND VGND VPWR VPWR hold771/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold782 _5420_/X VGND VGND VPWR VPWR _6993_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold793 hold793/A VGND VGND VPWR VPWR hold793/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1460 _6680_/Q VGND VGND VPWR VPWR _3979_/S sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1471 _6789_/Q VGND VGND VPWR VPWR _3412_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1482 hold11/A VGND VGND VPWR VPWR _3874_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1493 _6633_/Q VGND VGND VPWR VPWR _4173_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput309 _3380_/X VGND VGND VPWR VPWR serial_data_2 sky130_fd_sc_hd__buf_12
XFILLER_181_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6810_ _7033_/CLK _6810_/D fanout503/X VGND VGND VPWR VPWR _6810_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_63_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6741_ _7211_/CLK _6741_/D fanout488/X VGND VGND VPWR VPWR _6741_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_50_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3953_ _6459_/Q _3953_/B VGND VGND VPWR VPWR _3953_/X sky130_fd_sc_hd__and2b_4
XFILLER_189_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6672_ _6683_/CLK hold45/X fanout511/X VGND VGND VPWR VPWR _6672_/Q sky130_fd_sc_hd__dfstp_1
X_3884_ _3884_/A _3884_/B input131/X input169/X VGND VGND VPWR VPWR _3886_/C sky130_fd_sc_hd__or4bb_1
XFILLER_31_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5623_ _7151_/Q _5624_/B _5622_/B _5625_/S VGND VGND VPWR VPWR _7151_/D sky130_fd_sc_hd__a31o_1
XFILLER_136_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5554_ _5581_/A0 _5554_/A1 _5561_/S VGND VGND VPWR VPWR _5554_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4505_ _4738_/A _4424_/Y _4503_/X _4504_/X VGND VGND VPWR VPWR _4505_/X sky130_fd_sc_hd__o211a_1
X_5485_ _5536_/A1 _5485_/A1 _5492_/S VGND VGND VPWR VPWR _5485_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4436_ _4793_/A _4436_/B VGND VGND VPWR VPWR _4744_/C sky130_fd_sc_hd__nor2_1
Xfanout503 fanout504/X VGND VGND VPWR VPWR fanout503/X sky130_fd_sc_hd__buf_4
XFILLER_120_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7155_ _7181_/CLK _7155_/D fanout502/X VGND VGND VPWR VPWR _7155_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout514 fanout526/X VGND VGND VPWR VPWR fanout514/X sky130_fd_sc_hd__buf_8
X_4367_ _4846_/B _4367_/B VGND VGND VPWR VPWR _4471_/B sky130_fd_sc_hd__nand2_2
XFILLER_86_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout525 fanout526/X VGND VGND VPWR VPWR fanout525/X sky130_fd_sc_hd__buf_6
X_3318_ _3528_/A hold68/X VGND VGND VPWR VPWR _3318_/Y sky130_fd_sc_hd__nor2_4
X_6106_ _6869_/Q _6199_/B1 _6027_/D _6885_/Q _6105_/X VGND VGND VPWR VPWR _6109_/C
+ sky130_fd_sc_hd__a221o_1
X_7086_ _7107_/CLK _7086_/D fanout515/X VGND VGND VPWR VPWR _7086_/Q sky130_fd_sc_hd__dfrtp_1
X_4298_ _6396_/A0 hold548/X _4299_/S VGND VGND VPWR VPWR _4298_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3249_ hold16/X hold72/X _3248_/Y VGND VGND VPWR VPWR hold17/A sky130_fd_sc_hd__a21bo_1
X_6037_ _7119_/Q _6323_/B1 _6329_/B1 _7034_/Q VGND VGND VPWR VPWR _6037_/X sky130_fd_sc_hd__a22o_1
XFILLER_73_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6939_ _7128_/CLK _6939_/D fanout514/X VGND VGND VPWR VPWR _6939_/Q sky130_fd_sc_hd__dfstp_1
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_csclk _3942_/X VGND VGND VPWR VPWR clkbuf_0_csclk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_136_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold590 _5274_/X VGND VGND VPWR VPWR _6863_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_173_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_1_0_1_csclk/A sky130_fd_sc_hd__clkbuf_8
XFILLER_18_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1290 _5530_/X VGND VGND VPWR VPWR _7090_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5270_ _5555_/A0 hold353/X _5276_/S VGND VGND VPWR VPWR _5270_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4221_ _5534_/A1 hold685/X _4221_/S VGND VGND VPWR VPWR _4221_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4152_ _5534_/A1 hold717/X _4152_/S VGND VGND VPWR VPWR _4152_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4083_ hold227/X _5569_/A0 _4083_/S VGND VGND VPWR VPWR _4083_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4985_ _4985_/A _4985_/B _4985_/C VGND VGND VPWR VPWR _4988_/B sky130_fd_sc_hd__or3_1
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6724_ _6725_/CLK _6724_/D fanout510/X VGND VGND VPWR VPWR _6724_/Q sky130_fd_sc_hd__dfrtp_4
X_3936_ _6573_/Q user_clock _6822_/Q VGND VGND VPWR VPWR _3936_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_3_2_0_csclk clkbuf_3_3_0_csclk/A VGND VGND VPWR VPWR clkbuf_3_2_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_149_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6655_ _6708_/CLK _6655_/D _6432_/A VGND VGND VPWR VPWR _6655_/Q sky130_fd_sc_hd__dfrtp_4
X_3867_ _6473_/Q _6471_/Q _6541_/Q VGND VGND VPWR VPWR _3868_/B sky130_fd_sc_hd__and3_1
XFILLER_31_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5606_ _5606_/A _5606_/B _5606_/C VGND VGND VPWR VPWR _7146_/D sky130_fd_sc_hd__and3_1
XFILLER_137_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6586_ _7136_/CLK hold98/X fanout520/X VGND VGND VPWR VPWR _6586_/Q sky130_fd_sc_hd__dfrtp_1
X_3798_ _3798_/A _3800_/A VGND VGND VPWR VPWR _6473_/D sky130_fd_sc_hd__xor2_1
XFILLER_118_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5537_ hold371/X _5555_/A0 _5543_/S VGND VGND VPWR VPWR _5537_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5468_ hold359/X _5555_/A0 _5474_/S VGND VGND VPWR VPWR _5468_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7207_ _7207_/CLK _7207_/D fanout485/X VGND VGND VPWR VPWR _7207_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_78_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4419_ _4846_/B _4846_/A _4667_/C VGND VGND VPWR VPWR _4459_/B sky130_fd_sc_hd__and3b_4
XFILLER_99_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5399_ hold705/X _5567_/A0 _5402_/S VGND VGND VPWR VPWR _5399_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7138_ _7138_/CLK _7138_/D fanout520/X VGND VGND VPWR VPWR _7138_/Q sky130_fd_sc_hd__dfrtp_2
Xfanout366 _6171_/S VGND VGND VPWR VPWR _6319_/S sky130_fd_sc_hd__buf_8
XFILLER_101_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7069_ _7134_/CLK _7069_/D fanout521/X VGND VGND VPWR VPWR _7069_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput19 mask_rev_in[23] VGND VGND VPWR VPWR input19/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_260 hold127/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4770_ _4822_/A _4770_/B _4770_/C _4882_/B VGND VGND VPWR VPWR _4770_/X sky130_fd_sc_hd__or4b_1
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3721_ _3721_/A _3721_/B _3721_/C _3721_/D VGND VGND VPWR VPWR _3722_/D sky130_fd_sc_hd__or4_1
XFILLER_158_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6440_ _6441_/A _6440_/B VGND VGND VPWR VPWR _6440_/X sky130_fd_sc_hd__and2_1
X_3652_ _6980_/Q _5403_/A _3471_/Y _6763_/Q VGND VGND VPWR VPWR _3652_/X sky130_fd_sc_hd__a22o_1
XFILLER_174_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3583_ _3583_/A _3583_/B _3583_/C _3583_/D VGND VGND VPWR VPWR _3601_/A sky130_fd_sc_hd__or4_2
XFILLER_127_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6371_ _6370_/X _6371_/A1 _6386_/S VGND VGND VPWR VPWR _7199_/D sky130_fd_sc_hd__mux2_1
XFILLER_173_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5322_ _5322_/A _5571_/B VGND VGND VPWR VPWR _5330_/S sky130_fd_sc_hd__and2_4
XFILLER_173_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5253_ hold217/X _5583_/A0 _5258_/S VGND VGND VPWR VPWR _5253_/X sky130_fd_sc_hd__mux2_1
X_4204_ _4204_/A _6392_/B VGND VGND VPWR VPWR _4209_/S sky130_fd_sc_hd__and2_2
X_5184_ _5184_/A _6392_/B VGND VGND VPWR VPWR _5186_/S sky130_fd_sc_hd__nand2_1
X_4135_ _4135_/A _6392_/B VGND VGND VPWR VPWR _4140_/S sky130_fd_sc_hd__and2_1
XFILLER_29_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_63_csclk _6753_/CLK VGND VGND VPWR VPWR _7074_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_113_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4066_ _4118_/A1 _5569_/A0 _4068_/S VGND VGND VPWR VPWR _4066_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_78_csclk _6753_/CLK VGND VGND VPWR VPWR _6664_/CLK sky130_fd_sc_hd__clkbuf_16
X_4968_ _4969_/B VGND VGND VPWR VPWR _5100_/A sky130_fd_sc_hd__clkinv_2
XFILLER_149_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6707_ _6707_/CLK _6707_/D fanout496/X VGND VGND VPWR VPWR _6707_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_165_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3919_ _6578_/Q input89/X _3921_/S VGND VGND VPWR VPWR _3919_/X sky130_fd_sc_hd__mux2_2
X_4899_ _5059_/A _4899_/B VGND VGND VPWR VPWR _5130_/B sky130_fd_sc_hd__or2_1
XFILLER_20_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6638_ _6709_/CLK _6638_/D fanout494/X VGND VGND VPWR VPWR _6638_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_192_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6569_ _6925_/CLK _6569_/D fanout516/X VGND VGND VPWR VPWR _6569_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_16_csclk _6882_/CLK VGND VGND VPWR VPWR _7082_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_79_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5940_ _6524_/Q _5694_/X _5703_/X _6604_/Q _5939_/X VGND VGND VPWR VPWR _5945_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_46_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5871_ _6634_/Q _5655_/X _5666_/X _6686_/Q _5870_/X VGND VGND VPWR VPWR _5879_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4822_ _4822_/A _4822_/B _4822_/C _4882_/A VGND VGND VPWR VPWR _4823_/C sky130_fd_sc_hd__or4b_1
X_4753_ _4981_/B _4996_/A VGND VGND VPWR VPWR _4753_/Y sky130_fd_sc_hd__nor2_1
XFILLER_147_634 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3704_ _6712_/Q _4258_/A _4159_/A _6622_/Q VGND VGND VPWR VPWR _3704_/X sky130_fd_sc_hd__a22o_1
X_4684_ _4684_/A _4684_/B VGND VGND VPWR VPWR _4860_/B sky130_fd_sc_hd__nand2_2
X_6423_ _6441_/A _6440_/B VGND VGND VPWR VPWR _6423_/X sky130_fd_sc_hd__and2_1
X_3635_ _7068_/Q _5502_/A _5448_/A _7020_/Q _3634_/X VGND VGND VPWR VPWR _3642_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6354_ _6354_/A0 _3447_/X _6356_/S VGND VGND VPWR VPWR _7194_/D sky130_fd_sc_hd__mux2_1
X_3566_ input46/X _3308_/Y _5562_/A _7122_/Q _3565_/X VGND VGND VPWR VPWR _3573_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5305_ _5581_/A0 _5305_/A1 _5312_/S VGND VGND VPWR VPWR _5305_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3497_ _6802_/Q _5193_/A _4129_/A _6600_/Q VGND VGND VPWR VPWR _3497_/X sky130_fd_sc_hd__a22o_1
X_6285_ _6688_/Q _6024_/A _6040_/X _6528_/Q VGND VGND VPWR VPWR _6285_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5236_ _5584_/A0 hold451/X _5240_/S VGND VGND VPWR VPWR _5236_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5167_ _5148_/Y _5151_/X _5166_/Y _5147_/X VGND VGND VPWR VPWR _5167_/X sky130_fd_sc_hd__a211o_1
XFILLER_29_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4118_ _5569_/A0 _4118_/A1 hold97/X VGND VGND VPWR VPWR hold98/A sky130_fd_sc_hd__mux2_1
XFILLER_56_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5098_ _4997_/A _4728_/Y _4989_/C _4618_/D VGND VGND VPWR VPWR _5142_/B sky130_fd_sc_hd__o211ai_1
X_4049_ _6395_/A0 _4049_/A1 _4051_/S VGND VGND VPWR VPWR _4049_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_692 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold8 hold8/A VGND VGND VPWR VPWR hold8/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_87_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire383 _3547_/B VGND VGND VPWR VPWR _3714_/B sky130_fd_sc_hd__buf_12
Xhold408 _5423_/X VGND VGND VPWR VPWR _6995_/D sky130_fd_sc_hd__dlygate4sd3_1
Xwire394 _6023_/D VGND VGND VPWR VPWR wire394/X sky130_fd_sc_hd__buf_8
Xhold419 _7087_/Q VGND VGND VPWR VPWR hold419/X sky130_fd_sc_hd__dlygate4sd3_1
X_3420_ _6479_/Q _3966_/A _5448_/A _7023_/Q VGND VGND VPWR VPWR _3420_/X sky130_fd_sc_hd__a22o_1
XFILLER_109_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3351_ _7118_/Q _5553_/A _5439_/A _7017_/Q VGND VGND VPWR VPWR _3351_/X sky130_fd_sc_hd__a22o_1
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6070_ _6843_/Q _6046_/B _6069_/X _6318_/S VGND VGND VPWR VPWR _6070_/X sky130_fd_sc_hd__o211a_1
X_3282_ hold74/X hold66/X VGND VGND VPWR VPWR _3283_/A sky130_fd_sc_hd__nand2_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1108 _3972_/X VGND VGND VPWR VPWR _6476_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5021_ _5021_/A _5021_/B _5021_/C VGND VGND VPWR VPWR _5021_/X sky130_fd_sc_hd__or3_1
XFILLER_112_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1119 _7129_/Q VGND VGND VPWR VPWR _5574_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6972_ _7075_/CLK _6972_/D fanout514/X VGND VGND VPWR VPWR _6972_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_19_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5923_ _5923_/A _5923_/B _5923_/C _5923_/D VGND VGND VPWR VPWR _5923_/X sky130_fd_sc_hd__or4_1
XFILLER_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5854_ _6993_/Q _5697_/X _5702_/X _6985_/Q _5853_/X VGND VGND VPWR VPWR _5857_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_110_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4805_ _4814_/A _4683_/A _5076_/B _4996_/A _4802_/A VGND VGND VPWR VPWR _4805_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_167_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5785_ _5785_/A _5785_/B _5785_/C _5785_/D VGND VGND VPWR VPWR _5785_/X sky130_fd_sc_hd__or4_1
XFILLER_166_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4736_ _4981_/B _4997_/A VGND VGND VPWR VPWR _5049_/B sky130_fd_sc_hd__nor2_1
XFILLER_159_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4667_ _4596_/A _4732_/A _4667_/C VGND VGND VPWR VPWR _4667_/X sky130_fd_sc_hd__and3b_1
XFILLER_134_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6406_ _6407_/A _6407_/B VGND VGND VPWR VPWR _6406_/X sky130_fd_sc_hd__and2_1
Xhold920 _6504_/Q VGND VGND VPWR VPWR hold920/X sky130_fd_sc_hd__dlygate4sd3_1
X_3618_ _7129_/Q _5571_/A _4288_/A _6738_/Q VGND VGND VPWR VPWR _3618_/X sky130_fd_sc_hd__a22o_1
XFILLER_162_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold931 _4248_/X VGND VGND VPWR VPWR _6702_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4598_ _4965_/A _4598_/B _4983_/A _4598_/D VGND VGND VPWR VPWR _4599_/B sky130_fd_sc_hd__or4_1
Xhold942 _6707_/Q VGND VGND VPWR VPWR hold942/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold953 _4061_/X VGND VGND VPWR VPWR _6549_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6337_ _6690_/Q _6024_/A wire394/X _6638_/Q VGND VGND VPWR VPWR _6337_/X sky130_fd_sc_hd__a22o_1
Xhold964 _6681_/Q VGND VGND VPWR VPWR hold964/X sky130_fd_sc_hd__dlygate4sd3_1
X_3549_ input38/X _3751_/A2 _4300_/A _6749_/Q VGND VGND VPWR VPWR _3549_/X sky130_fd_sc_hd__a22o_1
Xhold975 _6548_/Q VGND VGND VPWR VPWR hold975/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold986 _5445_/X VGND VGND VPWR VPWR _7015_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold997 _6855_/Q VGND VGND VPWR VPWR hold997/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6268_ _6597_/Q _6046_/B _6257_/X _6267_/X _6318_/S VGND VGND VPWR VPWR _6268_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_135_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5219_ _5587_/A0 hold876/X _5220_/S VGND VGND VPWR VPWR _5219_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6199_ _7057_/Q _5988_/X _6199_/B1 _6873_/Q VGND VGND VPWR VPWR _6216_/A sky130_fd_sc_hd__a22o_1
XFILLER_130_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_610 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5570_ _5579_/A0 hold393/X _5570_/S VGND VGND VPWR VPWR _5570_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4521_ _4657_/C _4524_/B VGND VGND VPWR VPWR _5054_/A sky130_fd_sc_hd__nand2_1
XFILLER_144_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold205 _6845_/Q VGND VGND VPWR VPWR hold205/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold216 _5320_/X VGND VGND VPWR VPWR _6904_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4452_ _4758_/A _5001_/A _4758_/B _4657_/C VGND VGND VPWR VPWR _5165_/D sky130_fd_sc_hd__nand4_1
Xhold227 hold227/A VGND VGND VPWR VPWR hold227/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold238 _4113_/X VGND VGND VPWR VPWR _6581_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 _7068_/Q VGND VGND VPWR VPWR hold249/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_618 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3403_ _6888_/Q _3318_/Y _5221_/B _3380_/X VGND VGND VPWR VPWR _3403_/X sky130_fd_sc_hd__a22o_1
X_7171_ _7187_/CLK _7171_/D fanout488/X VGND VGND VPWR VPWR _7171_/Q sky130_fd_sc_hd__dfrtp_1
X_4383_ _4846_/A _4846_/B VGND VGND VPWR VPWR _4385_/B sky130_fd_sc_hd__nand2_2
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6122_ _6145_/A0 _6121_/X _6319_/S VGND VGND VPWR VPWR _7178_/D sky130_fd_sc_hd__mux2_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3334_ _3334_/A hold76/X VGND VGND VPWR VPWR _3334_/Y sky130_fd_sc_hd__nor2_4
XFILLER_124_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6053_ _7003_/Q _6202_/B1 _6272_/B _7067_/Q _6049_/X VGND VGND VPWR VPWR _6058_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3265_ hold26/X _4776_/B2 _3971_/S VGND VGND VPWR VPWR hold27/A sky130_fd_sc_hd__mux2_4
XFILLER_105_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5004_ _4999_/B _4838_/B _5158_/A VGND VGND VPWR VPWR _5148_/B sky130_fd_sc_hd__a21o_1
XFILLER_38_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3196_ _6564_/Q VGND VGND VPWR VPWR _5650_/B sky130_fd_sc_hd__clkinv_2
XFILLER_38_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6955_ _7070_/CLK _6955_/D fanout510/X VGND VGND VPWR VPWR _6955_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_41_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5906_ _6703_/Q _5659_/X _5667_/X _6618_/Q _5905_/X VGND VGND VPWR VPWR _5913_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_22_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6886_ _7123_/CLK _6886_/D _6407_/A VGND VGND VPWR VPWR _6886_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_22_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5837_ _5650_/A _7167_/Q _5836_/X VGND VGND VPWR VPWR _5837_/X sky130_fd_sc_hd__a21o_1
XFILLER_10_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5768_ _6973_/Q _5691_/B _5699_/X _7053_/Q _5690_/X VGND VGND VPWR VPWR _5768_/X
+ sky130_fd_sc_hd__a221o_1
X_4719_ _4719_/A _5016_/A VGND VGND VPWR VPWR _4720_/C sky130_fd_sc_hd__nor2_1
XFILLER_108_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5699_ _7152_/Q _5699_/B _5699_/C VGND VGND VPWR VPWR _5699_/X sky130_fd_sc_hd__and3_4
XFILLER_107_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold750 _4315_/X VGND VGND VPWR VPWR _6758_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold761 _6539_/Q VGND VGND VPWR VPWR hold761/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold772 _5453_/X VGND VGND VPWR VPWR _7022_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap480 _4951_/B VGND VGND VPWR VPWR _4376_/B sky130_fd_sc_hd__clkbuf_2
Xhold783 hold783/A VGND VGND VPWR VPWR hold783/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold794 _4112_/X VGND VGND VPWR VPWR _6580_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1450 _7193_/Q VGND VGND VPWR VPWR _6353_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1461 _3979_/X VGND VGND VPWR VPWR hold100/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1472 _6776_/Q VGND VGND VPWR VPWR _4776_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1483 _7192_/Q VGND VGND VPWR VPWR _6352_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1494 _7177_/Q VGND VGND VPWR VPWR _6121_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6740_ _6740_/CLK _6740_/D fanout510/X VGND VGND VPWR VPWR _6740_/Q sky130_fd_sc_hd__dfrtp_2
X_3952_ _6460_/Q _3952_/B VGND VGND VPWR VPWR _3952_/X sky130_fd_sc_hd__and2b_4
XFILLER_189_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6671_ _7094_/CLK _6671_/D fanout494/X VGND VGND VPWR VPWR _6671_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_189_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3883_ _4390_/C _4390_/D VGND VGND VPWR VPWR _4654_/B sky130_fd_sc_hd__or2_1
X_5622_ _7151_/Q _5622_/B VGND VGND VPWR VPWR _5625_/S sky130_fd_sc_hd__nor2_1
XFILLER_149_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5553_ _5553_/A _5571_/B VGND VGND VPWR VPWR _5561_/S sky130_fd_sc_hd__nand2_8
XFILLER_157_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4504_ _4504_/A _4504_/B _4860_/A VGND VGND VPWR VPWR _4504_/X sky130_fd_sc_hd__and3_1
X_5484_ _5484_/A _5535_/B VGND VGND VPWR VPWR _5492_/S sky130_fd_sc_hd__nand2_8
XFILLER_144_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4435_ _4435_/A _4435_/B VGND VGND VPWR VPWR _4453_/C sky130_fd_sc_hd__nand2_2
XFILLER_160_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7154_ _7181_/CLK _7154_/D fanout500/X VGND VGND VPWR VPWR _7154_/Q sky130_fd_sc_hd__dfstp_1
Xfanout504 fanout508/X VGND VGND VPWR VPWR fanout504/X sky130_fd_sc_hd__buf_8
Xfanout515 fanout526/X VGND VGND VPWR VPWR fanout515/X sky130_fd_sc_hd__buf_4
X_4366_ _4369_/B VGND VGND VPWR VPWR _4367_/B sky130_fd_sc_hd__inv_2
Xfanout526 fanout527/X VGND VGND VPWR VPWR fanout526/X sky130_fd_sc_hd__buf_12
XFILLER_59_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6105_ _6853_/Q _6027_/A _5988_/X _7053_/Q VGND VGND VPWR VPWR _6105_/X sky130_fd_sc_hd__a22o_1
XFILLER_59_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3317_ hold21/X _5241_/B VGND VGND VPWR VPWR hold22/A sky130_fd_sc_hd__nor2_8
X_7085_ _7138_/CLK _7085_/D fanout524/X VGND VGND VPWR VPWR _7085_/Q sky130_fd_sc_hd__dfrtp_4
X_4297_ _6395_/A0 _4297_/A1 _4299_/S VGND VGND VPWR VPWR _4297_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6036_ _6040_/B _6039_/C _6040_/C VGND VGND VPWR VPWR _6036_/X sky130_fd_sc_hd__and3_4
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3248_ _3248_/A _3252_/B VGND VGND VPWR VPWR _3248_/Y sky130_fd_sc_hd__nand2_1
XFILLER_27_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6938_ _7123_/CLK _6938_/D fanout519/X VGND VGND VPWR VPWR _6938_/Q sky130_fd_sc_hd__dfstp_4
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6869_ _7049_/CLK _6869_/D fanout522/X VGND VGND VPWR VPWR _6869_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_10_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold580 _4305_/X VGND VGND VPWR VPWR _6750_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold591 _6485_/Q VGND VGND VPWR VPWR hold591/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1280 _4211_/X VGND VGND VPWR VPWR _6665_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1291 _6756_/Q VGND VGND VPWR VPWR _4313_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4220_ _5533_/A1 hold689/X _4221_/S VGND VGND VPWR VPWR _4220_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4151_ _5533_/A1 hold759/X _4152_/S VGND VGND VPWR VPWR _4151_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4082_ hold403/X _4081_/X _4086_/S VGND VGND VPWR VPWR _4082_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4984_ _4984_/A _4984_/B _4984_/C VGND VGND VPWR VPWR _5090_/B sky130_fd_sc_hd__or3_1
XFILLER_51_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6723_ _6725_/CLK _6723_/D fanout509/X VGND VGND VPWR VPWR _6723_/Q sky130_fd_sc_hd__dfstp_2
X_3935_ _3233_/Y input2/X input1/X VGND VGND VPWR VPWR _3935_/X sky130_fd_sc_hd__mux2_4
XFILLER_149_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6654_ _7193_/CLK _6654_/D VGND VGND VPWR VPWR _6654_/Q sky130_fd_sc_hd__dfxtp_1
X_3866_ input58/X _3866_/A1 _3866_/S VGND VGND VPWR VPWR _6446_/D sky130_fd_sc_hd__mux2_1
X_5605_ _5605_/A VGND VGND VPWR VPWR _5606_/C sky130_fd_sc_hd__clkinv_2
X_6585_ _7130_/CLK _6585_/D fanout519/X VGND VGND VPWR VPWR _6585_/Q sky130_fd_sc_hd__dfrtp_1
X_3797_ _6473_/Q _6472_/Q VGND VGND VPWR VPWR _3838_/B sky130_fd_sc_hd__and2_1
XFILLER_176_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5536_ _5536_/A0 _5536_/A1 _5543_/S VGND VGND VPWR VPWR _5536_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5467_ _5467_/A0 _5536_/A1 _5474_/S VGND VGND VPWR VPWR _5467_/X sky130_fd_sc_hd__mux2_1
X_7206_ _3937_/A1 _7206_/D fanout529/X VGND VGND VPWR VPWR _7206_/Q sky130_fd_sc_hd__dfrtp_1
X_4418_ _4742_/A _4876_/A VGND VGND VPWR VPWR _4503_/C sky130_fd_sc_hd__nand2_1
X_5398_ hold659/X _5557_/A0 _5402_/S VGND VGND VPWR VPWR _5398_/X sky130_fd_sc_hd__mux2_1
XFILLER_120_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7137_ _7137_/CLK _7137_/D fanout508/X VGND VGND VPWR VPWR _7137_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4349_ _4404_/B _4350_/B _4654_/A VGND VGND VPWR VPWR _4351_/A sky130_fd_sc_hd__a21o_1
XFILLER_86_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7068_ _7068_/CLK _7068_/D fanout505/X VGND VGND VPWR VPWR _7068_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_86_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6019_ _6019_/A _6019_/B VGND VGND VPWR VPWR _6025_/C sky130_fd_sc_hd__nor2_4
XFILLER_100_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_250 _6822_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_261 _4083_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3720_ _6867_/Q _5277_/A hold50/A hold87/A _3719_/X VGND VGND VPWR VPWR _3721_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_119_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3651_ _3651_/A _3651_/B _3651_/C _3651_/D VGND VGND VPWR VPWR _3659_/A sky130_fd_sc_hd__or4_1
XFILLER_158_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6370_ _6700_/Q _6370_/A2 _6370_/B1 _6390_/A2 _6369_/X VGND VGND VPWR VPWR _6370_/X
+ sky130_fd_sc_hd__a221o_1
X_3582_ _3582_/A _3582_/B _3582_/C _3582_/D VGND VGND VPWR VPWR _3583_/D sky130_fd_sc_hd__or4_1
XFILLER_127_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5321_ _5579_/A0 hold536/X hold23/X VGND VGND VPWR VPWR _5321_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5252_ hold347/X _5555_/A0 _5258_/S VGND VGND VPWR VPWR _5252_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4203_ hold365/X _5534_/A1 _4203_/S VGND VGND VPWR VPWR _4203_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5183_ _5183_/A _5183_/B _5183_/C VGND VGND VPWR VPWR _6782_/D sky130_fd_sc_hd__or3_1
XFILLER_3_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4134_ hold463/X _6397_/A0 _4134_/S VGND VGND VPWR VPWR _4134_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4065_ hold956/X _4064_/X _4069_/S VGND VGND VPWR VPWR _4065_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4967_ _4794_/A _4784_/A _5016_/A _4810_/D _4887_/D VGND VGND VPWR VPWR _4969_/B
+ sky130_fd_sc_hd__o311a_1
X_6706_ _6708_/CLK _6706_/D fanout496/X VGND VGND VPWR VPWR _6706_/Q sky130_fd_sc_hd__dfrtp_4
X_3918_ _6579_/Q input91/X _3921_/S VGND VGND VPWR VPWR _3918_/X sky130_fd_sc_hd__mux2_4
XFILLER_20_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4898_ _5042_/A _4873_/Y _4875_/X _4897_/X _4992_/C VGND VGND VPWR VPWR _4928_/C
+ sky130_fd_sc_hd__o41a_1
XFILLER_177_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6637_ _7094_/CLK _6637_/D fanout494/X VGND VGND VPWR VPWR _6637_/Q sky130_fd_sc_hd__dfrtp_4
X_3849_ _6473_/Q _6472_/Q _6541_/Q _3848_/Y VGND VGND VPWR VPWR _3856_/B sky130_fd_sc_hd__o211a_1
XFILLER_192_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6568_ _6925_/CLK _6568_/D fanout516/X VGND VGND VPWR VPWR _6568_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5519_ _5552_/A0 hold757/X _5519_/S VGND VGND VPWR VPWR _5519_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6499_ _7128_/CLK _6499_/D fanout514/X VGND VGND VPWR VPWR _6499_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_105_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_76 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5870_ _6771_/Q _5663_/X _5664_/X _6751_/Q VGND VGND VPWR VPWR _5870_/X sky130_fd_sc_hd__a22o_1
X_4821_ _4982_/B _4821_/B _4821_/C _4821_/D VGND VGND VPWR VPWR _4822_/B sky130_fd_sc_hd__or4_1
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4752_ _4996_/A _5036_/A VGND VGND VPWR VPWR _4986_/B sky130_fd_sc_hd__nor2_1
X_3703_ _6843_/Q _5250_/A _4198_/A _6656_/Q _3702_/X VGND VGND VPWR VPWR _3710_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_119_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_646 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4683_ _4683_/A _4683_/B VGND VGND VPWR VPWR _4699_/B sky130_fd_sc_hd__or2_1
X_6422_ _6441_/A _6440_/B VGND VGND VPWR VPWR _6422_/X sky130_fd_sc_hd__and2_1
X_3634_ _7060_/Q _5493_/A _4028_/A _6523_/Q VGND VGND VPWR VPWR _3634_/X sky130_fd_sc_hd__a22o_1
X_6353_ _6353_/A0 _6353_/A1 _6356_/S VGND VGND VPWR VPWR _7193_/D sky130_fd_sc_hd__mux2_1
X_3565_ _6739_/Q _4288_/A _4270_/A _6724_/Q VGND VGND VPWR VPWR _3565_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5304_ _5304_/A _5580_/B VGND VGND VPWR VPWR _5312_/S sky130_fd_sc_hd__nand2_8
X_6284_ _6672_/Q _6340_/A2 wire394/X _6636_/Q _6283_/X VGND VGND VPWR VPWR _6291_/A
+ sky130_fd_sc_hd__a221o_1
X_3496_ _3714_/B _4120_/B VGND VGND VPWR VPWR _4129_/A sky130_fd_sc_hd__nor2_4
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5235_ _5574_/A0 _5235_/A1 _5240_/S VGND VGND VPWR VPWR _5235_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5166_ _5128_/C _5163_/X _5180_/C _5160_/X VGND VGND VPWR VPWR _5166_/Y sky130_fd_sc_hd__a31oi_2
XFILLER_68_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4117_ hold127/X _4117_/A1 hold97/X VGND VGND VPWR VPWR _4117_/X sky130_fd_sc_hd__mux2_1
X_5097_ _4870_/B _4783_/Y _5096_/X VGND VGND VPWR VPWR _5112_/D sky130_fd_sc_hd__a21o_1
XFILLER_83_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4048_ _6394_/A0 _4048_/A1 _4051_/S VGND VGND VPWR VPWR _4048_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5999_ _6986_/Q _6203_/A2 _5998_/Y _7010_/Q _5995_/X VGND VGND VPWR VPWR _6012_/B
+ sky130_fd_sc_hd__a221o_1
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput290 _6481_/Q VGND VGND VPWR VPWR pll_trim[23] sky130_fd_sc_hd__buf_12
Xhold9 hold9/A VGND VGND VPWR VPWR hold9/X sky130_fd_sc_hd__buf_6
XFILLER_47_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_62_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7115_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_116_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire362 _6069_/A VGND VGND VPWR VPWR _6168_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_128_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold409 _6560_/Q VGND VGND VPWR VPWR hold409/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_183_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3350_ input10/X _3295_/Y _3751_/A2 input42/X _3349_/X VGND VGND VPWR VPWR _3355_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_124_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_77_csclk _6753_/CLK VGND VGND VPWR VPWR _7209_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3281_ hold18/X _3301_/C hold94/X VGND VGND VPWR VPWR _3281_/X sky130_fd_sc_hd__or3_4
XFILLER_97_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ _4814_/A _4396_/X _4919_/X VGND VGND VPWR VPWR _5073_/B sky130_fd_sc_hd__o21ai_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1109 _6842_/Q VGND VGND VPWR VPWR _5251_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_65_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6971_ _7043_/CLK _6971_/D fanout514/X VGND VGND VPWR VPWR _6971_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_53_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5922_ _6623_/Q _5661_/X _5955_/A2 _6672_/Q _5921_/X VGND VGND VPWR VPWR _5923_/D
+ sky130_fd_sc_hd__a221o_2
XFILLER_179_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5853_ _7001_/Q _5656_/X _5670_/X _6937_/Q VGND VGND VPWR VPWR _5853_/X sky130_fd_sc_hd__a22o_1
XFILLER_110_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_15_csclk _6882_/CLK VGND VGND VPWR VPWR _7123_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_22_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4804_ _4674_/A _4569_/Y _4622_/Y _4746_/Y VGND VGND VPWR VPWR _4813_/C sky130_fd_sc_hd__a31o_1
X_5784_ _6878_/Q _5667_/X _5675_/X _6966_/Q _5783_/X VGND VGND VPWR VPWR _5785_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_166_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4735_ _4759_/A _4876_/A VGND VGND VPWR VPWR _4810_/C sky130_fd_sc_hd__nand2_1
XFILLER_147_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4666_ _5023_/A _4666_/B VGND VGND VPWR VPWR _4666_/Y sky130_fd_sc_hd__nor2_1
XFILLER_119_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6405_ _6407_/A _6407_/B VGND VGND VPWR VPWR _6405_/X sky130_fd_sc_hd__and2_1
X_3617_ _6988_/Q _5412_/A _4330_/A _6773_/Q VGND VGND VPWR VPWR _3658_/B sky130_fd_sc_hd__a22o_1
Xhold910 _7040_/Q VGND VGND VPWR VPWR hold910/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold921 _4008_/X VGND VGND VPWR VPWR _6504_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4597_ _4569_/B _5021_/B _4659_/B VGND VGND VPWR VPWR _4598_/D sky130_fd_sc_hd__a21oi_1
Xhold932 _6656_/Q VGND VGND VPWR VPWR hold932/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold943 _4254_/X VGND VGND VPWR VPWR _6707_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6336_ _6705_/Q _6336_/A2 _6272_/B _6535_/Q _6335_/X VGND VGND VPWR VPWR _6341_/C
+ sky130_fd_sc_hd__a221o_1
Xhold954 _6670_/Q VGND VGND VPWR VPWR hold954/X sky130_fd_sc_hd__dlygate4sd3_1
X_3548_ _6933_/Q _5349_/A _5358_/A _6941_/Q VGND VGND VPWR VPWR _3548_/X sky130_fd_sc_hd__a22o_1
Xhold965 _4235_/X VGND VGND VPWR VPWR _6681_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold976 _4059_/X VGND VGND VPWR VPWR _6548_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold987 _7124_/Q VGND VGND VPWR VPWR hold987/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_142_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold998 _5265_/X VGND VGND VPWR VPWR _6855_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6267_ _6292_/A _6267_/B _6267_/C VGND VGND VPWR VPWR _6267_/X sky130_fd_sc_hd__or3_1
XFILLER_88_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3479_ _6674_/Q _4216_/A _4246_/A _6705_/Q VGND VGND VPWR VPWR _3479_/X sky130_fd_sc_hd__a22o_1
XFILLER_130_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5218_ hold127/X hold251/X _5220_/S VGND VGND VPWR VPWR _5218_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6198_ _7089_/Q _5977_/X _6323_/B1 _7126_/Q VGND VGND VPWR VPWR _6198_/X sky130_fd_sc_hd__a22o_1
Xhold1610 _6574_/Q VGND VGND VPWR VPWR hold1610/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5149_ _4999_/B _4446_/Y _4843_/A _4965_/B _5009_/A VGND VGND VPWR VPWR _5151_/C
+ sky130_fd_sc_hd__a2111o_1
XFILLER_151_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4520_ _4739_/A _5002_/A VGND VGND VPWR VPWR _4520_/X sky130_fd_sc_hd__or2_1
XFILLER_156_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold206 _5254_/X VGND VGND VPWR VPWR _6845_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4451_ _4667_/C _4999_/B VGND VGND VPWR VPWR _4942_/A sky130_fd_sc_hd__nand2_2
Xhold217 _6844_/Q VGND VGND VPWR VPWR hold217/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 _4127_/X VGND VGND VPWR VPWR _6594_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold239 _6996_/Q VGND VGND VPWR VPWR hold239/X sky130_fd_sc_hd__dlygate4sd3_1
X_3402_ _6848_/Q _5250_/A _3308_/Y input50/X _3401_/X VGND VGND VPWR VPWR _3408_/A
+ sky130_fd_sc_hd__a221o_1
X_7170_ _7187_/CLK _7170_/D fanout488/X VGND VGND VPWR VPWR _7170_/Q sky130_fd_sc_hd__dfrtp_1
X_4382_ _5023_/A _4719_/A VGND VGND VPWR VPWR _4952_/A sky130_fd_sc_hd__nor2_1
XFILLER_171_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6121_ _5650_/A _6121_/A2 _6120_/X VGND VGND VPWR VPWR _6121_/X sky130_fd_sc_hd__a21o_1
XFILLER_98_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3333_ hold96/X _5241_/B VGND VGND VPWR VPWR _3333_/Y sky130_fd_sc_hd__nor2_2
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6052_ _7075_/Q _5994_/X _5998_/Y _7011_/Q _6051_/X VGND VGND VPWR VPWR _6058_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3264_ hold25/X input58/X hold72/A VGND VGND VPWR VPWR hold26/A sky130_fd_sc_hd__mux2_1
XFILLER_100_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5003_ _5003_/A _5036_/B VGND VGND VPWR VPWR _5008_/C sky130_fd_sc_hd__nor2_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3195_ _5650_/A VGND VGND VPWR VPWR _3195_/Y sky130_fd_sc_hd__inv_6
XFILLER_39_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6954_ _6990_/CLK _6954_/D _3873_/A VGND VGND VPWR VPWR _6954_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_41_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5905_ _6667_/Q _5677_/X _5694_/X _6523_/Q VGND VGND VPWR VPWR _5905_/X sky130_fd_sc_hd__a22o_1
X_6885_ _7140_/CLK _6885_/D fanout522/X VGND VGND VPWR VPWR _6885_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5836_ _6848_/Q _5691_/Y _5825_/X _5835_/X _6318_/S VGND VGND VPWR VPWR _5836_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_167_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5767_ _7021_/Q _5663_/X _5683_/X _6869_/Q _5755_/X VGND VGND VPWR VPWR _5770_/C
+ sky130_fd_sc_hd__a221o_1
X_4718_ _4745_/A _4718_/B VGND VGND VPWR VPWR _4899_/B sky130_fd_sc_hd__nor2_1
X_5698_ _7034_/Q _5966_/B1 _5697_/X _6986_/Q VGND VGND VPWR VPWR _5698_/X sky130_fd_sc_hd__a22o_1
XFILLER_147_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4649_ _4719_/A _4814_/B _4228_/Y VGND VGND VPWR VPWR _5031_/A sky130_fd_sc_hd__o21ai_1
XFILLER_190_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold740 _5492_/X VGND VGND VPWR VPWR _7057_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold751 _6926_/Q VGND VGND VPWR VPWR hold751/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold762 _4050_/X VGND VGND VPWR VPWR _6539_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold773 _6870_/Q VGND VGND VPWR VPWR hold773/X sky130_fd_sc_hd__dlygate4sd3_1
X_6319_ _6319_/A0 _6318_/X _6319_/S VGND VGND VPWR VPWR _7186_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold784 _4114_/X VGND VGND VPWR VPWR _6582_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold795 _7051_/Q VGND VGND VPWR VPWR hold795/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1440 _3471_/Y VGND VGND VPWR VPWR _4318_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1451 _6662_/Q VGND VGND VPWR VPWR hold1451/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1462 _6786_/Q VGND VGND VPWR VPWR _3603_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1473 _3330_/B VGND VGND VPWR VPWR _3299_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1484 _7168_/Q VGND VGND VPWR VPWR _5838_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_176_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1495 _6097_/X VGND VGND VPWR VPWR _7177_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3951_ input85/X input58/X _6460_/Q VGND VGND VPWR VPWR _3951_/X sky130_fd_sc_hd__mux2_2
XFILLER_50_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6670_ _6683_/CLK _6670_/D fanout511/X VGND VGND VPWR VPWR _6670_/Q sky130_fd_sc_hd__dfrtp_4
X_3882_ _4390_/A _4654_/A VGND VGND VPWR VPWR _4467_/A sky130_fd_sc_hd__and2_1
X_5621_ _7151_/Q _7150_/Q VGND VGND VPWR VPWR _5703_/B sky130_fd_sc_hd__nor2_2
X_5552_ _5552_/A0 hold500/X _5552_/S VGND VGND VPWR VPWR _5552_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4503_ _4502_/X _4887_/C _4503_/C _4503_/D VGND VGND VPWR VPWR _4503_/X sky130_fd_sc_hd__and4b_1
XFILLER_172_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5483_ hold40/X _5483_/A1 hold79/X VGND VGND VPWR VPWR hold80/A sky130_fd_sc_hd__mux2_1
XFILLER_144_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4434_ _4453_/A _4434_/B _4444_/B _4724_/A VGND VGND VPWR VPWR _4995_/A sky130_fd_sc_hd__or4_4
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7153_ _7182_/CLK _7153_/D fanout500/X VGND VGND VPWR VPWR _7153_/Q sky130_fd_sc_hd__dfstp_1
X_4365_ _4846_/A _4570_/B VGND VGND VPWR VPWR _4369_/B sky130_fd_sc_hd__nand2b_2
Xfanout505 fanout508/X VGND VGND VPWR VPWR fanout505/X sky130_fd_sc_hd__buf_8
Xfanout516 fanout517/X VGND VGND VPWR VPWR fanout516/X sky130_fd_sc_hd__buf_8
Xfanout527 input75/X VGND VGND VPWR VPWR fanout527/X sky130_fd_sc_hd__buf_12
X_6104_ _6933_/Q _6024_/B _6203_/A2 _6989_/Q _6103_/X VGND VGND VPWR VPWR _6109_/B
+ sky130_fd_sc_hd__a221o_1
X_3316_ _3546_/B _3334_/A VGND VGND VPWR VPWR _5394_/A sky130_fd_sc_hd__nor2_8
X_7084_ _7110_/CLK _7084_/D fanout508/X VGND VGND VPWR VPWR _7084_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_113_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4296_ _6394_/A0 _4296_/A1 _4299_/S VGND VGND VPWR VPWR _4296_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6035_ _6938_/Q _6024_/D wire394/X _6890_/Q _6034_/X VGND VGND VPWR VPWR _6044_/C
+ sky130_fd_sc_hd__a221o_1
X_3247_ _3971_/S hold93/X hold47/X VGND VGND VPWR VPWR hold48/A sky130_fd_sc_hd__o21bai_1
XFILLER_100_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_731 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6937_ _6977_/CLK _6937_/D fanout507/X VGND VGND VPWR VPWR _6937_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6868_ _7075_/CLK _6868_/D fanout514/X VGND VGND VPWR VPWR _6868_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_167_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5819_ _6960_/Q _5659_/X _5663_/X _7024_/Q VGND VGND VPWR VPWR _5819_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6799_ _7207_/CLK _6799_/D fanout484/X VGND VGND VPWR VPWR _6799_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_41_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold570 _5373_/X VGND VGND VPWR VPWR _6951_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold581 _7047_/Q VGND VGND VPWR VPWR hold581/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 _3987_/X VGND VGND VPWR VPWR _6485_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1270 _4253_/X VGND VGND VPWR VPWR _6706_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1281 _7042_/Q VGND VGND VPWR VPWR _5476_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1292 _4313_/X VGND VGND VPWR VPWR _6756_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4150_ _4327_/A1 hold807/X _4152_/S VGND VGND VPWR VPWR _4150_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4081_ hold193/X hold127/X _4085_/S VGND VGND VPWR VPWR _4081_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4983_ _4983_/A _4983_/B _4983_/C VGND VGND VPWR VPWR _4989_/C sky130_fd_sc_hd__nor3_1
XFILLER_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6722_ _6725_/CLK _6722_/D fanout509/X VGND VGND VPWR VPWR _6722_/Q sky130_fd_sc_hd__dfrtp_4
X_3934_ _3232_/Y _6443_/Q _6407_/B VGND VGND VPWR VPWR _3934_/X sky130_fd_sc_hd__mux2_8
XFILLER_189_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6653_ _7193_/CLK _6653_/D VGND VGND VPWR VPWR _6653_/Q sky130_fd_sc_hd__dfxtp_1
X_3865_ _3866_/A1 _3865_/A1 _3866_/S VGND VGND VPWR VPWR _6447_/D sky130_fd_sc_hd__mux2_1
X_5604_ _7144_/Q _7145_/Q _7146_/Q _5604_/D VGND VGND VPWR VPWR _5605_/A sky130_fd_sc_hd__and4_1
XFILLER_164_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3796_ _6472_/Q _6471_/Q _3801_/B VGND VGND VPWR VPWR _3800_/A sky130_fd_sc_hd__and3_1
X_6584_ _7130_/CLK _6584_/D fanout519/X VGND VGND VPWR VPWR _6584_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_191_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5535_ _5535_/A _5535_/B VGND VGND VPWR VPWR _5543_/S sky130_fd_sc_hd__and2_4
XFILLER_11_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5466_ _5466_/A _5535_/B VGND VGND VPWR VPWR _5474_/S sky130_fd_sc_hd__and2_4
XFILLER_145_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7205_ _3937_/A1 _7205_/D _6348_/B VGND VGND VPWR VPWR _7205_/Q sky130_fd_sc_hd__dfrtp_2
X_4417_ _4758_/A _5001_/A _4758_/B VGND VGND VPWR VPWR _4876_/A sky130_fd_sc_hd__and3_2
XFILLER_99_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5397_ hold819/X _5496_/A0 _5402_/S VGND VGND VPWR VPWR _5397_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7136_ _7136_/CLK hold6/X fanout519/X VGND VGND VPWR VPWR _7136_/Q sky130_fd_sc_hd__dfstp_2
X_4348_ _4348_/A _4348_/B _4348_/C VGND VGND VPWR VPWR _4542_/A sky130_fd_sc_hd__and3_1
XFILLER_98_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7067_ _7136_/CLK _7067_/D fanout521/X VGND VGND VPWR VPWR _7067_/Q sky130_fd_sc_hd__dfstp_2
X_4279_ hold44/X hold303/X _4281_/S VGND VGND VPWR VPWR _4279_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6018_ _6018_/A _6021_/A VGND VGND VPWR VPWR _6023_/D sky130_fd_sc_hd__nor2_8
XFILLER_55_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_240 hold36/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_251 _6613_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_262 input58/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3650_ _7076_/Q _5511_/A _3983_/A _6484_/Q _3649_/X VGND VGND VPWR VPWR _3651_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_9_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3581_ _6965_/Q _5385_/A _4104_/A input64/X _3580_/X VGND VGND VPWR VPWR _3582_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5320_ _5569_/A0 hold215/X hold23/X VGND VGND VPWR VPWR _5320_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5251_ _5251_/A0 _5536_/A1 _5258_/S VGND VGND VPWR VPWR _5251_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4202_ hold385/X _5533_/A1 _4203_/S VGND VGND VPWR VPWR _4202_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5182_ _6782_/Q _6362_/A _5156_/Y _5178_/X _5181_/Y VGND VGND VPWR VPWR _5183_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_142_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4133_ hold498/X _6396_/A0 _4134_/S VGND VGND VPWR VPWR _4133_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4064_ _4117_/A1 _5550_/A0 _4068_/S VGND VGND VPWR VPWR _4064_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4966_ _5016_/A _4694_/B _4758_/Y _4786_/Y VGND VGND VPWR VPWR _4969_/A sky130_fd_sc_hd__o211a_1
XFILLER_51_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6705_ _6755_/CLK _6705_/D fanout497/X VGND VGND VPWR VPWR _6705_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_189_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3917_ _3917_/A _3917_/B VGND VGND VPWR VPWR _6443_/D sky130_fd_sc_hd__and2_2
XFILLER_177_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4897_ _5158_/A _4897_/B _4897_/C _4530_/B VGND VGND VPWR VPWR _4897_/X sky130_fd_sc_hd__or4b_1
XFILLER_22_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6636_ _7094_/CLK _6636_/D fanout494/X VGND VGND VPWR VPWR _6636_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_165_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3848_ _6472_/Q _6471_/Q _6473_/Q VGND VGND VPWR VPWR _3848_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_165_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6567_ _6925_/CLK _6567_/D fanout516/X VGND VGND VPWR VPWR _6567_/Q sky130_fd_sc_hd__dfrtp_1
X_3779_ _7082_/Q _5520_/A _5403_/A _6978_/Q VGND VGND VPWR VPWR _3779_/X sky130_fd_sc_hd__a22o_2
XFILLER_164_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5518_ _5587_/A0 hold926/X _5519_/S VGND VGND VPWR VPWR _5518_/X sky130_fd_sc_hd__mux2_1
X_6498_ _7002_/CLK _6498_/D fanout498/X VGND VGND VPWR VPWR _6498_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_145_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5449_ _5536_/A1 _5449_/A1 _5456_/S VGND VGND VPWR VPWR _5449_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7119_ _7123_/CLK _7119_/D fanout527/X VGND VGND VPWR VPWR _7119_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_wbbd_sck clkbuf_0_wbbd_sck/X VGND VGND VPWR VPWR _3942_/A2 sky130_fd_sc_hd__clkbuf_16
XFILLER_179_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_506 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4820_ _4935_/A _4819_/C _4971_/B _4797_/A _4607_/X VGND VGND VPWR VPWR _4821_/D
+ sky130_fd_sc_hd__a41o_1
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4751_ _4994_/A _5036_/A VGND VGND VPWR VPWR _4987_/B sky130_fd_sc_hd__nor2_1
XFILLER_193_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3702_ _6491_/Q _3992_/A _4040_/A _6532_/Q VGND VGND VPWR VPWR _3702_/X sky130_fd_sc_hd__a22o_1
XFILLER_147_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4682_ _5023_/A _5023_/B _4582_/B VGND VGND VPWR VPWR _4699_/A sky130_fd_sc_hd__a21o_1
XFILLER_119_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6421_ _6441_/A _6440_/B VGND VGND VPWR VPWR _6421_/X sky130_fd_sc_hd__and2_1
X_3633_ _3633_/A _3633_/B _3633_/C _3633_/D VGND VGND VPWR VPWR _3660_/A sky130_fd_sc_hd__or4_2
XFILLER_174_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6352_ _6352_/A0 _3601_/X _6356_/S VGND VGND VPWR VPWR _7192_/D sky130_fd_sc_hd__mux2_1
X_3564_ _6917_/Q _5331_/A _3562_/X _3563_/X VGND VGND VPWR VPWR _3583_/B sky130_fd_sc_hd__a211o_1
XFILLER_108_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5303_ _5579_/A0 hold524/X _5303_/S VGND VGND VPWR VPWR _5303_/X sky130_fd_sc_hd__mux2_1
X_6283_ _6667_/Q wire412/X _6016_/X _6683_/Q VGND VGND VPWR VPWR _6283_/X sky130_fd_sc_hd__a22o_1
XFILLER_142_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3495_ _3495_/A _3528_/B VGND VGND VPWR VPWR _4028_/A sky130_fd_sc_hd__nor2_4
X_5234_ _5459_/A0 hold203/X _5240_/S VGND VGND VPWR VPWR _5234_/X sky130_fd_sc_hd__mux2_1
X_5165_ _4502_/A _5067_/A _5165_/C _5165_/D VGND VGND VPWR VPWR _5180_/C sky130_fd_sc_hd__and4bb_1
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4116_ hold85/X hold179/X hold97/X VGND VGND VPWR VPWR _4116_/X sky130_fd_sc_hd__mux2_1
X_5096_ _4993_/A _4870_/B _4971_/B _4778_/B VGND VGND VPWR VPWR _5096_/X sky130_fd_sc_hd__o31a_1
XFILLER_84_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4047_ _6393_/A0 _4047_/A1 _4051_/S VGND VGND VPWR VPWR _4047_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5998_ _6038_/A _6021_/B VGND VGND VPWR VPWR _5998_/Y sky130_fd_sc_hd__nor2_8
XFILLER_52_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4949_ _4932_/A _4933_/A _4944_/B _4932_/B _4837_/X VGND VGND VPWR VPWR _4950_/C
+ sky130_fd_sc_hd__o41a_1
XFILLER_33_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6619_ _6740_/CLK _6619_/D _3873_/A VGND VGND VPWR VPWR _6619_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_193_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput280 _6488_/Q VGND VGND VPWR VPWR pll_trim[14] sky130_fd_sc_hd__buf_12
Xoutput291 _6804_/Q VGND VGND VPWR VPWR pll_trim[24] sky130_fd_sc_hd__buf_12
XFILLER_121_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_615 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3280_ _5212_/B _3528_/A VGND VGND VPWR VPWR _3280_/Y sky130_fd_sc_hd__nor2_2
XFILLER_97_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6970_ _6970_/CLK _6970_/D fanout505/X VGND VGND VPWR VPWR _6970_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5921_ _6763_/Q _5686_/X _5705_/X _6683_/Q VGND VGND VPWR VPWR _5921_/X sky130_fd_sc_hd__a22o_1
XFILLER_80_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5852_ _7065_/Q _5671_/X _5693_/X _6905_/Q _5851_/X VGND VGND VPWR VPWR _5857_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_61_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4803_ _4674_/A _4569_/Y _4592_/Y _5049_/B VGND VGND VPWR VPWR _4817_/B sky130_fd_sc_hd__a31o_1
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5783_ _6974_/Q _5691_/B _5699_/X _7054_/Q _5690_/X VGND VGND VPWR VPWR _5783_/X
+ sky130_fd_sc_hd__a221o_1
X_4734_ _4872_/A _4802_/A VGND VGND VPWR VPWR _4770_/C sky130_fd_sc_hd__nor2_1
XFILLER_119_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4665_ _5021_/C _4665_/B VGND VGND VPWR VPWR _4665_/Y sky130_fd_sc_hd__nor2_1
XFILLER_190_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6404_ _6407_/A _6407_/B VGND VGND VPWR VPWR _6404_/X sky130_fd_sc_hd__and2_1
Xhold900 _6984_/Q VGND VGND VPWR VPWR hold900/X sky130_fd_sc_hd__dlygate4sd3_1
X_3616_ input58/X _4083_/S _5544_/A _7105_/Q VGND VGND VPWR VPWR _3616_/X sky130_fd_sc_hd__a22o_1
Xhold911 _5473_/X VGND VGND VPWR VPWR _7040_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold922 hold922/A VGND VGND VPWR VPWR hold922/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_134_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4596_ _4596_/A _4596_/B VGND VGND VPWR VPWR _4596_/X sky130_fd_sc_hd__or2_2
Xhold933 _4200_/X VGND VGND VPWR VPWR _6656_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6335_ _6540_/Q _5988_/X _6023_/C _6615_/Q VGND VGND VPWR VPWR _6335_/X sky130_fd_sc_hd__a22o_1
Xhold944 _6675_/Q VGND VGND VPWR VPWR hold944/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3547_ _5212_/B _3547_/B VGND VGND VPWR VPWR _3547_/Y sky130_fd_sc_hd__nor2_1
Xhold955 _4217_/X VGND VGND VPWR VPWR _6670_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold966 _6819_/Q VGND VGND VPWR VPWR _5221_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold977 hold977/A VGND VGND VPWR VPWR hold977/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold988 _5568_/X VGND VGND VPWR VPWR _7124_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6266_ _6266_/A _6266_/B _6266_/C _6266_/D VGND VGND VPWR VPWR _6267_/C sky130_fd_sc_hd__or4_1
X_3478_ _3530_/B _3729_/B VGND VGND VPWR VPWR _4246_/A sky130_fd_sc_hd__nor2_4
Xhold999 _7140_/Q VGND VGND VPWR VPWR hold999/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5217_ _5583_/A0 hold283/X _5220_/S VGND VGND VPWR VPWR _5217_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1600 _6572_/Q VGND VGND VPWR VPWR hold349/A sky130_fd_sc_hd__dlygate4sd3_1
X_6197_ _7134_/Q _6320_/A2 _6320_/B1 _6881_/Q VGND VGND VPWR VPWR _6197_/X sky130_fd_sc_hd__a22o_1
Xhold1611 _6716_/Q VGND VGND VPWR VPWR hold1611/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5148_ _5148_/A _5148_/B _5148_/C _5148_/D VGND VGND VPWR VPWR _5148_/Y sky130_fd_sc_hd__nor4_1
X_5079_ _5079_/A _5079_/B VGND VGND VPWR VPWR _5106_/C sky130_fd_sc_hd__or2_1
XFILLER_71_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4450_ _4570_/B _5035_/A VGND VGND VPWR VPWR _4657_/C sky130_fd_sc_hd__nor2_8
Xhold207 _7098_/Q VGND VGND VPWR VPWR hold207/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 _5253_/X VGND VGND VPWR VPWR _6844_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold229 _6553_/Q VGND VGND VPWR VPWR hold229/X sky130_fd_sc_hd__dlygate4sd3_1
X_3401_ _7064_/Q _5493_/A _5322_/A _6912_/Q VGND VGND VPWR VPWR _3401_/X sky130_fd_sc_hd__a22o_1
XFILLER_132_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4381_ _4657_/A _4999_/A VGND VGND VPWR VPWR _4719_/A sky130_fd_sc_hd__nand2_1
XFILLER_98_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3332_ hold29/X _3534_/A VGND VGND VPWR VPWR _5430_/A sky130_fd_sc_hd__nor2_8
X_6120_ _6845_/Q _6046_/B _6110_/X _6119_/X _3195_/Y VGND VGND VPWR VPWR _6120_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_171_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3263_ hold54/X _4929_/A1 _3971_/S VGND VGND VPWR VPWR hold55/A sky130_fd_sc_hd__mux2_4
X_6051_ _7083_/Q _5977_/X _6323_/B1 _7120_/Q VGND VGND VPWR VPWR _6051_/X sky130_fd_sc_hd__a22o_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _5002_/A _5036_/B VGND VGND VPWR VPWR _5049_/D sky130_fd_sc_hd__nor2_1
XFILLER_85_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3194_ _6565_/Q VGND VGND VPWR VPWR _5648_/C sky130_fd_sc_hd__inv_2
XFILLER_39_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6953_ _6992_/CLK _6953_/D fanout517/X VGND VGND VPWR VPWR _6953_/Q sky130_fd_sc_hd__dfrtp_1
X_5904_ _5904_/A0 _5903_/X _6319_/S VGND VGND VPWR VPWR _7171_/D sky130_fd_sc_hd__mux2_1
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6884_ _7136_/CLK _6884_/D fanout520/X VGND VGND VPWR VPWR _6884_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_62_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5835_ _5835_/A _5835_/B _5835_/C _5835_/D VGND VGND VPWR VPWR _5835_/X sky130_fd_sc_hd__or4_1
XFILLER_61_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5766_ _6949_/Q _5666_/X _5685_/X _6909_/Q _5765_/X VGND VGND VPWR VPWR _5770_/B
+ sky130_fd_sc_hd__a221o_1
X_4717_ _4745_/A _5035_/B VGND VGND VPWR VPWR _5050_/B sky130_fd_sc_hd__or2_1
XFILLER_148_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5697_ _7152_/Q _5703_/B _5699_/B VGND VGND VPWR VPWR _5697_/X sky130_fd_sc_hd__and3_4
XFILLER_108_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4648_ _4963_/A _4648_/B VGND VGND VPWR VPWR _4648_/Y sky130_fd_sc_hd__nor2_1
XFILLER_107_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold730 _5543_/X VGND VGND VPWR VPWR _7102_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold741 _6509_/Q VGND VGND VPWR VPWR hold741/X sky130_fd_sc_hd__dlygate4sd3_1
X_4579_ _4814_/A _5016_/A VGND VGND VPWR VPWR _4639_/A sky130_fd_sc_hd__or2_4
Xhold752 _5345_/X VGND VGND VPWR VPWR _6926_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 _6958_/Q VGND VGND VPWR VPWR hold763/X sky130_fd_sc_hd__dlygate4sd3_1
X_6318_ _6318_/A0 _6317_/X _6318_/S VGND VGND VPWR VPWR _6318_/X sky130_fd_sc_hd__mux2_1
Xhold774 _5282_/X VGND VGND VPWR VPWR _6870_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold785 _6720_/Q VGND VGND VPWR VPWR hold785/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold796 _5486_/X VGND VGND VPWR VPWR _7051_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6249_ _6537_/Q _5988_/X _6022_/B _6656_/Q VGND VGND VPWR VPWR _6249_/X sky130_fd_sc_hd__a22o_1
XFILLER_77_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1430 _7034_/Q VGND VGND VPWR VPWR hold1430/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1441 _4321_/X VGND VGND VPWR VPWR _6763_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1452 _4207_/X VGND VGND VPWR VPWR _6662_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1463 _3603_/X VGND VGND VPWR VPWR _6786_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1474 _6627_/Q VGND VGND VPWR VPWR _4167_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1485 _5838_/X VGND VGND VPWR VPWR _7168_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_61_csclk _6753_/CLK VGND VGND VPWR VPWR _7002_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1496 _7163_/Q VGND VGND VPWR VPWR _5731_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_55_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_76_csclk _6753_/CLK VGND VGND VPWR VPWR _7207_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_14_csclk _6882_/CLK VGND VGND VPWR VPWR _6579_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_96_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold90 hold90/A VGND VGND VPWR VPWR hold90/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_29_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7138_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_90_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3950_ _3950_/A VGND VGND VPWR VPWR _3950_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3881_ _4338_/C _4338_/D _4337_/A _4337_/B VGND VGND VPWR VPWR _3887_/C sky130_fd_sc_hd__or4_1
X_5620_ _5620_/A1 _5618_/B _5624_/B _5619_/Y VGND VGND VPWR VPWR _7150_/D sky130_fd_sc_hd__a31o_1
XFILLER_188_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5551_ _5578_/A0 hold860/X _5552_/S VGND VGND VPWR VPWR _5551_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4502_ _4502_/A _5053_/A _5165_/D VGND VGND VPWR VPWR _4502_/X sky130_fd_sc_hd__or3b_1
X_5482_ _5587_/A0 hold886/X hold79/X VGND VGND VPWR VPWR _5482_/X sky130_fd_sc_hd__mux2_1
X_4433_ _4758_/A _4436_/B _4433_/C _4758_/B VGND VGND VPWR VPWR _4759_/B sky130_fd_sc_hd__and4_2
XFILLER_144_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7152_ _7183_/CLK _7152_/D fanout500/X VGND VGND VPWR VPWR _7152_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_116_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4364_ _4474_/A _4489_/A VGND VGND VPWR VPWR _4745_/A sky130_fd_sc_hd__or2_4
Xfanout506 fanout508/X VGND VGND VPWR VPWR fanout506/X sky130_fd_sc_hd__buf_8
Xfanout517 fanout526/X VGND VGND VPWR VPWR fanout517/X sky130_fd_sc_hd__buf_8
X_6103_ _6901_/Q _6022_/B _6212_/B1 _7045_/Q VGND VGND VPWR VPWR _6103_/X sky130_fd_sc_hd__a22o_1
X_3315_ _3534_/A hold68/X VGND VGND VPWR VPWR _5439_/A sky130_fd_sc_hd__nor2_8
XFILLER_112_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout528 fanout529/X VGND VGND VPWR VPWR _6348_/B sky130_fd_sc_hd__buf_6
X_4295_ _6393_/A0 _4295_/A1 _4299_/S VGND VGND VPWR VPWR _4295_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7083_ _7139_/CLK _7083_/D fanout518/X VGND VGND VPWR VPWR _7083_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_113_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3246_ hold46/X _3971_/S _3244_/X _3245_/Y VGND VGND VPWR VPWR hold47/A sky130_fd_sc_hd__o31a_1
XFILLER_100_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6034_ _6914_/Q wire412/X _6205_/B1 _7058_/Q VGND VGND VPWR VPWR _6034_/X sky130_fd_sc_hd__a22o_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6936_ _6977_/CLK _6936_/D fanout507/X VGND VGND VPWR VPWR _6936_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6867_ _7043_/CLK _6867_/D fanout514/X VGND VGND VPWR VPWR _6867_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_179_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5818_ _6880_/Q _5667_/X _5682_/X _7088_/Q _5817_/X VGND VGND VPWR VPWR _5825_/A
+ sky130_fd_sc_hd__a221o_1
X_6798_ _7207_/CLK _6798_/D fanout484/X VGND VGND VPWR VPWR _6798_/Q sky130_fd_sc_hd__dfrtp_2
X_5749_ _6996_/Q _5656_/X _5694_/X _7076_/Q _5748_/X VGND VGND VPWR VPWR _5750_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_136_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold560 _6515_/Q VGND VGND VPWR VPWR hold560/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold571 _6725_/Q VGND VGND VPWR VPWR hold571/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold582 _5481_/X VGND VGND VPWR VPWR _7047_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_173_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold593 _6801_/Q VGND VGND VPWR VPWR hold593/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_173_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1260 _5449_/X VGND VGND VPWR VPWR _7018_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1271 _6655_/Q VGND VGND VPWR VPWR _4199_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1282 _5476_/X VGND VGND VPWR VPWR _7042_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1293 _6490_/Q VGND VGND VPWR VPWR _3993_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4080_ hold417/X _4079_/X _4086_/S VGND VGND VPWR VPWR _4080_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4982_ _4982_/A _4982_/B _4982_/C VGND VGND VPWR VPWR _5119_/B sky130_fd_sc_hd__or3_1
X_6721_ _6725_/CLK _6721_/D fanout509/X VGND VGND VPWR VPWR _6721_/Q sky130_fd_sc_hd__dfrtp_4
X_3933_ _6554_/Q input3/X input1/X VGND VGND VPWR VPWR _3933_/X sky130_fd_sc_hd__mux2_4
X_6652_ _7193_/CLK _6652_/D VGND VGND VPWR VPWR _6652_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3864_ _3865_/A1 _3864_/A1 _3866_/S VGND VGND VPWR VPWR _6448_/D sky130_fd_sc_hd__mux2_1
X_5603_ _7144_/Q _7145_/Q _5604_/D _7146_/Q VGND VGND VPWR VPWR _5606_/B sky130_fd_sc_hd__a31o_1
XFILLER_118_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6583_ _7142_/CLK _6583_/D fanout525/X VGND VGND VPWR VPWR _6583_/Q sky130_fd_sc_hd__dfrtp_1
X_3795_ _3801_/B VGND VGND VPWR VPWR _3795_/Y sky130_fd_sc_hd__inv_2
X_5534_ hold695/X _5534_/A1 _5534_/S VGND VGND VPWR VPWR _5534_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5465_ _5552_/A0 hold745/X _5465_/S VGND VGND VPWR VPWR _5465_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7204_ _3937_/A1 _7204_/D fanout529/X VGND VGND VPWR VPWR _7204_/Q sky130_fd_sc_hd__dfrtp_1
X_4416_ _4434_/B _4444_/B VGND VGND VPWR VPWR _4758_/B sky130_fd_sc_hd__nor2_4
X_5396_ hold848/X _5573_/A0 _5402_/S VGND VGND VPWR VPWR _5396_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7135_ _7135_/CLK _7135_/D fanout519/X VGND VGND VPWR VPWR _7135_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_160_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4347_ _4935_/A _4819_/C _4781_/A VGND VGND VPWR VPWR _4350_/B sky130_fd_sc_hd__and3_1
XFILLER_113_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7066_ _7123_/CLK _7066_/D _6407_/A VGND VGND VPWR VPWR _7066_/Q sky130_fd_sc_hd__dfstp_4
X_4278_ _5459_/A0 hold343/X _4281_/S VGND VGND VPWR VPWR _4278_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6017_ _6019_/A _6033_/A _6030_/C VGND VGND VPWR VPWR _6022_/D sky130_fd_sc_hd__and3b_4
X_3229_ _6885_/Q VGND VGND VPWR VPWR _3229_/Y sky130_fd_sc_hd__clkinv_2
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f_wbbd_sck clkbuf_0_wbbd_sck/X VGND VGND VPWR VPWR _6387_/A1 sky130_fd_sc_hd__clkbuf_16
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6919_ _7108_/CLK _6919_/D fanout523/X VGND VGND VPWR VPWR _6919_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold390 _5447_/X VGND VGND VPWR VPWR _7017_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1090 _6660_/Q VGND VGND VPWR VPWR _4205_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_230 _5569_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_241 hold79/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_252 _7214_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_263 _5581_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3580_ _6619_/Q _4153_/A hold50/A _6678_/Q VGND VGND VPWR VPWR _3580_/X sky130_fd_sc_hd__a22o_2
XFILLER_139_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5250_ _5250_/A _5535_/B VGND VGND VPWR VPWR _5258_/S sky130_fd_sc_hd__and2_4
XFILLER_142_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4201_ hold827/X _4327_/A1 _4203_/S VGND VGND VPWR VPWR _4201_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5181_ _5123_/X _5180_/X _5160_/X VGND VGND VPWR VPWR _5181_/Y sky130_fd_sc_hd__a21oi_2
X_4132_ _4132_/A0 _6395_/A0 _4134_/S VGND VGND VPWR VPWR _4132_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4063_ hold381/X _4062_/X _4069_/S VGND VGND VPWR VPWR _4063_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4965_ _4965_/A _4965_/B _4816_/X VGND VGND VPWR VPWR _5142_/A sky130_fd_sc_hd__or3b_1
XFILLER_51_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6704_ _6708_/CLK _6704_/D fanout496/X VGND VGND VPWR VPWR _6704_/Q sky130_fd_sc_hd__dfrtp_2
X_3916_ _6542_/Q _6545_/Q _3850_/B VGND VGND VPWR VPWR _3917_/B sky130_fd_sc_hd__o21ai_1
XFILLER_149_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4896_ _5134_/A _4896_/B _4896_/C _5045_/A VGND VGND VPWR VPWR _4897_/B sky130_fd_sc_hd__or4_1
X_6635_ _7093_/CLK _6635_/D _6432_/A VGND VGND VPWR VPWR _6635_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3847_ input58/X _3847_/A1 _3847_/S VGND VGND VPWR VPWR _6456_/D sky130_fd_sc_hd__mux2_1
XFILLER_137_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6566_ _6925_/CLK _6566_/D fanout516/X VGND VGND VPWR VPWR _6566_/Q sky130_fd_sc_hd__dfrtp_1
X_3778_ _6498_/Q _3778_/A2 _5484_/A _7050_/Q _3777_/X VGND VGND VPWR VPWR _3781_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_152_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5517_ _5550_/A0 hold599/X _5519_/S VGND VGND VPWR VPWR _5517_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6497_ _6760_/CLK _6497_/D fanout488/X VGND VGND VPWR VPWR _6497_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_106_726 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5448_ _5448_/A _5535_/B VGND VGND VPWR VPWR _5456_/S sky130_fd_sc_hd__nand2_8
XFILLER_160_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5379_ _5574_/A0 _5379_/A1 _5384_/S VGND VGND VPWR VPWR _5379_/X sky130_fd_sc_hd__mux2_1
X_7118_ _7132_/CLK _7118_/D fanout525/X VGND VGND VPWR VPWR _7118_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7049_ _7049_/CLK hold80/X fanout522/X VGND VGND VPWR VPWR _7049_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4750_ _5002_/A _5036_/A VGND VGND VPWR VPWR _4983_/B sky130_fd_sc_hd__nor2_1
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3701_ _3701_/A _3701_/B _3701_/C _3701_/D VGND VGND VPWR VPWR _3722_/B sky130_fd_sc_hd__or4_1
XFILLER_186_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4681_ _4832_/B _5024_/A _5017_/A _5076_/A VGND VGND VPWR VPWR _4681_/X sky130_fd_sc_hd__o22a_1
XFILLER_159_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6420_ _6441_/A _6440_/B VGND VGND VPWR VPWR _6420_/X sky130_fd_sc_hd__and2_1
X_3632_ _3632_/A _3632_/B _3632_/C _3632_/D VGND VGND VPWR VPWR _3633_/D sky130_fd_sc_hd__or4_1
XFILLER_134_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6351_ _6351_/A0 _3660_/X _6356_/S VGND VGND VPWR VPWR _7191_/D sky130_fd_sc_hd__mux2_1
X_3563_ _6668_/Q _4210_/A _4198_/A _6658_/Q _3549_/X VGND VGND VPWR VPWR _3563_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_127_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5302_ _5578_/A0 hold825/X _5303_/S VGND VGND VPWR VPWR _5302_/X sky130_fd_sc_hd__mux2_1
X_6282_ _6748_/Q _6322_/B1 _6030_/X _6743_/Q _6281_/X VGND VGND VPWR VPWR _6292_/B
+ sky130_fd_sc_hd__a221o_1
X_3494_ input56/X _5232_/A _3340_/Y input24/X _3493_/X VGND VGND VPWR VPWR _3499_/C
+ sky130_fd_sc_hd__a221o_2
XFILLER_88_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5233_ _5581_/A0 hold971/X _5240_/S VGND VGND VPWR VPWR _5233_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5164_ _4932_/A _4784_/A _5016_/B _4950_/C VGND VGND VPWR VPWR _5165_/C sky130_fd_sc_hd__o31a_1
XFILLER_111_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4115_ _5584_/A0 hold472/X hold97/X VGND VGND VPWR VPWR _4115_/X sky130_fd_sc_hd__mux2_1
X_5095_ _5095_/A _5095_/B _5095_/C _5095_/D VGND VGND VPWR VPWR _5145_/B sky130_fd_sc_hd__or4_1
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4046_ _4046_/A _6392_/B VGND VGND VPWR VPWR _4051_/S sky130_fd_sc_hd__nand2_2
XFILLER_17_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5997_ _6038_/A _6019_/B VGND VGND VPWR VPWR _5997_/Y sky130_fd_sc_hd__nor2_8
XFILLER_52_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4948_ _4932_/A _4947_/A _4933_/A _4932_/B _4857_/A VGND VGND VPWR VPWR _4950_/B
+ sky130_fd_sc_hd__o41a_1
X_4879_ _4996_/A _5036_/A _4510_/B VGND VGND VPWR VPWR _5174_/A sky130_fd_sc_hd__o21ai_1
XFILLER_138_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6618_ _6963_/CLK _6618_/D fanout509/X VGND VGND VPWR VPWR _6618_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_192_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6549_ _7142_/CLK _6549_/D fanout525/X VGND VGND VPWR VPWR _6549_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput270 _6797_/Q VGND VGND VPWR VPWR pll_div[4] sky130_fd_sc_hd__buf_12
Xoutput281 _6489_/Q VGND VGND VPWR VPWR pll_trim[15] sky130_fd_sc_hd__buf_12
XFILLER_121_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput292 _6805_/Q VGND VGND VPWR VPWR pll_trim[25] sky130_fd_sc_hd__buf_12
XFILLER_121_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5920_ _6533_/Q _5678_/X _5702_/X _6723_/Q _5919_/X VGND VGND VPWR VPWR _5923_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5851_ _6913_/Q _5685_/X _5691_/B _5850_/X VGND VGND VPWR VPWR _5851_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4802_ _4802_/A _4802_/B _4802_/C _4802_/D VGND VGND VPWR VPWR _4822_/C sky130_fd_sc_hd__nor4_1
X_5782_ _6982_/Q _5702_/X _5706_/X _6502_/Q _5781_/X VGND VGND VPWR VPWR _5785_/C
+ sky130_fd_sc_hd__a221o_1
X_4733_ _4656_/Y _4667_/X _5039_/A _4758_/A VGND VGND VPWR VPWR _4761_/A sky130_fd_sc_hd__o22a_1
XFILLER_159_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4664_ _4664_/A _4814_/B VGND VGND VPWR VPWR _4665_/B sky130_fd_sc_hd__or2_1
XFILLER_174_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6403_ _6407_/A _6407_/B VGND VGND VPWR VPWR _6403_/X sky130_fd_sc_hd__and2_1
X_3615_ _6932_/Q _5349_/A _3320_/Y _6956_/Q VGND VGND VPWR VPWR _3615_/X sky130_fd_sc_hd__a22o_1
XFILLER_135_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold901 _5410_/X VGND VGND VPWR VPWR _6984_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4595_ _4674_/A _4595_/B VGND VGND VPWR VPWR _4659_/B sky130_fd_sc_hd__nand2_8
Xhold912 _7091_/Q VGND VGND VPWR VPWR hold912/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold923 _4122_/X VGND VGND VPWR VPWR _6589_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold934 _6507_/Q VGND VGND VPWR VPWR hold934/X sky130_fd_sc_hd__dlygate4sd3_1
X_6334_ _6515_/Q _5977_/X _5997_/Y _6735_/Q _6333_/X VGND VGND VPWR VPWR _6341_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_162_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3546_ _3546_/A _3546_/B VGND VGND VPWR VPWR _5205_/A sky130_fd_sc_hd__nor2_8
Xhold945 _4223_/X VGND VGND VPWR VPWR _6675_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold956 _6551_/Q VGND VGND VPWR VPWR hold956/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold967 _5221_/X VGND VGND VPWR VPWR hold967/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold978 _4121_/X VGND VGND VPWR VPWR _6588_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6265_ _6612_/Q _6023_/C _6020_/X _6707_/Q _6249_/X VGND VGND VPWR VPWR _6266_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold989 _6935_/Q VGND VGND VPWR VPWR hold989/X sky130_fd_sc_hd__dlygate4sd3_1
X_3477_ hold49/X _3525_/B VGND VGND VPWR VPWR _4216_/A sky130_fd_sc_hd__nor2_4
XFILLER_115_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5216_ _5539_/A1 hold231/X _5220_/S VGND VGND VPWR VPWR _5216_/X sky130_fd_sc_hd__mux2_1
X_6196_ _6196_/A1 _5652_/Y _6194_/X _6195_/X VGND VGND VPWR VPWR _7181_/D sky130_fd_sc_hd__a22o_1
XFILLER_130_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1601 _7107_/Q VGND VGND VPWR VPWR hold653/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1612 _6767_/Q VGND VGND VPWR VPWR hold301/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5147_ _5172_/B _5147_/B VGND VGND VPWR VPWR _5147_/X sky130_fd_sc_hd__and2b_1
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5078_ _4659_/B _5108_/B _5077_/X VGND VGND VPWR VPWR _5178_/A sky130_fd_sc_hd__o21ai_1
XFILLER_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4029_ _4029_/A0 _5476_/A0 _4033_/S VGND VGND VPWR VPWR _4029_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold208 _5539_/X VGND VGND VPWR VPWR _7098_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold219 _6618_/Q VGND VGND VPWR VPWR hold219/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3400_ _6896_/Q _5304_/A _3397_/X _3399_/X VGND VGND VPWR VPWR _3409_/C sky130_fd_sc_hd__a211o_1
XFILLER_125_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4380_ _4588_/A _4935_/A _4605_/A _4621_/B VGND VGND VPWR VPWR _5021_/A sky130_fd_sc_hd__or4_4
XFILLER_98_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3331_ _3536_/A hold76/X VGND VGND VPWR VPWR hold77/A sky130_fd_sc_hd__nor2_8
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6050_ _7136_/Q _6308_/A2 _6338_/B1 _7096_/Q VGND VGND VPWR VPWR _6050_/X sky130_fd_sc_hd__a22o_1
XFILLER_112_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ hold53/X hold25/X hold72/A VGND VGND VPWR VPWR hold54/A sky130_fd_sc_hd__mux2_1
XFILLER_140_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5001_ _5001_/A _5001_/B _5001_/C VGND VGND VPWR VPWR _5042_/C sky130_fd_sc_hd__and3_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3193_ _3193_/A VGND VGND VPWR VPWR _5615_/A sky130_fd_sc_hd__inv_2
XFILLER_66_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6952_ _7031_/CLK _6952_/D fanout517/X VGND VGND VPWR VPWR _6952_/Q sky130_fd_sc_hd__dfrtp_4
X_5903_ _6563_/Q _7170_/Q _5902_/X VGND VGND VPWR VPWR _5903_/X sky130_fd_sc_hd__a21o_1
XFILLER_179_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6883_ _6883_/CLK _6883_/D fanout505/X VGND VGND VPWR VPWR _6883_/Q sky130_fd_sc_hd__dfstp_1
X_5834_ _6992_/Q _5697_/X _5700_/X _7032_/Q _5833_/X VGND VGND VPWR VPWR _5835_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_179_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5765_ _6957_/Q _5659_/X _5705_/X _6941_/Q VGND VGND VPWR VPWR _5765_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4716_ _4745_/A _5035_/B VGND VGND VPWR VPWR _5031_/B sky130_fd_sc_hd__nor2_1
X_5696_ _7152_/Q _5705_/B _5699_/C VGND VGND VPWR VPWR _5696_/X sky130_fd_sc_hd__and3_4
XFILLER_163_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4647_ _4647_/A _4647_/B VGND VGND VPWR VPWR _4648_/B sky130_fd_sc_hd__nor2_1
XFILLER_162_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold720 _4310_/X VGND VGND VPWR VPWR _6754_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold731 _6854_/Q VGND VGND VPWR VPWR hold731/X sky130_fd_sc_hd__dlygate4sd3_1
X_4578_ _4588_/A _4605_/A _4621_/B _4935_/A VGND VGND VPWR VPWR _4646_/A sky130_fd_sc_hd__or4b_4
Xhold742 _4014_/X VGND VGND VPWR VPWR _6509_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold753 _6519_/Q VGND VGND VPWR VPWR hold753/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6317_ _6301_/X _6307_/X _6316_/X _6046_/B _6599_/Q VGND VGND VPWR VPWR _6317_/X
+ sky130_fd_sc_hd__o32a_1
Xhold764 _5381_/X VGND VGND VPWR VPWR _6958_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3529_ _6894_/Q _3280_/Y _4159_/A _6625_/Q _3527_/X VGND VGND VPWR VPWR _3541_/A
+ sky130_fd_sc_hd__a221o_1
Xhold775 _6874_/Q VGND VGND VPWR VPWR hold775/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold786 _4269_/X VGND VGND VPWR VPWR _6720_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold797 _7011_/Q VGND VGND VPWR VPWR hold797/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6248_ _6532_/Q _6272_/B VGND VGND VPWR VPWR _6248_/X sky130_fd_sc_hd__and2_1
XFILLER_77_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6179_ _6928_/Q _6027_/B _6023_/D _6896_/Q _6178_/X VGND VGND VPWR VPWR _6180_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1420 _6626_/Q VGND VGND VPWR VPWR _4166_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1431 _5467_/X VGND VGND VPWR VPWR _7034_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1442 _6592_/Q VGND VGND VPWR VPWR hold209/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1453 _7058_/Q VGND VGND VPWR VPWR hold1453/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1464 _6785_/Q VGND VGND VPWR VPWR _3662_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1475 _6790_/Q VGND VGND VPWR VPWR _3376_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1486 _7162_/Q VGND VGND VPWR VPWR _5710_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1497 _5731_/X VGND VGND VPWR VPWR _7163_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_730 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold80 hold80/A VGND VGND VPWR VPWR hold80/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 hold91/A VGND VGND VPWR VPWR hold91/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_36_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3880_ _4337_/C _4337_/D _3880_/C input116/X VGND VGND VPWR VPWR _3887_/B sky130_fd_sc_hd__or4b_1
XFILLER_149_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5550_ _5550_/A0 hold423/X _5552_/S VGND VGND VPWR VPWR _5550_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4501_ _4489_/A _4981_/B _4932_/A _4500_/X VGND VGND VPWR VPWR _5053_/A sky130_fd_sc_hd__o31ai_1
X_5481_ _5550_/A0 hold581/X hold79/X VGND VGND VPWR VPWR _5481_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4432_ _4436_/B _4433_/C VGND VGND VPWR VPWR _4724_/A sky130_fd_sc_hd__nand2_1
X_7151_ _7183_/CLK _7151_/D fanout500/X VGND VGND VPWR VPWR _7151_/Q sky130_fd_sc_hd__dfrtp_1
X_4363_ _4944_/A _4428_/B _4426_/B VGND VGND VPWR VPWR _4489_/A sky130_fd_sc_hd__or3_1
XFILLER_98_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout507 fanout508/X VGND VGND VPWR VPWR fanout507/X sky130_fd_sc_hd__clkbuf_8
X_6102_ _7114_/Q _6322_/B1 _6206_/B1 _6981_/Q _6101_/X VGND VGND VPWR VPWR _6109_/A
+ sky130_fd_sc_hd__a221o_1
X_3314_ _3731_/A _4120_/B VGND VGND VPWR VPWR _3992_/A sky130_fd_sc_hd__nor2_8
XFILLER_140_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout518 fanout526/X VGND VGND VPWR VPWR fanout518/X sky130_fd_sc_hd__buf_8
Xfanout529 input164/X VGND VGND VPWR VPWR fanout529/X sky130_fd_sc_hd__buf_6
X_7082_ _7082_/CLK _7082_/D fanout527/X VGND VGND VPWR VPWR _7082_/Q sky130_fd_sc_hd__dfstp_2
X_4294_ _4294_/A _6392_/B VGND VGND VPWR VPWR _4299_/S sky130_fd_sc_hd__nand2_2
XFILLER_98_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6033_ _6033_/A _6040_/B _6040_/C VGND VGND VPWR VPWR _6033_/X sky130_fd_sc_hd__and3_4
X_3245_ _6782_/Q _3971_/S VGND VGND VPWR VPWR _3245_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_67_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_560 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6935_ _7134_/CLK _6935_/D fanout524/X VGND VGND VPWR VPWR _6935_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_35_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6866_ _7107_/CLK _6866_/D fanout511/X VGND VGND VPWR VPWR _6866_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5817_ _6904_/Q _5693_/X _5699_/X _7056_/Q VGND VGND VPWR VPWR _5817_/X sky130_fd_sc_hd__a22o_1
X_6797_ _7207_/CLK _6797_/D fanout484/X VGND VGND VPWR VPWR _6797_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_167_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5748_ _6956_/Q _5659_/X _5682_/X _7084_/Q VGND VGND VPWR VPWR _5748_/X sky130_fd_sc_hd__a22o_1
XFILLER_157_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5679_ _6914_/Q _5677_/X _5678_/X _7066_/Q VGND VGND VPWR VPWR _5679_/X sky130_fd_sc_hd__a22o_1
XFILLER_135_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold550 _6556_/Q VGND VGND VPWR VPWR hold550/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 _4021_/X VGND VGND VPWR VPWR _6515_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold572 _4275_/X VGND VGND VPWR VPWR _6725_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 _6497_/Q VGND VGND VPWR VPWR hold583/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold594 _5197_/X VGND VGND VPWR VPWR _6801_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1250 _6711_/Q VGND VGND VPWR VPWR _4259_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1261 _6906_/Q VGND VGND VPWR VPWR _5323_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1272 _4199_/X VGND VGND VPWR VPWR _6655_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1283 _6766_/Q VGND VGND VPWR VPWR _4325_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1294 _3993_/X VGND VGND VPWR VPWR _6490_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_696 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput170 wb_we_i VGND VGND VPWR VPWR _6358_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4981_ _5021_/A _4981_/B _4981_/C VGND VGND VPWR VPWR _4982_/C sky130_fd_sc_hd__nor3_1
XFILLER_23_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3932_ _3931_/X _3953_/B _6459_/Q VGND VGND VPWR VPWR _3932_/X sky130_fd_sc_hd__mux2_4
X_6720_ _7115_/CLK _6720_/D fanout501/X VGND VGND VPWR VPWR _6720_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_16_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6651_ _7193_/CLK _6651_/D VGND VGND VPWR VPWR _6651_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3863_ _3864_/A1 hold83/A _3866_/S VGND VGND VPWR VPWR _6449_/D sky130_fd_sc_hd__mux2_1
XFILLER_149_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5602_ _7145_/Q _5595_/Y _5600_/Y _5601_/X VGND VGND VPWR VPWR _7145_/D sky130_fd_sc_hd__a22o_1
X_6582_ _7142_/CLK _6582_/D fanout525/X VGND VGND VPWR VPWR _6582_/Q sky130_fd_sc_hd__dfrtp_1
X_3794_ _6541_/Q _3794_/B VGND VGND VPWR VPWR _3801_/B sky130_fd_sc_hd__or2_2
XFILLER_176_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5533_ hold791/X _5533_/A1 _5534_/S VGND VGND VPWR VPWR _5533_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5464_ _5587_/A0 hold882/X _5465_/S VGND VGND VPWR VPWR _5464_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_60_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7050_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_133_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7203_ _3937_/A1 _7203_/D fanout529/X VGND VGND VPWR VPWR hold99/A sky130_fd_sc_hd__dfrtp_1
X_4415_ _4415_/A _4435_/B VGND VGND VPWR VPWR _4444_/B sky130_fd_sc_hd__or2_2
X_5395_ _5395_/A0 _5536_/A1 _5402_/S VGND VGND VPWR VPWR _5395_/X sky130_fd_sc_hd__mux2_1
X_7134_ _7134_/CLK _7134_/D fanout524/X VGND VGND VPWR VPWR _7134_/Q sky130_fd_sc_hd__dfrtp_1
X_4346_ _4819_/C _4781_/A VGND VGND VPWR VPWR _4354_/A sky130_fd_sc_hd__nand2_1
XFILLER_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_75_csclk _6753_/CLK VGND VGND VPWR VPWR _7211_/CLK sky130_fd_sc_hd__clkbuf_16
X_7065_ _7065_/CLK _7065_/D fanout517/X VGND VGND VPWR VPWR _7065_/Q sky130_fd_sc_hd__dfrtp_2
X_4277_ _5581_/A0 _4277_/A1 _4281_/S VGND VGND VPWR VPWR _4277_/X sky130_fd_sc_hd__mux2_1
X_6016_ _6039_/A _6039_/C _6020_/C VGND VGND VPWR VPWR _6016_/X sky130_fd_sc_hd__and3_4
X_3228_ _6893_/Q VGND VGND VPWR VPWR _3228_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6918_ _7123_/CLK _6918_/D _6407_/A VGND VGND VPWR VPWR _6918_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_70_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6849_ _7098_/CLK _6849_/D fanout506/X VGND VGND VPWR VPWR _6849_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_168_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_28_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7136_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_136_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold380 _4097_/X VGND VGND VPWR VPWR _6570_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold391 _6808_/Q VGND VGND VPWR VPWR hold391/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1080 _5231_/X VGND VGND VPWR VPWR _6825_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1091 _4205_/X VGND VGND VPWR VPWR _6660_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_220 _6489_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_231 _5558_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_242 hold127/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_253 input58/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_264 _5581_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4200_ hold932/X _5531_/A1 _4203_/S VGND VGND VPWR VPWR _4200_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5180_ _4939_/C _5066_/C _5180_/C _5180_/D VGND VGND VPWR VPWR _5180_/X sky130_fd_sc_hd__and4bb_1
XFILLER_3_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4131_ _4131_/A0 _6394_/A0 _4134_/S VGND VGND VPWR VPWR _4131_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4062_ hold179/X hold85/X _4068_/S VGND VGND VPWR VPWR _4062_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4964_ _4964_/A _5112_/B VGND VGND VPWR VPWR _5103_/A sky130_fd_sc_hd__or2_1
X_6703_ _6755_/CLK _6703_/D fanout497/X VGND VGND VPWR VPWR _6703_/Q sky130_fd_sc_hd__dfstp_1
X_3915_ _3850_/B _3890_/Y _3834_/B hold72/A VGND VGND VPWR VPWR _6543_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_189_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4895_ _4742_/A _4742_/C _4741_/C _4741_/X VGND VGND VPWR VPWR _5045_/A sky130_fd_sc_hd__a31o_1
X_3846_ _6473_/Q _6472_/Q _6471_/Q _6541_/Q VGND VGND VPWR VPWR _3847_/S sky130_fd_sc_hd__or4bb_1
X_6634_ _7094_/CLK _6634_/D fanout494/X VGND VGND VPWR VPWR _6634_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_165_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3777_ input34/X _3295_/Y _3340_/Y input20/X VGND VGND VPWR VPWR _3777_/X sky130_fd_sc_hd__a22o_1
X_6565_ _7181_/CLK _6565_/D fanout499/X VGND VGND VPWR VPWR _6565_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_192_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5516_ hold85/X hold142/X _5519_/S VGND VGND VPWR VPWR _5516_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6496_ _6759_/CLK _6496_/D fanout488/X VGND VGND VPWR VPWR _6496_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_133_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5447_ _5579_/A0 hold389/X _5447_/S VGND VGND VPWR VPWR _5447_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5378_ _5459_/A0 hold337/X _5384_/S VGND VGND VPWR VPWR _5378_/X sky130_fd_sc_hd__mux2_1
X_4329_ hold453/X _6397_/A0 _4329_/S VGND VGND VPWR VPWR _4329_/X sky130_fd_sc_hd__mux2_1
X_7117_ _7133_/CLK _7117_/D fanout506/X VGND VGND VPWR VPWR _7117_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_113_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7048_ _7141_/CLK _7048_/D fanout504/X VGND VGND VPWR VPWR _7048_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_170_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3700_ _7035_/Q _5466_/A _4264_/A _6717_/Q _3699_/X VGND VGND VPWR VPWR _3701_/D
+ sky130_fd_sc_hd__a221o_1
X_4680_ _4784_/A _4692_/B VGND VGND VPWR VPWR _5083_/B sky130_fd_sc_hd__nor2_1
XFILLER_174_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3631_ _6884_/Q _5295_/A _5259_/A _6852_/Q _3608_/X VGND VGND VPWR VPWR _3632_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6350_ _6350_/A0 _3723_/X _6356_/S VGND VGND VPWR VPWR _7190_/D sky130_fd_sc_hd__mux2_1
X_3562_ _6901_/Q hold22/A _5376_/A _6957_/Q _3548_/X VGND VGND VPWR VPWR _3562_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_155_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5301_ _5550_/A0 hold532/X _5303_/S VGND VGND VPWR VPWR _5301_/X sky130_fd_sc_hd__mux2_1
X_6281_ _6718_/Q _6023_/B _6338_/B1 _6768_/Q _6271_/X VGND VGND VPWR VPWR _6281_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_142_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3493_ _6870_/Q _5277_/A _4016_/A _6515_/Q VGND VGND VPWR VPWR _3493_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5232_ _5232_/A _5571_/B VGND VGND VPWR VPWR _5240_/S sky130_fd_sc_hd__nand2_4
XFILLER_142_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5163_ _5163_/A _5163_/B _5163_/C VGND VGND VPWR VPWR _5163_/X sky130_fd_sc_hd__and3_1
XFILLER_96_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4114_ _5574_/A0 hold783/X hold97/X VGND VGND VPWR VPWR _4114_/X sky130_fd_sc_hd__mux2_1
X_5094_ _5094_/A _5094_/B VGND VGND VPWR VPWR _5095_/D sky130_fd_sc_hd__nor2_1
XFILLER_68_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4045_ _6397_/A0 hold671/X _4045_/S VGND VGND VPWR VPWR _4045_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5996_ _6014_/A _6030_/C VGND VGND VPWR VPWR _6019_/B sky130_fd_sc_hd__nand2_4
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4947_ _4947_/A _4947_/B VGND VGND VPWR VPWR _5064_/C sky130_fd_sc_hd__nor2_1
XFILLER_177_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4878_ _5124_/A _4987_/B VGND VGND VPWR VPWR _4878_/X sky130_fd_sc_hd__or2_1
X_6617_ _6617_/CLK _6617_/D _3873_/A VGND VGND VPWR VPWR _6617_/Q sky130_fd_sc_hd__dfrtp_4
X_3829_ _3252_/B _6541_/Q hold53/A VGND VGND VPWR VPWR _3831_/A sky130_fd_sc_hd__o21ai_1
XFILLER_118_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6548_ _7142_/CLK _6548_/D fanout525/X VGND VGND VPWR VPWR _6548_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6479_ _7002_/CLK _6479_/D fanout498/X VGND VGND VPWR VPWR _6479_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_106_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput260 _3950_/A VGND VGND VPWR VPWR pad_flash_io1_oeb sky130_fd_sc_hd__buf_12
Xoutput271 _6791_/Q VGND VGND VPWR VPWR pll_ena sky130_fd_sc_hd__buf_12
Xoutput282 _6474_/Q VGND VGND VPWR VPWR pll_trim[16] sky130_fd_sc_hd__buf_12
Xoutput293 _6492_/Q VGND VGND VPWR VPWR pll_trim[2] sky130_fd_sc_hd__buf_12
XFILLER_59_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire365 _6028_/Y VGND VGND VPWR VPWR _6094_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_156_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5850_ _6977_/Q _5960_/B VGND VGND VPWR VPWR _5850_/X sky130_fd_sc_hd__or2_1
X_4801_ _4674_/A _4595_/B _4569_/Y _4764_/A VGND VGND VPWR VPWR _4813_/B sky130_fd_sc_hd__a31o_1
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5781_ _7022_/Q _5663_/X _5683_/X _6870_/Q VGND VGND VPWR VPWR _5781_/X sky130_fd_sc_hd__a22o_1
XFILLER_9_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4732_ _4732_/A _4742_/A _4741_/C VGND VGND VPWR VPWR _5039_/A sky130_fd_sc_hd__and3_1
XFILLER_187_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4663_ _4664_/A _4814_/B VGND VGND VPWR VPWR _4663_/Y sky130_fd_sc_hd__nor2_1
XFILLER_174_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3614_ _6868_/Q _5277_/A hold31/A _6876_/Q VGND VGND VPWR VPWR _3614_/X sky130_fd_sc_hd__a22o_1
X_6402_ _6407_/A _6407_/B VGND VGND VPWR VPWR _6402_/X sky130_fd_sc_hd__and2_1
X_4594_ _5016_/A _5108_/A VGND VGND VPWR VPWR _4983_/A sky130_fd_sc_hd__nor2_1
Xhold902 hold902/A VGND VGND VPWR VPWR hold902/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold913 _5531_/X VGND VGND VPWR VPWR _7091_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3545_ _3544_/X _6787_/Q _3917_/A VGND VGND VPWR VPWR _6787_/D sky130_fd_sc_hd__mux2_1
X_6333_ _6715_/Q _6009_/X wire412/X _6669_/Q VGND VGND VPWR VPWR _6333_/X sky130_fd_sc_hd__a22o_1
Xhold924 _6923_/Q VGND VGND VPWR VPWR hold924/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold935 _4012_/X VGND VGND VPWR VPWR _6507_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_127_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold946 _6512_/Q VGND VGND VPWR VPWR hold946/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 _4065_/X VGND VGND VPWR VPWR _6551_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold968 hold968/A VGND VGND VPWR VPWR _6819_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6264_ _6602_/Q _5980_/Y _6036_/X _6517_/Q _6247_/X VGND VGND VPWR VPWR _6266_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3476_ _3476_/A _4111_/B VGND VGND VPWR VPWR _4010_/A sky130_fd_sc_hd__nor2_4
XFILLER_142_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold979 _6823_/Q VGND VGND VPWR VPWR hold979/X sky130_fd_sc_hd__dlygate4sd3_1
X_5215_ _5558_/A0 hold191/X _5220_/S VGND VGND VPWR VPWR _5215_/X sky130_fd_sc_hd__mux2_1
X_6195_ _6318_/S _6195_/A2 _6171_/S VGND VGND VPWR VPWR _6195_/X sky130_fd_sc_hd__o21a_1
Xhold1602 _7149_/Q VGND VGND VPWR VPWR _5617_/B1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5146_ _5172_/A _5172_/C _5170_/C VGND VGND VPWR VPWR _5147_/B sky130_fd_sc_hd__or3_1
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1613 _6542_/Q VGND VGND VPWR VPWR _3837_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5077_ _4659_/B _5021_/B _5027_/B _4582_/B _4860_/B VGND VGND VPWR VPWR _5077_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_151_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4028_ _4028_/A _4330_/B VGND VGND VPWR VPWR _4033_/S sky130_fd_sc_hd__and2_2
XFILLER_44_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5979_ _6040_/A _6030_/C VGND VGND VPWR VPWR _6038_/B sky130_fd_sc_hd__nand2_8
XFILLER_40_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold209 hold209/A VGND VGND VPWR VPWR hold209/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_125_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3330_ hold75/X _3330_/B VGND VGND VPWR VPWR hold76/A sky130_fd_sc_hd__nand2_8
XFILLER_124_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3261_ hold74/X hold66/X VGND VGND VPWR VPWR _3299_/A sky130_fd_sc_hd__and2b_4
XFILLER_124_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _4740_/Y _4999_/Y _4453_/A VGND VGND VPWR VPWR _5039_/B sky130_fd_sc_hd__a21oi_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3192_ _6543_/Q VGND VGND VPWR VPWR _3850_/B sky130_fd_sc_hd__inv_2
XFILLER_39_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6951_ _7079_/CLK _6951_/D fanout517/X VGND VGND VPWR VPWR _6951_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5902_ _6597_/Q _5691_/Y _5891_/X _5901_/X _6318_/S VGND VGND VPWR VPWR _5902_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_46_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6882_ _6882_/CLK _6882_/D _6407_/A VGND VGND VPWR VPWR _6882_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5833_ _6872_/Q _5683_/X _5685_/X _6912_/Q VGND VGND VPWR VPWR _5833_/X sky130_fd_sc_hd__a22o_1
XFILLER_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5764_ _6925_/Q _5955_/A2 _5700_/X _7029_/Q _5763_/X VGND VGND VPWR VPWR _5770_/A
+ sky130_fd_sc_hd__a221o_1
X_4715_ _4478_/Y _4563_/B _4670_/Y _4714_/X VGND VGND VPWR VPWR _4722_/B sky130_fd_sc_hd__a211o_1
X_5695_ _6898_/Q _5693_/X _5694_/X _7074_/Q _5692_/X VGND VGND VPWR VPWR _5708_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_135_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4646_ _4646_/A _4646_/B VGND VGND VPWR VPWR _4646_/X sky130_fd_sc_hd__or2_1
XFILLER_163_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold710 _5353_/X VGND VGND VPWR VPWR _6933_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold721 _6525_/Q VGND VGND VPWR VPWR hold721/X sky130_fd_sc_hd__dlygate4sd3_1
X_4577_ _4814_/B _5027_/A VGND VGND VPWR VPWR _5115_/A sky130_fd_sc_hd__nor2_1
XFILLER_162_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold732 _5264_/X VGND VGND VPWR VPWR _6854_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold743 _6524_/Q VGND VGND VPWR VPWR hold743/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold754 _4026_/X VGND VGND VPWR VPWR _6519_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6316_ _6341_/A _6316_/B _6316_/C VGND VGND VPWR VPWR _6316_/X sky130_fd_sc_hd__or3_1
XFILLER_116_674 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3528_ _3528_/A _3528_/B VGND VGND VPWR VPWR _4159_/A sky130_fd_sc_hd__nor2_2
XFILLER_143_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold765 _6966_/Q VGND VGND VPWR VPWR hold765/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold776 _5287_/X VGND VGND VPWR VPWR _6874_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 _6636_/Q VGND VGND VPWR VPWR hold787/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold798 _5441_/X VGND VGND VPWR VPWR _7011_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6247_ _7091_/Q _5642_/X _5992_/X hold87/A VGND VGND VPWR VPWR _6247_/X sky130_fd_sc_hd__a22o_1
X_3459_ _6950_/Q _5367_/A _5439_/A _7014_/Q VGND VGND VPWR VPWR _3459_/X sky130_fd_sc_hd__a22o_1
XFILLER_103_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6178_ _7101_/Q _6029_/B _6038_/Y _6984_/Q VGND VGND VPWR VPWR _6178_/X sky130_fd_sc_hd__a22o_1
Xhold1410 _6643_/Q VGND VGND VPWR VPWR hold1410/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1421 _6647_/Q VGND VGND VPWR VPWR _4190_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1432 _6781_/Q VGND VGND VPWR VPWR _5168_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5129_ _5123_/X _5128_/X _5160_/A VGND VGND VPWR VPWR _5139_/C sky130_fd_sc_hd__a21oi_2
Xhold1443 _7066_/Q VGND VGND VPWR VPWR hold1443/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1454 _5494_/X VGND VGND VPWR VPWR _7058_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1465 _3662_/X VGND VGND VPWR VPWR _6785_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1476 _6632_/Q VGND VGND VPWR VPWR _4172_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1487 _6694_/Q VGND VGND VPWR VPWR _3893_/B1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1498 _6652_/Q VGND VGND VPWR VPWR _4195_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold70 hold70/A VGND VGND VPWR VPWR hold70/X sky130_fd_sc_hd__buf_6
XFILLER_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold81 hold81/A VGND VGND VPWR VPWR hold81/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_63_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold92 hold92/A VGND VGND VPWR VPWR hold92/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4500_ _4351_/A _4351_/B _5076_/A _5021_/A _4391_/Y VGND VGND VPWR VPWR _4500_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_129_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5480_ _5549_/A0 hold639/X hold79/X VGND VGND VPWR VPWR _5480_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1 _5960_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4431_ _4846_/C _4459_/B VGND VGND VPWR VPWR _4871_/A sky130_fd_sc_hd__nand2_4
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7150_ _7183_/CLK _7150_/D fanout499/X VGND VGND VPWR VPWR _7150_/Q sky130_fd_sc_hd__dfrtp_1
X_4362_ _4428_/B _4426_/B VGND VGND VPWR VPWR _4957_/A sky130_fd_sc_hd__nor2_1
X_3313_ hold56/X _3313_/B VGND VGND VPWR VPWR _4120_/B sky130_fd_sc_hd__nand2_8
X_6101_ _6949_/Q _6024_/A _6205_/B1 _7061_/Q VGND VGND VPWR VPWR _6101_/X sky130_fd_sc_hd__a22o_1
Xfanout508 fanout527/X VGND VGND VPWR VPWR fanout508/X sky130_fd_sc_hd__buf_8
X_7081_ _7102_/CLK _7081_/D fanout502/X VGND VGND VPWR VPWR _7081_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_59_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4293_ _5549_/A0 hold631/X _4293_/S VGND VGND VPWR VPWR _4293_/X sky130_fd_sc_hd__mux2_1
Xfanout519 fanout521/X VGND VGND VPWR VPWR fanout519/X sky130_fd_sc_hd__buf_8
XFILLER_98_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3244_ _6468_/Q hold72/X VGND VGND VPWR VPWR _3244_/X sky130_fd_sc_hd__and2_1
X_6032_ _7111_/Q _6322_/B1 _6027_/D _6882_/Q _6031_/X VGND VGND VPWR VPWR _6044_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_591 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6934_ _7139_/CLK _6934_/D fanout518/X VGND VGND VPWR VPWR _6934_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6865_ _7088_/CLK _6865_/D fanout507/X VGND VGND VPWR VPWR _6865_/Q sky130_fd_sc_hd__dfrtp_2
X_5816_ _5816_/A0 _5815_/X _6171_/S VGND VGND VPWR VPWR _5816_/X sky130_fd_sc_hd__mux2_1
X_6796_ _7207_/CLK _6796_/D fanout484/X VGND VGND VPWR VPWR _6796_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_167_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5747_ _7044_/Q _5848_/B1 _5677_/X _6916_/Q _5746_/X VGND VGND VPWR VPWR _5750_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_157_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5678_ _7152_/Q _5705_/B _5706_/C VGND VGND VPWR VPWR _5678_/X sky130_fd_sc_hd__and3_4
XFILLER_163_522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4629_ _4814_/A _4784_/A VGND VGND VPWR VPWR _5017_/A sky130_fd_sc_hd__or2_1
Xhold540 _6734_/Q VGND VGND VPWR VPWR hold540/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold551 _4076_/X VGND VGND VPWR VPWR _6556_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold562 _7065_/Q VGND VGND VPWR VPWR hold562/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 _6895_/Q VGND VGND VPWR VPWR hold573/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold584 _4000_/X VGND VGND VPWR VPWR _6497_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 _6849_/Q VGND VGND VPWR VPWR hold595/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1240 _6686_/Q VGND VGND VPWR VPWR _4241_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1251 _4259_/X VGND VGND VPWR VPWR _6711_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1262 _5323_/X VGND VGND VPWR VPWR _6906_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1273 _6701_/Q VGND VGND VPWR VPWR _4247_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1284 _4325_/X VGND VGND VPWR VPWR _6766_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1295 _6516_/Q VGND VGND VPWR VPWR _4023_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput160 wb_dat_i[6] VGND VGND VPWR VPWR _6382_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_63_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4980_ _5059_/A _5130_/A _5158_/B VGND VGND VPWR VPWR _4980_/X sky130_fd_sc_hd__or3_1
X_3931_ _3930_/X input38/X _6461_/Q VGND VGND VPWR VPWR _3931_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6650_ _7187_/CLK _6650_/D VGND VGND VPWR VPWR _6650_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3862_ hold83/A _3862_/A1 _3866_/S VGND VGND VPWR VPWR _6450_/D sky130_fd_sc_hd__mux2_1
XFILLER_32_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5601_ _7144_/Q _7145_/Q _6565_/Q _5650_/A _5592_/Y VGND VGND VPWR VPWR _5601_/X
+ sky130_fd_sc_hd__o221a_1
X_6581_ _7142_/CLK _6581_/D fanout525/X VGND VGND VPWR VPWR _6581_/Q sky130_fd_sc_hd__dfrtp_1
X_3793_ hold72/A _6543_/Q VGND VGND VPWR VPWR _3794_/B sky130_fd_sc_hd__or2_1
XFILLER_145_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5532_ _5532_/A0 _6395_/A0 _5534_/S VGND VGND VPWR VPWR _5532_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_9_csclk _6820_/CLK VGND VGND VPWR VPWR _6725_/CLK sky130_fd_sc_hd__clkbuf_16
X_5463_ _5550_/A0 hold673/X _5465_/S VGND VGND VPWR VPWR _5463_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7202_ _3937_/A1 _7202_/D fanout529/X VGND VGND VPWR VPWR _7202_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_132_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4414_ _4819_/C _4538_/B _4935_/A VGND VGND VPWR VPWR _4435_/B sky130_fd_sc_hd__a21oi_1
X_5394_ _5394_/A _5571_/B VGND VGND VPWR VPWR _5402_/S sky130_fd_sc_hd__and2_4
X_7133_ _7133_/CLK _7133_/D fanout506/X VGND VGND VPWR VPWR _7133_/Q sky130_fd_sc_hd__dfrtp_1
X_4345_ _4846_/A _4570_/B _4846_/B _4570_/D VGND VGND VPWR VPWR _4781_/A sky130_fd_sc_hd__o211a_4
XFILLER_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4276_ _4276_/A _5580_/B VGND VGND VPWR VPWR _4281_/S sky130_fd_sc_hd__nand2_2
X_7064_ _7126_/CLK _7064_/D fanout524/X VGND VGND VPWR VPWR _7064_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6015_ _6039_/C _6020_/C _6040_/C VGND VGND VPWR VPWR _6015_/X sky130_fd_sc_hd__and3_4
X_3227_ _6901_/Q VGND VGND VPWR VPWR _3227_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6917_ _7140_/CLK _6917_/D fanout522/X VGND VGND VPWR VPWR _6917_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_52_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6848_ _7110_/CLK _6848_/D fanout506/X VGND VGND VPWR VPWR _6848_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6779_ _3937_/A1 _6779_/D fanout529/X VGND VGND VPWR VPWR _6779_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_183_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold370 _4015_/X VGND VGND VPWR VPWR _6510_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 _6550_/Q VGND VGND VPWR VPWR hold381/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold392 _5207_/X VGND VGND VPWR VPWR _6808_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1070 _5545_/X VGND VGND VPWR VPWR _7103_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1081 _6828_/Q VGND VGND VPWR VPWR _5235_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1092 _6661_/Q VGND VGND VPWR VPWR _4206_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_210 _6981_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_221 _4085_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_232 _5539_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_243 _5466_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_254 input38/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__1134_ clkbuf_0__1134_/X VGND VGND VPWR VPWR _6353_/A1 sky130_fd_sc_hd__clkbuf_16
XFILLER_114_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4130_ _4130_/A0 _6393_/A0 _4134_/S VGND VGND VPWR VPWR _4130_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4061_ hold952/X _4060_/X _4069_/S VGND VGND VPWR VPWR _4061_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4963_ _4963_/A _4963_/B VGND VGND VPWR VPWR _5112_/B sky130_fd_sc_hd__or2_1
XFILLER_51_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6702_ _6707_/CLK _6702_/D _6432_/A VGND VGND VPWR VPWR _6702_/Q sky130_fd_sc_hd__dfrtp_1
X_3914_ _3914_/A1 _3914_/A2 _3835_/S _3834_/B _3252_/B VGND VGND VPWR VPWR _6544_/D
+ sky130_fd_sc_hd__o32ai_1
X_4894_ _4965_/B _4894_/B _4894_/C _4490_/X VGND VGND VPWR VPWR _4896_/C sky130_fd_sc_hd__or4b_1
XFILLER_149_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6633_ _7196_/CLK _6633_/D VGND VGND VPWR VPWR _6633_/Q sky130_fd_sc_hd__dfxtp_1
X_3845_ input58/X _3845_/A1 _3845_/S VGND VGND VPWR VPWR _6457_/D sky130_fd_sc_hd__mux2_1
XFILLER_20_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6564_ _7182_/CLK _6564_/D fanout499/X VGND VGND VPWR VPWR _6564_/Q sky130_fd_sc_hd__dfrtp_4
X_3776_ _7143_/Q _5221_/B _6392_/A _7207_/Q _3775_/X VGND VGND VPWR VPWR _3781_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_138_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5515_ _5539_/A1 _5515_/A1 _5519_/S VGND VGND VPWR VPWR _5515_/X sky130_fd_sc_hd__mux2_1
X_6495_ _6759_/CLK _6495_/D fanout488/X VGND VGND VPWR VPWR _6495_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_173_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5446_ _5587_/A0 hold821/X _5447_/S VGND VGND VPWR VPWR _5446_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5377_ _5521_/A0 _5377_/A1 _5384_/S VGND VGND VPWR VPWR _5377_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7116_ _7134_/CLK _7116_/D fanout525/X VGND VGND VPWR VPWR _7116_/Q sky130_fd_sc_hd__dfrtp_1
X_4328_ hold235/X _5539_/A1 _4329_/S VGND VGND VPWR VPWR _4328_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7047_ _7079_/CLK _7047_/D fanout516/X VGND VGND VPWR VPWR _7047_/Q sky130_fd_sc_hd__dfrtp_4
X_4259_ _4259_/A0 _5521_/A0 _4263_/S VGND VGND VPWR VPWR _4259_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_534 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3630_ _6636_/Q _4174_/A _4258_/A _6713_/Q _3610_/X VGND VGND VPWR VPWR _3632_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_186_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3561_ _7053_/Q _3684_/B1 _4028_/A _6524_/Q VGND VGND VPWR VPWR _3561_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5300_ _5567_/A0 hold647/X _5303_/S VGND VGND VPWR VPWR _5300_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3492_ _3536_/A _3729_/B VGND VGND VPWR VPWR _4016_/A sky130_fd_sc_hd__nor2_4
X_6280_ _6280_/A _6280_/B _6280_/C _6280_/D VGND VGND VPWR VPWR _6280_/X sky130_fd_sc_hd__or4_1
XFILLER_142_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5231_ _6394_/A0 _5231_/A1 _5231_/S VGND VGND VPWR VPWR _5231_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5162_ _5162_/A _5162_/B _5162_/C _5162_/D VGND VGND VPWR VPWR _5163_/C sky130_fd_sc_hd__nor4_1
Xclkbuf_leaf_12_csclk _6882_/CLK VGND VGND VPWR VPWR _6617_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_111_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4113_ _5459_/A0 hold237/X hold97/X VGND VGND VPWR VPWR _4113_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5093_ _4485_/A _4870_/B _5083_/A _4785_/X VGND VGND VPWR VPWR _5114_/C sky130_fd_sc_hd__a211o_1
XFILLER_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4044_ _6396_/A0 hold747/X _4045_/S VGND VGND VPWR VPWR _4044_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_27_csclk _6882_/CLK VGND VGND VPWR VPWR _7130_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_52_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5995_ _6498_/Q _5642_/X _5994_/X _7074_/Q VGND VGND VPWR VPWR _5995_/X sky130_fd_sc_hd__a22o_1
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4946_ _5064_/B _5126_/C _5053_/B _4945_/X VGND VGND VPWR VPWR _4960_/A sky130_fd_sc_hd__or4b_1
XFILLER_193_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4877_ _4657_/C _4524_/B _4983_/B VGND VGND VPWR VPWR _5049_/C sky130_fd_sc_hd__a21o_1
X_6616_ _6617_/CLK _6616_/D _3873_/A VGND VGND VPWR VPWR _6616_/Q sky130_fd_sc_hd__dfrtp_4
X_3828_ _3827_/X _3828_/A1 _3833_/S VGND VGND VPWR VPWR _6465_/D sky130_fd_sc_hd__mux2_1
XFILLER_20_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6547_ _7142_/CLK _6547_/D fanout525/X VGND VGND VPWR VPWR _6547_/Q sky130_fd_sc_hd__dfrtp_1
X_3759_ _7119_/Q _5562_/A hold31/A _6874_/Q _3737_/X VGND VGND VPWR VPWR _3760_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_192_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6478_ _6825_/CLK _6478_/D fanout490/X VGND VGND VPWR VPWR _6478_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_133_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5429_ _5552_/A0 hold723/X _5429_/S VGND VGND VPWR VPWR _5429_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput250 _3927_/X VGND VGND VPWR VPWR mgmt_gpio_out[9] sky130_fd_sc_hd__clkbuf_1
Xoutput261 _6801_/Q VGND VGND VPWR VPWR pll90_sel[0] sky130_fd_sc_hd__buf_12
XFILLER_121_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput272 _6798_/Q VGND VGND VPWR VPWR pll_sel[0] sky130_fd_sc_hd__buf_12
Xoutput283 _6475_/Q VGND VGND VPWR VPWR pll_trim[17] sky130_fd_sc_hd__buf_12
XFILLER_59_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput294 _6493_/Q VGND VGND VPWR VPWR pll_trim[3] sky130_fd_sc_hd__buf_12
XFILLER_114_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_1_1_1_wb_clk_i clkbuf_1_1_1_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_2_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_8
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4800_ _4569_/Y _4684_/B _4753_/Y VGND VGND VPWR VPWR _5090_/A sky130_fd_sc_hd__a21o_1
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5780_ _6958_/Q _5659_/X _5705_/X _6942_/Q _5779_/X VGND VGND VPWR VPWR _5785_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4731_ _4484_/B _4731_/B _4731_/C VGND VGND VPWR VPWR _4741_/C sky130_fd_sc_hd__and3b_1
XFILLER_187_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4662_ _4931_/A _4674_/A VGND VGND VPWR VPWR _4683_/B sky130_fd_sc_hd__nand2_2
X_6401_ _6407_/A _6407_/B VGND VGND VPWR VPWR _6401_/X sky130_fd_sc_hd__and2_1
X_3613_ _6948_/Q _5367_/A _5385_/A _6964_/Q VGND VGND VPWR VPWR _3613_/X sky130_fd_sc_hd__a22o_1
X_4593_ _4814_/A _4707_/A VGND VGND VPWR VPWR _5108_/A sky130_fd_sc_hd__or2_4
Xhold903 _5542_/X VGND VGND VPWR VPWR _7101_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_134_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6332_ _6332_/A _6332_/B _6332_/C VGND VGND VPWR VPWR _6332_/X sky130_fd_sc_hd__or3_1
Xhold914 _6916_/Q VGND VGND VPWR VPWR hold914/X sky130_fd_sc_hd__dlygate4sd3_1
X_3544_ _6353_/A1 _3603_/A1 _3791_/A VGND VGND VPWR VPWR _3544_/X sky130_fd_sc_hd__mux2_1
Xhold925 _5342_/X VGND VGND VPWR VPWR _6923_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold936 _7024_/Q VGND VGND VPWR VPWR hold936/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold947 _4018_/X VGND VGND VPWR VPWR _6512_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold958 _6532_/Q VGND VGND VPWR VPWR hold958/X sky130_fd_sc_hd__dlygate4sd3_1
X_6263_ _6607_/Q _6326_/A2 _6021_/Y _6622_/Q _6262_/X VGND VGND VPWR VPWR _6266_/B
+ sky130_fd_sc_hd__a221o_1
Xhold969 _7207_/Q VGND VGND VPWR VPWR hold969/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3475_ input16/X _3268_/Y _4264_/A _6720_/Q _3473_/X VGND VGND VPWR VPWR _3484_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_103_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5214_ _5221_/B _5535_/B VGND VGND VPWR VPWR _5220_/S sky130_fd_sc_hd__nand2_2
X_6194_ _6848_/Q _6094_/A _6193_/X _5650_/A VGND VGND VPWR VPWR _6194_/X sky130_fd_sc_hd__a211o_1
XFILLER_130_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1603 _7141_/Q VGND VGND VPWR VPWR hold906/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5145_ _5145_/A _5145_/B _5144_/X VGND VGND VPWR VPWR _5170_/C sky130_fd_sc_hd__or3b_1
Xhold1614 _7185_/Q VGND VGND VPWR VPWR _6318_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5076_ _5076_/A _5076_/B VGND VGND VPWR VPWR _5108_/B sky130_fd_sc_hd__and2_2
XFILLER_44_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4027_ hold715/X _5534_/A1 _4027_/S VGND VGND VPWR VPWR _4027_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5978_ _7156_/Q _7155_/Q VGND VGND VPWR VPWR _6030_/C sky130_fd_sc_hd__nor2_4
X_4929_ _4929_/A1 _4232_/X _4825_/X _4928_/X VGND VGND VPWR VPWR _6777_/D sky130_fd_sc_hd__o22a_1
XFILLER_166_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ hold65/X _5034_/B2 _3971_/S VGND VGND VPWR VPWR hold66/A sky130_fd_sc_hd__mux2_2
XFILLER_140_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3191_ _3191_/A VGND VGND VPWR VPWR _3191_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6950_ _7078_/CLK _6950_/D fanout514/X VGND VGND VPWR VPWR _6950_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_53_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5901_ _5901_/A _5901_/B _5901_/C _5901_/D VGND VGND VPWR VPWR _5901_/X sky130_fd_sc_hd__or4_1
XFILLER_34_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6881_ _7126_/CLK _6881_/D fanout523/X VGND VGND VPWR VPWR _6881_/Q sky130_fd_sc_hd__dfrtp_4
X_5832_ _6952_/Q _5666_/X _5705_/X _6944_/Q _5831_/X VGND VGND VPWR VPWR _5835_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_34_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5763_ _7037_/Q _5696_/X _5697_/X _6989_/Q VGND VGND VPWR VPWR _5763_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4714_ _4714_/A _4714_/B _4822_/A _4882_/B VGND VGND VPWR VPWR _4714_/X sky130_fd_sc_hd__or4b_1
X_5694_ _7152_/Q _5706_/C _5703_/C VGND VGND VPWR VPWR _5694_/X sky130_fd_sc_hd__and3_4
XFILLER_187_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4645_ _5076_/B _4653_/C VGND VGND VPWR VPWR _4645_/X sky130_fd_sc_hd__or2_1
XFILLER_30_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold700 _4108_/X VGND VGND VPWR VPWR _6577_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold711 _6764_/Q VGND VGND VPWR VPWR hold711/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_146_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4576_ _4814_/A _4814_/C VGND VGND VPWR VPWR _5027_/A sky130_fd_sc_hd__or2_4
Xhold722 _4033_/X VGND VGND VPWR VPWR _6525_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap430 _5203_/B VGND VGND VPWR VPWR hold113/A sky130_fd_sc_hd__buf_12
Xhold733 _7041_/Q VGND VGND VPWR VPWR hold733/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold744 _4032_/X VGND VGND VPWR VPWR _6524_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6315_ _6315_/A _6315_/B _6315_/C _6315_/D VGND VGND VPWR VPWR _6316_/C sky130_fd_sc_hd__or4_1
Xhold755 hold755/A VGND VGND VPWR VPWR hold755/X sky130_fd_sc_hd__dlygate4sd3_1
X_3527_ _6540_/Q _4046_/A _5187_/A _6797_/Q VGND VGND VPWR VPWR _3527_/X sky130_fd_sc_hd__a22o_1
XFILLER_190_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold766 _5390_/X VGND VGND VPWR VPWR _6966_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 _6705_/Q VGND VGND VPWR VPWR hold777/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 _4177_/X VGND VGND VPWR VPWR _6636_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6246_ _6727_/Q _6320_/A2 _6320_/B1 _6617_/Q VGND VGND VPWR VPWR _6246_/X sky130_fd_sc_hd__a22o_2
Xhold799 hold799/A VGND VGND VPWR VPWR hold799/X sky130_fd_sc_hd__dlygate4sd3_1
X_3458_ _6690_/Q _4240_/A _4040_/A _6535_/Q _3457_/X VGND VGND VPWR VPWR _3468_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_76_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6177_ _7008_/Q _6202_/B1 _6176_/X VGND VGND VPWR VPWR _6180_/C sky130_fd_sc_hd__a21o_1
XFILLER_162_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3389_ _6928_/Q _5340_/A _5358_/A _6944_/Q VGND VGND VPWR VPWR _3389_/X sky130_fd_sc_hd__a22o_1
Xhold1400 _6645_/Q VGND VGND VPWR VPWR hold1400/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1411 _6654_/Q VGND VGND VPWR VPWR hold1411/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1422 _7194_/Q VGND VGND VPWR VPWR _6354_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1433 _3300_/A VGND VGND VPWR VPWR _3462_/B sky130_fd_sc_hd__dlygate4sd3_1
X_5128_ _5160_/B _5128_/B _5128_/C _5159_/B VGND VGND VPWR VPWR _5128_/X sky130_fd_sc_hd__and4b_1
XFILLER_111_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1444 _5503_/X VGND VGND VPWR VPWR _7066_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1455 _7201_/Q VGND VGND VPWR VPWR _6377_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_55_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1466 _6784_/Q VGND VGND VPWR VPWR _3725_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1477 _6584_/Q VGND VGND VPWR VPWR hold179/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5059_ _5059_/A _5059_/B _5059_/C VGND VGND VPWR VPWR _5159_/A sky130_fd_sc_hd__nor3_1
Xhold1488 hold38/A VGND VGND VPWR VPWR _3860_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1499 _6693_/Q VGND VGND VPWR VPWR _3892_/B1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold60 hold60/A VGND VGND VPWR VPWR hold60/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 hold71/A VGND VGND VPWR VPWR hold71/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_36_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold82 hold82/A VGND VGND VPWR VPWR hold82/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 hold93/A VGND VGND VPWR VPWR hold93/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_662 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4430_ _4570_/D _4738_/A VGND VGND VPWR VPWR _4931_/B sky130_fd_sc_hd__nor2_4
XFILLER_6_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_2 _3278_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4361_ _4341_/X _4781_/A _4360_/B _4605_/A VGND VGND VPWR VPWR _4426_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_98_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6100_ _7130_/Q _6320_/A2 _6320_/B1 _6877_/Q _6099_/X VGND VGND VPWR VPWR _6110_/A
+ sky130_fd_sc_hd__a221o_1
X_3312_ _3526_/A _3528_/A VGND VGND VPWR VPWR _5268_/A sky130_fd_sc_hd__nor2_8
XFILLER_98_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7080_ _7080_/CLK _7080_/D fanout502/X VGND VGND VPWR VPWR _7080_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_112_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout509 fanout510/X VGND VGND VPWR VPWR fanout509/X sky130_fd_sc_hd__buf_8
X_4292_ hold36/X hold150/X _4293_/S VGND VGND VPWR VPWR _4292_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6031_ _6906_/Q _6024_/C _6030_/X _6994_/Q VGND VGND VPWR VPWR _6031_/X sky130_fd_sc_hd__a22o_1
X_3243_ hold46/X hold72/X hold92/X VGND VGND VPWR VPWR hold93/A sky130_fd_sc_hd__a21oi_1
XFILLER_98_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6933_ _7049_/CLK _6933_/D fanout522/X VGND VGND VPWR VPWR _6933_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6864_ _7088_/CLK _6864_/D fanout506/X VGND VGND VPWR VPWR _6864_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_179_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5815_ _5650_/A _7166_/Q _5814_/X VGND VGND VPWR VPWR _5815_/X sky130_fd_sc_hd__a21o_1
XFILLER_179_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6795_ _7207_/CLK _6795_/D fanout484/X VGND VGND VPWR VPWR _6795_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_148_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5746_ _6876_/Q _5667_/X _5703_/X _6852_/Q VGND VGND VPWR VPWR _5746_/X sky130_fd_sc_hd__a22o_1
XFILLER_182_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5677_ _5938_/B _5703_/C _5699_/C VGND VGND VPWR VPWR _5677_/X sky130_fd_sc_hd__and3_4
XFILLER_108_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4628_ _4675_/A _4646_/B VGND VGND VPWR VPWR _5083_/A sky130_fd_sc_hd__nor2_2
Xhold530 _6775_/Q VGND VGND VPWR VPWR hold530/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold541 _4286_/X VGND VGND VPWR VPWR _6734_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4559_ _4560_/A _4573_/B VGND VGND VPWR VPWR _4797_/A sky130_fd_sc_hd__and2_2
Xhold552 _6802_/Q VGND VGND VPWR VPWR hold552/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold563 _5501_/X VGND VGND VPWR VPWR _7065_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 _5310_/X VGND VGND VPWR VPWR _6895_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold585 _6610_/Q VGND VGND VPWR VPWR hold585/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 _5258_/X VGND VGND VPWR VPWR _6849_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6229_ _6771_/Q _6002_/Y _6007_/Y _6756_/Q _6228_/X VGND VGND VPWR VPWR _6232_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_77_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1230 _6850_/Q VGND VGND VPWR VPWR _5260_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1241 _4241_/X VGND VGND VPWR VPWR _6686_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1252 _6531_/Q VGND VGND VPWR VPWR _4041_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1263 _6596_/Q VGND VGND VPWR VPWR _4130_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1274 _4247_/X VGND VGND VPWR VPWR _6701_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1285 hold1611/X VGND VGND VPWR VPWR _4265_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1296 _4023_/X VGND VGND VPWR VPWR _6516_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput150 wb_dat_i[26] VGND VGND VPWR VPWR _6370_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput161 wb_dat_i[7] VGND VGND VPWR VPWR _6385_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3930_ _6555_/Q _6790_/Q _6440_/B VGND VGND VPWR VPWR _3930_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3861_ _3862_/A1 hold1/A _3866_/S VGND VGND VPWR VPWR _3861_/X sky130_fd_sc_hd__mux2_1
XFILLER_189_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5600_ _7144_/Q _7145_/Q VGND VGND VPWR VPWR _5600_/Y sky130_fd_sc_hd__nand2_1
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6580_ _7142_/CLK _6580_/D fanout525/X VGND VGND VPWR VPWR _6580_/Q sky130_fd_sc_hd__dfrtp_1
X_3792_ _3792_/A1 _3917_/A _3790_/X _3791_/Y VGND VGND VPWR VPWR _6783_/D sky130_fd_sc_hd__a22o_1
XFILLER_192_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5531_ hold912/X _5531_/A1 _5534_/S VGND VGND VPWR VPWR _5531_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5462_ _5549_/A0 hold623/X _5465_/S VGND VGND VPWR VPWR _5462_/X sky130_fd_sc_hd__mux2_1
X_7201_ _3937_/A1 _7201_/D fanout529/X VGND VGND VPWR VPWR _7201_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4413_ _4819_/C _4538_/B _4435_/A VGND VGND VPWR VPWR _4434_/B sky130_fd_sc_hd__a21boi_2
X_5393_ _5552_/A0 hold601/X _5393_/S VGND VGND VPWR VPWR _5393_/X sky130_fd_sc_hd__mux2_1
X_7132_ _7132_/CLK _7132_/D fanout525/X VGND VGND VPWR VPWR _7132_/Q sky130_fd_sc_hd__dfrtp_1
X_4344_ _4846_/A _4570_/B VGND VGND VPWR VPWR _4596_/B sky130_fd_sc_hd__or2_1
XFILLER_86_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7063_ _7108_/CLK _7063_/D fanout523/X VGND VGND VPWR VPWR _7063_/Q sky130_fd_sc_hd__dfrtp_2
X_4275_ hold571/X _5549_/A0 _4275_/S VGND VGND VPWR VPWR _4275_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6014_ _6014_/A _6039_/A _6020_/C VGND VGND VPWR VPWR _6022_/C sky130_fd_sc_hd__and3_1
XFILLER_140_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3226_ _6909_/Q VGND VGND VPWR VPWR _3226_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_278 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6916_ _7128_/CLK _6916_/D fanout514/X VGND VGND VPWR VPWR _6916_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_70_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6847_ _7065_/CLK _6847_/D fanout517/X VGND VGND VPWR VPWR _6847_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6778_ _3937_/A1 _6778_/D fanout529/X VGND VGND VPWR VPWR _6778_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_139_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5729_ _6843_/Q _5691_/Y _5719_/X _5728_/X _3195_/Y VGND VGND VPWR VPWR _5729_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_182_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold360 _5468_/X VGND VGND VPWR VPWR _7035_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold371 _7096_/Q VGND VGND VPWR VPWR hold371/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 _4063_/X VGND VGND VPWR VPWR _6550_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 _7126_/Q VGND VGND VPWR VPWR hold393/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1060 _5186_/X VGND VGND VPWR VPWR _6792_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1071 _7127_/Q VGND VGND VPWR VPWR _5572_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1082 _5235_/X VGND VGND VPWR VPWR _6828_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1093 _4206_/X VGND VGND VPWR VPWR _6661_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_200 _5411_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_211 _6762_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_222 _5571_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_233 _5583_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_244 _4028_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_255 _5583_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4060_ hold472/X _5557_/A0 _4068_/S VGND VGND VPWR VPWR _4060_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4962_ _5068_/B _4962_/B VGND VGND VPWR VPWR _4962_/Y sky130_fd_sc_hd__nor2_1
X_3913_ _3913_/A1 _6541_/Q _3834_/B _3913_/B1 VGND VGND VPWR VPWR _6545_/D sky130_fd_sc_hd__a31o_1
X_6701_ _6707_/CLK _6701_/D _6432_/A VGND VGND VPWR VPWR _6701_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_51_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4893_ _4524_/B _4871_/Y _4892_/X VGND VGND VPWR VPWR _4894_/B sky130_fd_sc_hd__a21o_1
X_6632_ _7196_/CLK _6632_/D VGND VGND VPWR VPWR _6632_/Q sky130_fd_sc_hd__dfxtp_1
X_3844_ _6473_/Q _6472_/Q _6471_/Q _6541_/Q VGND VGND VPWR VPWR _3845_/S sky130_fd_sc_hd__or4b_1
XFILLER_20_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6563_ _7181_/CLK _6563_/D fanout502/X VGND VGND VPWR VPWR _6563_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_158_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3775_ _6798_/Q _5193_/A _5529_/A _7090_/Q VGND VGND VPWR VPWR _3775_/X sky130_fd_sc_hd__a22o_1
XFILLER_164_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5514_ _5583_/A0 hold307/X _5519_/S VGND VGND VPWR VPWR _5514_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6494_ _6759_/CLK _6494_/D fanout488/X VGND VGND VPWR VPWR _6494_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_145_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5445_ _5586_/A0 hold985/X _5447_/S VGND VGND VPWR VPWR _5445_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5376_ _5376_/A _5580_/B VGND VGND VPWR VPWR _5384_/S sky130_fd_sc_hd__nand2_8
XFILLER_154_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7115_ _7115_/CLK _7115_/D fanout508/X VGND VGND VPWR VPWR _7115_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4327_ hold683/X _4327_/A1 _4329_/S VGND VGND VPWR VPWR _4327_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7046_ _7070_/CLK _7046_/D fanout510/X VGND VGND VPWR VPWR _7046_/Q sky130_fd_sc_hd__dfrtp_4
X_4258_ _4258_/A _5580_/B VGND VGND VPWR VPWR _4263_/S sky130_fd_sc_hd__and2_1
XFILLER_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3209_ _7045_/Q VGND VGND VPWR VPWR _3209_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4189_ _6694_/Q _6348_/B VGND VGND VPWR VPWR _4197_/S sky130_fd_sc_hd__and2_4
XFILLER_28_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold190 _5291_/X VGND VGND VPWR VPWR _6878_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_8_csclk _6820_/CLK VGND VGND VPWR VPWR _6963_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_160_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3560_ _6989_/Q _3298_/Y _3471_/Y _6764_/Q VGND VGND VPWR VPWR _3560_/X sky130_fd_sc_hd__a22o_1
XFILLER_10_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3491_ _6715_/Q _4258_/A _4300_/A _6750_/Q _3488_/X VGND VGND VPWR VPWR _3499_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_5_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5230_ _5212_/C _5230_/A1 _5231_/S VGND VGND VPWR VPWR _5230_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5161_ _4638_/B _4704_/B _4490_/X VGND VGND VPWR VPWR _5162_/D sky130_fd_sc_hd__o21ai_1
XFILLER_68_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4112_ _5581_/A0 hold793/X hold97/X VGND VGND VPWR VPWR _4112_/X sky130_fd_sc_hd__mux2_1
X_5092_ _5119_/A _5119_/B _5170_/B _5092_/D VGND VGND VPWR VPWR _5102_/A sky130_fd_sc_hd__or4_1
XFILLER_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4043_ _6395_/A0 _4043_/A1 _4045_/S VGND VGND VPWR VPWR _4043_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5994_ _6040_/A _6039_/A _6040_/B VGND VGND VPWR VPWR _5994_/X sky130_fd_sc_hd__and3_4
X_4945_ _4846_/A _4483_/A _4944_/X _4839_/A _4847_/A VGND VGND VPWR VPWR _4945_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_177_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4876_ _4876_/A _4971_/B VGND VGND VPWR VPWR _4887_/D sky130_fd_sc_hd__nand2_1
XFILLER_177_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6615_ _6708_/CLK _6615_/D fanout494/X VGND VGND VPWR VPWR _6615_/Q sky130_fd_sc_hd__dfrtp_2
X_3827_ hold53/A hold72/A _3820_/Y _3826_/X VGND VGND VPWR VPWR _3827_/X sky130_fd_sc_hd__a22o_1
XFILLER_137_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6546_ _7140_/CLK _6546_/D fanout525/X VGND VGND VPWR VPWR _6546_/Q sky130_fd_sc_hd__dfrtp_1
X_3758_ _6906_/Q _5322_/A _4300_/A _6746_/Q _3728_/X VGND VGND VPWR VPWR _3760_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_180_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6477_ _6825_/CLK _6477_/D fanout490/X VGND VGND VPWR VPWR _6477_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_118_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3689_ _3689_/A _3689_/B VGND VGND VPWR VPWR _3723_/B sky130_fd_sc_hd__or2_1
XFILLER_133_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5428_ _5587_/A0 hold892/X _5429_/S VGND VGND VPWR VPWR _5428_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput240 _6576_/Q VGND VGND VPWR VPWR mgmt_gpio_out[34] sky130_fd_sc_hd__buf_12
Xoutput251 _3945_/X VGND VGND VPWR VPWR pad_flash_clk sky130_fd_sc_hd__clkbuf_1
Xoutput262 _6802_/Q VGND VGND VPWR VPWR pll90_sel[1] sky130_fd_sc_hd__buf_12
Xoutput273 _6799_/Q VGND VGND VPWR VPWR pll_sel[1] sky130_fd_sc_hd__buf_12
XFILLER_121_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput284 _6476_/Q VGND VGND VPWR VPWR pll_trim[18] sky130_fd_sc_hd__buf_12
X_5359_ _5521_/A0 _5359_/A1 _5366_/S VGND VGND VPWR VPWR _5359_/X sky130_fd_sc_hd__mux2_1
Xoutput295 _6494_/Q VGND VGND VPWR VPWR pll_trim[4] sky130_fd_sc_hd__buf_12
XFILLER_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7029_ _7037_/CLK _7029_/D fanout515/X VGND VGND VPWR VPWR _7029_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_74_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4730_ _4981_/B _5002_/A VGND VGND VPWR VPWR _4815_/A sky130_fd_sc_hd__nor2_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4661_ _5023_/A _4693_/A VGND VGND VPWR VPWR _4704_/B sky130_fd_sc_hd__or2_2
XFILLER_187_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6400_ _6433_/A _6441_/B VGND VGND VPWR VPWR _6400_/X sky130_fd_sc_hd__and2_1
X_3612_ _6940_/Q _5358_/A _4264_/A _6718_/Q VGND VGND VPWR VPWR _3612_/X sky130_fd_sc_hd__a22o_1
X_4592_ _4707_/A VGND VGND VPWR VPWR _4592_/Y sky130_fd_sc_hd__inv_2
XFILLER_190_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6331_ _6331_/A _6331_/B _6331_/C _6331_/D VGND VGND VPWR VPWR _6332_/C sky130_fd_sc_hd__or4_1
Xhold904 _6939_/Q VGND VGND VPWR VPWR hold904/X sky130_fd_sc_hd__dlygate4sd3_1
X_3543_ _3543_/A _3543_/B _3543_/C VGND VGND VPWR VPWR _3543_/X sky130_fd_sc_hd__or3_2
XFILLER_127_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold915 _5334_/X VGND VGND VPWR VPWR _6916_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold926 _7080_/Q VGND VGND VPWR VPWR hold926/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold937 _5455_/X VGND VGND VPWR VPWR _7024_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold948 _6752_/Q VGND VGND VPWR VPWR hold948/X sky130_fd_sc_hd__dlygate4sd3_1
X_6262_ _6687_/Q _5982_/X _6040_/X _6527_/Q VGND VGND VPWR VPWR _6262_/X sky130_fd_sc_hd__a22o_1
Xhold959 _4042_/X VGND VGND VPWR VPWR _6532_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3474_ _3546_/A _3528_/B VGND VGND VPWR VPWR _4264_/A sky130_fd_sc_hd__nor2_4
XFILLER_115_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5213_ hold962/X _3727_/Y _4330_/B _5212_/X VGND VGND VPWR VPWR _5213_/X sky130_fd_sc_hd__o211a_1
XFILLER_103_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6193_ _6193_/A _6193_/B _6193_/C VGND VGND VPWR VPWR _6193_/X sky130_fd_sc_hd__or3_1
XFILLER_142_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5144_ _4794_/A _5143_/Y _4810_/C _4631_/B VGND VGND VPWR VPWR _5144_/X sky130_fd_sc_hd__o211a_1
Xhold1604 hold25/A VGND VGND VPWR VPWR _3833_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5075_ _5018_/A _5074_/X _5029_/B _5013_/X _4911_/X VGND VGND VPWR VPWR _5156_/B
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_151_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4026_ hold753/X _5533_/A1 _4027_/S VGND VGND VPWR VPWR _4026_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5977_ _6014_/A _6039_/A _6040_/B VGND VGND VPWR VPWR _5977_/X sky130_fd_sc_hd__and3_4
X_4928_ _6362_/A _4928_/B _4928_/C _4928_/D VGND VGND VPWR VPWR _4928_/X sky130_fd_sc_hd__or4_1
XFILLER_21_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4859_ _5023_/B _4582_/B _4858_/X _4504_/A VGND VGND VPWR VPWR _4860_/D sky130_fd_sc_hd__o211a_1
XFILLER_166_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6529_ _7207_/CLK _6529_/D fanout484/X VGND VGND VPWR VPWR _6529_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_180_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_73_csclk _6753_/CLK VGND VGND VPWR VPWR _6759_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_11_csclk clkbuf_opt_2_0_csclk/X VGND VGND VPWR VPWR _6683_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_7_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_26_csclk _6882_/CLK VGND VGND VPWR VPWR _7135_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_124_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3190_ hold72/X VGND VGND VPWR VPWR _3252_/B sky130_fd_sc_hd__clkinv_2
XFILLER_94_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5900_ _6702_/Q _5659_/X _5700_/X _6507_/Q _5899_/X VGND VGND VPWR VPWR _5901_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_93_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6880_ _7126_/CLK _6880_/D fanout524/X VGND VGND VPWR VPWR _6880_/Q sky130_fd_sc_hd__dfrtp_4
X_5831_ _6888_/Q _5846_/A2 _5848_/B1 _7048_/Q VGND VGND VPWR VPWR _5831_/X sky130_fd_sc_hd__a22o_1
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5762_ _6933_/Q _5670_/X _5686_/X _7013_/Q _5761_/X VGND VGND VPWR VPWR _5771_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4713_ _4713_/A _4713_/B _4713_/C _4713_/D VGND VGND VPWR VPWR _4714_/B sky130_fd_sc_hd__nand4_1
X_5693_ _5938_/B _5706_/B _5700_/C VGND VGND VPWR VPWR _5693_/X sky130_fd_sc_hd__and3_4
XFILLER_147_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4644_ _5059_/A _4644_/B _5095_/A _4643_/X VGND VGND VPWR VPWR _4647_/B sky130_fd_sc_hd__or4b_1
Xhold701 _7054_/Q VGND VGND VPWR VPWR hold701/X sky130_fd_sc_hd__dlygate4sd3_1
X_4575_ _4605_/A _4610_/A _4621_/C VGND VGND VPWR VPWR _4814_/C sky130_fd_sc_hd__or3_4
Xhold712 _4322_/X VGND VGND VPWR VPWR _6764_/D sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap420 _5676_/X VGND VGND VPWR VPWR _5848_/B1 sky130_fd_sc_hd__buf_12
Xhold723 _7001_/Q VGND VGND VPWR VPWR hold723/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3526_ _3526_/A _3714_/B VGND VGND VPWR VPWR _5187_/A sky130_fd_sc_hd__nor2_8
Xhold734 _5474_/X VGND VGND VPWR VPWR _7041_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6314_ _6604_/Q _5980_/Y _6036_/X _6519_/Q _6298_/X VGND VGND VPWR VPWR _6315_/D
+ sky130_fd_sc_hd__a221o_1
Xhold745 _7033_/Q VGND VGND VPWR VPWR hold745/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold756 _4128_/X VGND VGND VPWR VPWR _6595_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold767 _6755_/Q VGND VGND VPWR VPWR hold767/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold778 _4251_/X VGND VGND VPWR VPWR _6705_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6245_ _6245_/A1 _6319_/S _6243_/X _6244_/X VGND VGND VPWR VPWR _7183_/D sky130_fd_sc_hd__o22a_1
X_3457_ _7022_/Q _5448_/A _4282_/A _6735_/Q VGND VGND VPWR VPWR _3457_/X sky130_fd_sc_hd__a22o_1
Xhold789 _6688_/Q VGND VGND VPWR VPWR hold789/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6176_ _7141_/Q _6023_/B _6204_/A2 _7024_/Q VGND VGND VPWR VPWR _6176_/X sky130_fd_sc_hd__a22o_1
XFILLER_162_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3388_ _7032_/Q _5457_/A _5259_/A _6856_/Q _3387_/X VGND VGND VPWR VPWR _3392_/B
+ sky130_fd_sc_hd__a221o_1
Xhold1401 _6629_/Q VGND VGND VPWR VPWR hold1401/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1412 _6640_/Q VGND VGND VPWR VPWR hold1412/X sky130_fd_sc_hd__dlygate4sd3_1
X_5127_ _5148_/A _5127_/B _5127_/C VGND VGND VPWR VPWR _5159_/B sky130_fd_sc_hd__nor3_1
Xhold1423 _6449_/Q VGND VGND VPWR VPWR hold83/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1434 _3300_/Y VGND VGND VPWR VPWR _5421_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1445 _7191_/Q VGND VGND VPWR VPWR _6351_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1456 _6492_/Q VGND VGND VPWR VPWR hold1456/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1467 _3725_/X VGND VGND VPWR VPWR _6784_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5058_ _4931_/A _4951_/B _4846_/D VGND VGND VPWR VPWR _5059_/C sky130_fd_sc_hd__o21a_1
XFILLER_55_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1478 _6646_/Q VGND VGND VPWR VPWR _4188_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1489 _3860_/X VGND VGND VPWR VPWR _6452_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4009_ _5552_/A0 hold737/X _4009_/S VGND VGND VPWR VPWR _4009_/X sky130_fd_sc_hd__mux2_1
XTAP_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold50 hold50/A VGND VGND VPWR VPWR hold50/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 hold61/A VGND VGND VPWR VPWR hold61/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 hold72/A VGND VGND VPWR VPWR hold72/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 hold83/A VGND VGND VPWR VPWR hold83/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 hold94/A VGND VGND VPWR VPWR hold94/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_35_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_674 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_3 _3966_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4360_ _4360_/A _4360_/B VGND VGND VPWR VPWR _4462_/B sky130_fd_sc_hd__or2_1
XFILLER_125_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3311_ _3340_/B _3530_/B VGND VGND VPWR VPWR _5349_/A sky130_fd_sc_hd__nor2_8
XFILLER_125_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4291_ hold44/X hold253/X _4293_/S VGND VGND VPWR VPWR _4291_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6030_ _6033_/A _6040_/B _6030_/C VGND VGND VPWR VPWR _6030_/X sky130_fd_sc_hd__and3_4
X_3242_ hold91/X _3252_/B VGND VGND VPWR VPWR hold92/A sky130_fd_sc_hd__and2_1
XFILLER_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6932_ _7136_/CLK _6932_/D fanout521/X VGND VGND VPWR VPWR _6932_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_47_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6863_ _7079_/CLK _6863_/D fanout516/X VGND VGND VPWR VPWR _6863_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5814_ _6847_/Q _5691_/Y _5804_/X _5813_/X _6318_/S VGND VGND VPWR VPWR _5814_/X
+ sky130_fd_sc_hd__o221a_2
X_6794_ _7209_/CLK _6794_/D fanout484/X VGND VGND VPWR VPWR _6794_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_167_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5745_ _6924_/Q _5955_/A2 _5693_/X _6900_/Q _5744_/X VGND VGND VPWR VPWR _5750_/B
+ sky130_fd_sc_hd__a221o_1
X_5676_ _7152_/Q _5703_/C _5699_/C VGND VGND VPWR VPWR _5676_/X sky130_fd_sc_hd__and3_4
XFILLER_148_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4627_ _4986_/A _5115_/B _4627_/C _5177_/A VGND VGND VPWR VPWR _4634_/A sky130_fd_sc_hd__or4_1
XFILLER_163_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold520 _6929_/Q VGND VGND VPWR VPWR hold520/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold531 _4335_/X VGND VGND VPWR VPWR _6775_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4558_ _4802_/B _4609_/B VGND VGND VPWR VPWR _4778_/B sky130_fd_sc_hd__nor2_2
XFILLER_190_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold542 _7053_/Q VGND VGND VPWR VPWR hold542/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold553 _5198_/X VGND VGND VPWR VPWR _6802_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold564 _7197_/Q VGND VGND VPWR VPWR hold564/X sky130_fd_sc_hd__dlygate4sd3_1
X_3509_ _7099_/Q _5535_/A _5571_/A _7131_/Q _3508_/X VGND VGND VPWR VPWR _3515_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold575 _7114_/Q VGND VGND VPWR VPWR hold575/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold586 _4146_/X VGND VGND VPWR VPWR _6610_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4489_ _4489_/A _4932_/A _5023_/B VGND VGND VPWR VPWR _4489_/X sky130_fd_sc_hd__or3_1
XFILLER_104_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold597 _6949_/Q VGND VGND VPWR VPWR hold597/X sky130_fd_sc_hd__dlygate4sd3_1
X_6228_ _6731_/Q _5997_/Y _6015_/X _6660_/Q VGND VGND VPWR VPWR _6228_/X sky130_fd_sc_hd__a22o_1
XFILLER_131_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6159_ _6919_/Q wire412/X _6024_/D _6943_/Q VGND VGND VPWR VPWR _6159_/X sky130_fd_sc_hd__a22o_1
Xhold1220 _6741_/Q VGND VGND VPWR VPWR _4295_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_530 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1231 _5260_/X VGND VGND VPWR VPWR _6850_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1242 _6882_/Q VGND VGND VPWR VPWR _5296_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1253 _4041_/X VGND VGND VPWR VPWR _6531_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1264 _4130_/X VGND VGND VPWR VPWR _6596_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1275 _6521_/Q VGND VGND VPWR VPWR _4029_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1286 _4265_/X VGND VGND VPWR VPWR _6716_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1297 _6506_/Q VGND VGND VPWR VPWR _4011_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput140 wb_dat_i[17] VGND VGND VPWR VPWR _6367_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput151 wb_dat_i[27] VGND VGND VPWR VPWR _6373_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput162 wb_dat_i[8] VGND VGND VPWR VPWR _6364_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3860_ hold1/A _3860_/A1 _3866_/S VGND VGND VPWR VPWR _3860_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3791_ _3791_/A _3917_/A VGND VGND VPWR VPWR _3791_/Y sky130_fd_sc_hd__nor2_1
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5530_ _5530_/A0 _6393_/A0 _5534_/S VGND VGND VPWR VPWR _5530_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5461_ hold36/X hold275/X _5465_/S VGND VGND VPWR VPWR _5461_/X sky130_fd_sc_hd__mux2_1
X_4412_ _4341_/X _4538_/B _4588_/A VGND VGND VPWR VPWR _4435_/A sky130_fd_sc_hd__a21o_1
X_7200_ _7200_/CLK _7200_/D fanout529/X VGND VGND VPWR VPWR _7200_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5392_ _5587_/A0 hold836/X _5393_/S VGND VGND VPWR VPWR _5392_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7131_ _7139_/CLK _7131_/D fanout518/X VGND VGND VPWR VPWR _7131_/Q sky130_fd_sc_hd__dfrtp_4
X_4343_ _4846_/B _4570_/D VGND VGND VPWR VPWR _4596_/A sky130_fd_sc_hd__nand2_2
XFILLER_113_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7062_ _7075_/CLK _7062_/D fanout515/X VGND VGND VPWR VPWR _7062_/Q sky130_fd_sc_hd__dfrtp_1
X_4274_ hold146/X hold36/X _4275_/S VGND VGND VPWR VPWR _4274_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6013_ _6040_/A _6020_/C _6040_/C VGND VGND VPWR VPWR _6027_/C sky130_fd_sc_hd__and3_1
X_3225_ _6917_/Q VGND VGND VPWR VPWR _3225_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6915_ _7128_/CLK _6915_/D fanout514/X VGND VGND VPWR VPWR _6915_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_35_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6846_ _7068_/CLK _6846_/D fanout505/X VGND VGND VPWR VPWR _6846_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_167_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6777_ _3937_/A1 _6777_/D fanout529/X VGND VGND VPWR VPWR _6777_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_167_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3989_ hold140/X hold127/X _3991_/S VGND VGND VPWR VPWR _3989_/X sky130_fd_sc_hd__mux2_1
XFILLER_167_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5728_ _5728_/A _5728_/B _5728_/C _5728_/D VGND VGND VPWR VPWR _5728_/X sky130_fd_sc_hd__or4_1
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5659_ _5938_/B _5699_/B _5706_/C VGND VGND VPWR VPWR _5659_/X sky130_fd_sc_hd__and3_4
XFILLER_163_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold350 _4101_/X VGND VGND VPWR VPWR _6572_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 _6638_/Q VGND VGND VPWR VPWR hold361/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold372 _5537_/X VGND VGND VPWR VPWR _7096_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 _6709_/Q VGND VGND VPWR VPWR hold383/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 _5570_/X VGND VGND VPWR VPWR _7126_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1050 _5368_/X VGND VGND VPWR VPWR _6946_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1061 _6726_/Q VGND VGND VPWR VPWR _4277_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1072 _5572_/X VGND VGND VPWR VPWR _7127_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1083 _6858_/Q VGND VGND VPWR VPWR _5269_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1094 _7135_/Q VGND VGND VPWR VPWR _5581_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_201 _5655_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_212 _6613_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_223 _5331_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_234 _5496_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_245 _5655_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_256 _5581_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4961_ _4961_/A _4961_/B VGND VGND VPWR VPWR _4962_/B sky130_fd_sc_hd__nor2_1
XFILLER_17_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6700_ _7200_/CLK _6700_/D _6348_/B VGND VGND VPWR VPWR _6700_/Q sky130_fd_sc_hd__dfrtp_4
X_3912_ _3914_/A1 _3868_/A _6541_/Q _3834_/B _3912_/B1 VGND VGND VPWR VPWR _6542_/D
+ sky130_fd_sc_hd__a41o_1
X_4892_ _4454_/Y _4871_/Y _5049_/C _4878_/X _4891_/X VGND VGND VPWR VPWR _4892_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_189_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6631_ _7196_/CLK _6631_/D VGND VGND VPWR VPWR _6631_/Q sky130_fd_sc_hd__dfxtp_1
X_3843_ _3794_/B _3890_/A _3842_/Y _6541_/Q VGND VGND VPWR VPWR _6458_/D sky130_fd_sc_hd__a211oi_1
XFILLER_149_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3774_ _6596_/Q _4129_/A _4312_/A _6756_/Q _3773_/X VGND VGND VPWR VPWR _3781_/A
+ sky130_fd_sc_hd__a221o_1
X_6562_ _7182_/CLK _6562_/D fanout499/X VGND VGND VPWR VPWR _6562_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_164_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5513_ _5573_/A0 hold803/X _5519_/S VGND VGND VPWR VPWR _5513_/X sky130_fd_sc_hd__mux2_1
X_6493_ _6759_/CLK _6493_/D fanout488/X VGND VGND VPWR VPWR _6493_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_145_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5444_ _5567_/A0 hold707/X _5447_/S VGND VGND VPWR VPWR _5444_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5375_ _5579_/A0 hold514/X _5375_/S VGND VGND VPWR VPWR _5375_/X sky130_fd_sc_hd__mux2_1
X_7114_ _7134_/CLK _7114_/D fanout525/X VGND VGND VPWR VPWR _7114_/Q sky130_fd_sc_hd__dfrtp_4
X_4326_ hold301/X _5555_/A0 _4329_/S VGND VGND VPWR VPWR _4326_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4257_ hold687/X _5534_/A1 _4257_/S VGND VGND VPWR VPWR _4257_/X sky130_fd_sc_hd__mux2_1
X_7045_ _7108_/CLK _7045_/D fanout523/X VGND VGND VPWR VPWR _7045_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3208_ _7053_/Q VGND VGND VPWR VPWR _3208_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4188_ _4188_/A0 _3373_/X _4188_/S VGND VGND VPWR VPWR _6646_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6829_ _7138_/CLK _6829_/D fanout524/X VGND VGND VPWR VPWR _6829_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold180 _4116_/X VGND VGND VPWR VPWR _6584_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 _6813_/Q VGND VGND VPWR VPWR hold191/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_747 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3490_ hold95/X _3525_/B VGND VGND VPWR VPWR _4300_/A sky130_fd_sc_hd__nor2_4
XFILLER_6_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5160_ _5160_/A _5160_/B _5160_/C VGND VGND VPWR VPWR _5160_/X sky130_fd_sc_hd__or3_1
XFILLER_69_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4111_ hold96/X _4111_/B _6407_/B hold13/X VGND VGND VPWR VPWR hold97/A sky130_fd_sc_hd__or4_4
X_5091_ _4516_/B _4729_/Y _4988_/B _4627_/C _4635_/Y VGND VGND VPWR VPWR _5092_/D
+ sky130_fd_sc_hd__a2111o_1
XFILLER_96_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4042_ _5531_/A1 hold958/X _4045_/S VGND VGND VPWR VPWR _4042_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5993_ _7095_/Q _6338_/B1 _5992_/X _6930_/Q _5990_/X VGND VGND VPWR VPWR _6012_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_52_558 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4944_ _4944_/A _4944_/B VGND VGND VPWR VPWR _4944_/X sky130_fd_sc_hd__or2_1
XFILLER_178_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4875_ _4964_/A _4875_/B VGND VGND VPWR VPWR _4875_/X sky130_fd_sc_hd__or2_1
X_6614_ _6708_/CLK _6614_/D fanout494/X VGND VGND VPWR VPWR _6614_/Q sky130_fd_sc_hd__dfstp_2
X_3826_ hold53/A hold25/A hold64/A VGND VGND VPWR VPWR _3826_/X sky130_fd_sc_hd__a21o_1
XFILLER_20_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6545_ _3927_/A1 _6545_/D _6433_/X VGND VGND VPWR VPWR _6545_/Q sky130_fd_sc_hd__dfrtp_1
X_3757_ input43/X _4068_/S _5205_/A _6807_/Q _3740_/X VGND VGND VPWR VPWR _3760_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_173_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6476_ _6825_/CLK _6476_/D fanout490/X VGND VGND VPWR VPWR _6476_/Q sky130_fd_sc_hd__dfstp_1
X_3688_ _3688_/A _3688_/B _3688_/C _3688_/D VGND VGND VPWR VPWR _3689_/B sky130_fd_sc_hd__or4_1
X_5427_ hold127/X hold154/X _5429_/S VGND VGND VPWR VPWR _5427_/X sky130_fd_sc_hd__mux2_1
Xoutput230 _6827_/Q VGND VGND VPWR VPWR mgmt_gpio_out[25] sky130_fd_sc_hd__buf_12
Xoutput241 _3925_/X VGND VGND VPWR VPWR mgmt_gpio_out[35] sky130_fd_sc_hd__buf_12
XFILLER_133_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput252 _3946_/Y VGND VGND VPWR VPWR pad_flash_clk_oeb sky130_fd_sc_hd__buf_12
XFILLER_160_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput263 _6803_/Q VGND VGND VPWR VPWR pll90_sel[2] sky130_fd_sc_hd__buf_12
Xoutput274 _6800_/Q VGND VGND VPWR VPWR pll_sel[2] sky130_fd_sc_hd__buf_12
Xoutput285 _6477_/Q VGND VGND VPWR VPWR pll_trim[19] sky130_fd_sc_hd__buf_12
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5358_ _5358_/A _5580_/B VGND VGND VPWR VPWR _5366_/S sky130_fd_sc_hd__nand2_8
Xoutput296 _6495_/Q VGND VGND VPWR VPWR pll_trim[5] sky130_fd_sc_hd__buf_12
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4309_ _6395_/A0 _4309_/A1 _4311_/S VGND VGND VPWR VPWR _4309_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5289_ _5574_/A0 _5289_/A1 hold32/X VGND VGND VPWR VPWR _5289_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7028_ _7137_/CLK _7028_/D fanout501/X VGND VGND VPWR VPWR _7028_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_28_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7159__531 VGND VGND VPWR VPWR _7159_/D _7159__531/LO sky130_fd_sc_hd__conb_1
XFILLER_75_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire357 _3280_/Y VGND VGND VPWR VPWR _5304_/A sky130_fd_sc_hd__buf_8
XFILLER_136_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout490 fanout491/X VGND VGND VPWR VPWR fanout490/X sky130_fd_sc_hd__buf_6
XFILLER_48_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4660_ _5023_/A _5023_/B VGND VGND VPWR VPWR _5016_/B sky130_fd_sc_hd__and2_2
XFILLER_30_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3611_ _6924_/Q _5340_/A hold58/A _6683_/Q VGND VGND VPWR VPWR _3611_/X sky130_fd_sc_hd__a22o_1
XFILLER_175_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4591_ _4605_/A _4621_/B _4621_/C VGND VGND VPWR VPWR _4707_/A sky130_fd_sc_hd__or3_4
XFILLER_190_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6330_ _6510_/Q _6049_/B _6021_/Y _6625_/Q _6329_/X VGND VGND VPWR VPWR _6331_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_162_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3542_ _3542_/A _3542_/B _3542_/C _3542_/D VGND VGND VPWR VPWR _3543_/C sky130_fd_sc_hd__or4_2
Xhold905 _5360_/X VGND VGND VPWR VPWR _6939_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold916 _6480_/Q VGND VGND VPWR VPWR hold916/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold927 _5518_/X VGND VGND VPWR VPWR _7080_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold938 _7008_/Q VGND VGND VPWR VPWR hold938/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_142_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3473_ _6765_/Q _3471_/Y _3472_/Y _3658_/A VGND VGND VPWR VPWR _3473_/X sky130_fd_sc_hd__a211o_1
X_6261_ _6671_/Q _6340_/A2 _6023_/D _6635_/Q _6260_/X VGND VGND VPWR VPWR _6266_/A
+ sky130_fd_sc_hd__a221o_1
Xhold949 _4308_/X VGND VGND VPWR VPWR _6752_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5212_ _5212_/A _5212_/B _5212_/C VGND VGND VPWR VPWR _5212_/X sky130_fd_sc_hd__or3_1
X_6192_ _6192_/A _6192_/B _6192_/C _6192_/D VGND VGND VPWR VPWR _6193_/C sky130_fd_sc_hd__or4_1
XFILLER_123_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5143_ _4814_/B _4653_/C _4795_/Y _4870_/B VGND VGND VPWR VPWR _5143_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_96_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1605 _7113_/Q VGND VGND VPWR VPWR hold1605/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5074_ _5021_/A _4596_/X _4665_/B VGND VGND VPWR VPWR _5074_/X sky130_fd_sc_hd__o21a_1
XFILLER_57_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4025_ _4025_/A0 _6395_/A0 _4027_/S VGND VGND VPWR VPWR _4025_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5976_ _6006_/B _6021_/A VGND VGND VPWR VPWR _6022_/A sky130_fd_sc_hd__nor2_1
XFILLER_52_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4927_ _5130_/B _4925_/X _4650_/Y VGND VGND VPWR VPWR _4928_/D sky130_fd_sc_hd__o21a_1
XFILLER_33_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4858_ _4424_/Y _5035_/B _4694_/X _4857_/X VGND VGND VPWR VPWR _4858_/X sky130_fd_sc_hd__o211a_1
XFILLER_21_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3809_ hold46/A _6468_/Q _6467_/Q _3821_/S VGND VGND VPWR VPWR _3811_/S sky130_fd_sc_hd__nand4_1
XFILLER_165_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4789_ _5002_/A _4802_/A _5076_/B _5108_/A VGND VGND VPWR VPWR _4983_/C sky130_fd_sc_hd__o22ai_1
XFILLER_4_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6528_ _7207_/CLK _6528_/D fanout484/X VGND VGND VPWR VPWR _6528_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_180_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6459_ _3945_/A1 _6459_/D _6414_/X VGND VGND VPWR VPWR _6459_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_106_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5830_ _7072_/Q _5678_/X _5703_/X _6856_/Q _5829_/X VGND VGND VPWR VPWR _5835_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_61_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5761_ _6997_/Q _5656_/X _5671_/X _7061_/Q VGND VGND VPWR VPWR _5761_/X sky130_fd_sc_hd__a22o_1
X_4712_ _5018_/A _4814_/B _5018_/C VGND VGND VPWR VPWR _4713_/D sky130_fd_sc_hd__or3_1
X_5692_ _6858_/Q _5688_/X _5689_/X _6970_/Q _5690_/X VGND VGND VPWR VPWR _5692_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_187_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4643_ _4569_/B _5024_/A _4642_/X _4847_/A _4530_/B VGND VGND VPWR VPWR _4643_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_162_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap410 _6015_/X VGND VGND VPWR VPWR _6024_/C sky130_fd_sc_hd__buf_12
X_4574_ _5036_/A _4609_/B _4981_/C VGND VGND VPWR VPWR _4574_/Y sky130_fd_sc_hd__nor3_1
Xhold702 _5489_/X VGND VGND VPWR VPWR _7054_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 _6765_/Q VGND VGND VPWR VPWR hold713/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap421 _5672_/X VGND VGND VPWR VPWR _5955_/A2 sky130_fd_sc_hd__buf_12
XFILLER_162_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold724 _5429_/X VGND VGND VPWR VPWR _7001_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6313_ _6609_/Q _6326_/A2 _6021_/Y _6624_/Q _6312_/X VGND VGND VPWR VPWR _6315_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3525_ _3525_/A _3525_/B VGND VGND VPWR VPWR _4046_/A sky130_fd_sc_hd__nor2_4
Xhold735 _6990_/Q VGND VGND VPWR VPWR hold735/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold746 _5465_/X VGND VGND VPWR VPWR _7033_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold757 _7081_/Q VGND VGND VPWR VPWR hold757/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold768 _4311_/X VGND VGND VPWR VPWR _6755_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold779 _7009_/Q VGND VGND VPWR VPWR hold779/X sky130_fd_sc_hd__dlygate4sd3_1
X_6244_ _7182_/Q _5592_/Y _5650_/Y VGND VGND VPWR VPWR _6244_/X sky130_fd_sc_hd__o21ba_1
XFILLER_89_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3456_ _3507_/B _3525_/B VGND VGND VPWR VPWR _4282_/A sky130_fd_sc_hd__nor2_4
XFILLER_130_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3387_ _6992_/Q _5412_/A hold78/A _7048_/Q VGND VGND VPWR VPWR _3387_/X sky130_fd_sc_hd__a22o_1
X_6175_ _6992_/Q _6203_/A2 _6022_/D _7125_/Q _6174_/X VGND VGND VPWR VPWR _6180_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_97_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1402 _6627_/Q VGND VGND VPWR VPWR hold1402/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1413 _6639_/Q VGND VGND VPWR VPWR hold1413/X sky130_fd_sc_hd__dlygate4sd3_1
X_5126_ _5126_/A _5126_/B _5126_/C _4945_/X VGND VGND VPWR VPWR _5160_/B sky130_fd_sc_hd__or4b_1
Xhold1424 _6650_/Q VGND VGND VPWR VPWR _4193_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1435 _6489_/Q VGND VGND VPWR VPWR _3991_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1446 _6938_/Q VGND VGND VPWR VPWR hold1446/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1457 _3995_/X VGND VGND VPWR VPWR _6492_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1468 _6788_/Q VGND VGND VPWR VPWR _3449_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5057_ _4932_/A _5023_/B _4675_/A _5056_/X _4503_/C VGND VGND VPWR VPWR _5123_/B
+ sky130_fd_sc_hd__o311a_1
Xhold1479 _6631_/Q VGND VGND VPWR VPWR _4171_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_55_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4008_ _5587_/A0 hold920/X _4009_/S VGND VGND VPWR VPWR _4008_/X sky130_fd_sc_hd__mux2_1
XTAP_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5959_ _6620_/Q _5667_/X _5683_/X _6615_/Q _5958_/X VGND VGND VPWR VPWR _5967_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_139_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold40 hold40/A VGND VGND VPWR VPWR hold40/X sky130_fd_sc_hd__buf_6
Xhold51 hold51/A VGND VGND VPWR VPWR hold51/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold62 hold62/A VGND VGND VPWR VPWR hold62/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 hold73/A VGND VGND VPWR VPWR hold73/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 hold84/A VGND VGND VPWR VPWR hold84/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 hold95/A VGND VGND VPWR VPWR hold95/X sky130_fd_sc_hd__buf_8
XFILLER_152_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_4 _5520_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3310_ hold68/X _3334_/A VGND VGND VPWR VPWR _5367_/A sky130_fd_sc_hd__nor2_8
XFILLER_98_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4290_ _5459_/A0 hold327/X _4293_/S VGND VGND VPWR VPWR _4290_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3241_ _6473_/Q _6472_/Q _6471_/Q VGND VGND VPWR VPWR _3791_/A sky130_fd_sc_hd__or3_4
XFILLER_98_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6931_ _6931_/CLK _6931_/D fanout517/X VGND VGND VPWR VPWR _6931_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6862_ _7123_/CLK _6862_/D _6407_/A VGND VGND VPWR VPWR _6862_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_34_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5813_ _5813_/A _5813_/B _5813_/C _5813_/D VGND VGND VPWR VPWR _5813_/X sky130_fd_sc_hd__or4_1
XFILLER_179_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6793_ _7209_/CLK _6793_/D fanout484/X VGND VGND VPWR VPWR _6793_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_50_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5744_ _7052_/Q _5699_/X _5743_/X _5691_/B VGND VGND VPWR VPWR _5744_/X sky130_fd_sc_hd__a22o_1
XFILLER_148_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5675_ _5938_/B _5706_/B _5706_/C VGND VGND VPWR VPWR _5675_/X sky130_fd_sc_hd__and3_4
Xclkbuf_leaf_72_csclk _6753_/CLK VGND VGND VPWR VPWR _6760_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_108_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4626_ _5177_/A VGND VGND VPWR VPWR _4626_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold510 _6857_/Q VGND VGND VPWR VPWR hold510/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold521 _5348_/X VGND VGND VPWR VPWR _6929_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4557_ _4605_/A _4793_/B _4802_/C VGND VGND VPWR VPWR _4609_/B sky130_fd_sc_hd__or3_2
Xhold532 _6887_/Q VGND VGND VPWR VPWR hold532/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold543 _5488_/X VGND VGND VPWR VPWR _7053_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 _6897_/Q VGND VGND VPWR VPWR hold554/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3508_ _6486_/Q _3983_/A _4034_/A _6530_/Q VGND VGND VPWR VPWR _3508_/X sky130_fd_sc_hd__a22o_2
XFILLER_1_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold565 _3967_/X VGND VGND VPWR VPWR hold565/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4488_ _4759_/A _5060_/A VGND VGND VPWR VPWR _4847_/A sky130_fd_sc_hd__nand2_2
Xhold576 _5557_/X VGND VGND VPWR VPWR _7114_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold587 _6927_/Q VGND VGND VPWR VPWR hold587/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold598 _5371_/X VGND VGND VPWR VPWR _6949_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6227_ _6506_/Q _6049_/B _6006_/Y _6751_/Q _6222_/X VGND VGND VPWR VPWR _6232_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_104_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3439_ input8/X _3295_/Y _3340_/Y input25/X VGND VGND VPWR VPWR _3439_/X sky130_fd_sc_hd__a22o_2
XFILLER_58_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6158_ _7116_/Q _6322_/B1 _6030_/X _6999_/Q _6157_/X VGND VGND VPWR VPWR _6168_/B
+ sky130_fd_sc_hd__a221o_1
Xhold1210 _4105_/X VGND VGND VPWR VPWR _6574_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1221 _4295_/X VGND VGND VPWR VPWR _6741_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_10_csclk _6820_/CLK VGND VGND VPWR VPWR _6679_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_85_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1232 _6954_/Q VGND VGND VPWR VPWR _5377_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5109_ _5109_/A _5109_/B _5109_/C _5109_/D VGND VGND VPWR VPWR _5110_/C sky130_fd_sc_hd__or4_1
Xhold1243 _5296_/X VGND VGND VPWR VPWR _6882_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6089_ _7012_/Q _5998_/Y _6023_/C _6868_/Q _6088_/X VGND VGND VPWR VPWR _6094_/C
+ sky130_fd_sc_hd__a221o_1
Xhold1254 _6621_/Q VGND VGND VPWR VPWR _4160_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1265 _7082_/Q VGND VGND VPWR VPWR _5521_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1276 _4029_/X VGND VGND VPWR VPWR _6521_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1287 _6474_/Q VGND VGND VPWR VPWR _3968_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1298 _4011_/X VGND VGND VPWR VPWR _6506_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_25_csclk _6882_/CLK VGND VGND VPWR VPWR _7139_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_53_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput130 wb_adr_i[9] VGND VGND VPWR VPWR _4339_/A sky130_fd_sc_hd__clkbuf_1
Xinput141 wb_dat_i[18] VGND VGND VPWR VPWR _6369_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput152 wb_dat_i[28] VGND VGND VPWR VPWR _6376_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput163 wb_dat_i[9] VGND VGND VPWR VPWR _6366_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3790_ _3790_/A _3790_/B _3790_/C _3790_/D VGND VGND VPWR VPWR _3790_/X sky130_fd_sc_hd__or4_4
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5460_ _5583_/A0 hold305/X _5465_/S VGND VGND VPWR VPWR _5460_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4411_ _4758_/A _5001_/A VGND VGND VPWR VPWR _4445_/A sky130_fd_sc_hd__nand2_1
X_5391_ _5586_/A0 _5391_/A1 _5393_/S VGND VGND VPWR VPWR _5391_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7130_ _7130_/CLK _7130_/D fanout521/X VGND VGND VPWR VPWR _7130_/Q sky130_fd_sc_hd__dfrtp_4
X_4342_ _4588_/A _4605_/A _4621_/B VGND VGND VPWR VPWR _4819_/C sky130_fd_sc_hd__and3_2
XFILLER_98_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7061_ _7138_/CLK _7061_/D fanout521/X VGND VGND VPWR VPWR _7061_/Q sky130_fd_sc_hd__dfrtp_4
X_4273_ hold221/X hold44/X _4275_/S VGND VGND VPWR VPWR _4273_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6012_ _6012_/A _6012_/B _6012_/C _6012_/D VGND VGND VPWR VPWR _6045_/B sky130_fd_sc_hd__or4_1
X_3224_ _6925_/Q VGND VGND VPWR VPWR _3224_/Y sky130_fd_sc_hd__inv_2
.ends

