magic
tech sky130A
magscale 1 2
timestamp 1695840358
<< metal2 >>
rect 27498 953270 27558 953726
rect 29498 953270 29558 953726
rect 34360 953270 34416 953726
rect 34912 953270 34968 953726
rect 35556 953270 35612 953726
rect 36200 953270 36256 953726
rect 38040 953270 38096 953726
rect 38592 953270 38648 953726
rect 39236 953270 39292 953726
rect 39880 953270 39936 953726
rect 42364 953270 42420 953726
rect 42916 953270 42972 953726
rect 43560 953270 43616 953726
rect 44204 953270 44260 953726
rect 44677 953270 44891 953726
rect 45400 953270 45456 953726
rect 46560 953270 46688 953726
rect 47240 953270 47296 953726
rect 49080 953270 49136 953726
rect 78698 953270 78758 953726
rect 80698 953270 80758 953726
rect 85760 953270 85816 953726
rect 86312 953270 86368 953726
rect 86956 953270 87012 953726
rect 87600 953270 87656 953726
rect 89440 953270 89496 953726
rect 89992 953270 90048 953726
rect 90636 953270 90692 953726
rect 91280 953270 91336 953726
rect 93764 953270 93820 953726
rect 94316 953270 94372 953726
rect 94960 953270 95016 953726
rect 95604 953270 95660 953726
rect 96077 953270 96291 953726
rect 96800 953270 96856 953726
rect 97960 953270 98088 953726
rect 98640 953270 98696 953726
rect 100480 953270 100536 953726
rect 129898 953270 129958 953726
rect 131898 953270 131958 953726
rect 137160 953270 137216 953726
rect 137712 953270 137768 953726
rect 138356 953270 138412 953726
rect 139000 953270 139056 953726
rect 140840 953270 140896 953726
rect 141392 953270 141448 953726
rect 142036 953270 142092 953726
rect 142680 953270 142736 953726
rect 145164 953270 145220 953726
rect 145716 953270 145772 953726
rect 146360 953270 146416 953726
rect 147004 953270 147060 953726
rect 147477 953270 147691 953726
rect 148200 953270 148256 953726
rect 149360 953270 149488 953726
rect 150040 953270 150096 953726
rect 151880 953270 151936 953726
rect 181098 953270 181158 953726
rect 183098 953270 183158 953726
rect 188560 953270 188616 953726
rect 189112 953270 189168 953726
rect 189756 953270 189812 953726
rect 190400 953270 190456 953726
rect 192240 953270 192296 953726
rect 192792 953270 192848 953726
rect 193436 953270 193492 953726
rect 194080 953270 194136 953726
rect 196564 953270 196620 953726
rect 197116 953270 197172 953726
rect 197760 953270 197816 953726
rect 198404 953270 198460 953726
rect 198877 953270 199091 953726
rect 199600 953270 199656 953726
rect 200760 953270 200888 953726
rect 201440 953270 201496 953726
rect 203280 953270 203336 953726
rect 232298 953270 232358 953726
rect 234298 953270 234358 953726
rect 240160 953270 240216 953726
rect 240712 953270 240768 953726
rect 241356 953270 241412 953726
rect 242000 953270 242056 953726
rect 243840 953270 243896 953726
rect 244392 953270 244448 953726
rect 245036 953270 245092 953726
rect 245680 953270 245736 953726
rect 248164 953270 248220 953726
rect 248716 953270 248772 953726
rect 249360 953270 249416 953726
rect 250004 953270 250060 953726
rect 250477 953270 250691 953726
rect 251200 953270 251256 953726
rect 252360 953270 252488 953726
rect 253040 953270 253096 953726
rect 254880 953270 254936 953726
rect 336698 953270 336758 953726
rect 338698 953270 338758 953726
rect 341960 953270 342016 953726
rect 342512 953270 342568 953726
rect 343156 953270 343212 953726
rect 343800 953270 343856 953726
rect 345640 953270 345696 953726
rect 346192 953270 346248 953726
rect 346836 953270 346892 953726
rect 347480 953270 347536 953726
rect 349964 953270 350020 953726
rect 350516 953270 350572 953726
rect 351160 953270 351216 953726
rect 351804 953270 351860 953726
rect 352277 953270 352491 953726
rect 353000 953270 353056 953726
rect 354160 953270 354288 953726
rect 354840 953270 354896 953726
rect 356680 953270 356736 953726
rect 425698 953270 425758 953726
rect 427698 953270 427758 953726
rect 430960 953270 431016 953726
rect 431512 953270 431568 953726
rect 432156 953270 432212 953726
rect 432800 953270 432856 953726
rect 434640 953270 434696 953726
rect 435192 953270 435248 953726
rect 435836 953270 435892 953726
rect 436480 953270 436536 953726
rect 438964 953270 439020 953726
rect 439516 953270 439572 953726
rect 440160 953270 440216 953726
rect 440804 953270 440860 953726
rect 441277 953270 441491 953726
rect 442000 953270 442056 953726
rect 443160 953270 443288 953726
rect 443840 953270 443896 953726
rect 445680 953270 445736 953726
rect 476898 953270 476958 953726
rect 478898 953270 478958 953726
rect 482360 953270 482416 953726
rect 482912 953270 482968 953726
rect 483556 953270 483612 953726
rect 484200 953270 484256 953726
rect 486040 953270 486096 953726
rect 486592 953270 486648 953726
rect 487236 953270 487292 953726
rect 487880 953270 487936 953726
rect 490364 953270 490420 953726
rect 490916 953270 490972 953726
rect 491560 953270 491616 953726
rect 492204 953270 492260 953726
rect 492677 953270 492891 953726
rect 493400 953270 493456 953726
rect 494560 953270 494688 953726
rect 495240 953270 495296 953726
rect 497080 953270 497136 953726
rect 576298 953270 576358 953726
rect 578298 953270 578358 953726
rect 584160 953270 584216 953726
rect 584712 953270 584768 953726
rect 585356 953270 585412 953726
rect 586000 953270 586056 953726
rect 587840 953270 587896 953726
rect 588392 953270 588448 953726
rect 589036 953270 589092 953726
rect 589680 953270 589736 953726
rect 592164 953270 592220 953726
rect 592716 953270 592772 953726
rect 593360 953270 593416 953726
rect 594004 953270 594060 953726
rect 594477 953270 594691 953726
rect 595200 953270 595256 953726
rect 596360 953270 596488 953726
rect 597040 953270 597096 953726
rect 598880 953270 598936 953726
rect 99576 -400 99632 56
rect 110164 -400 110220 56
rect 145190 -400 145246 56
rect 147030 -400 147086 56
rect 147638 -400 147766 56
rect 148870 -400 148926 56
rect 149435 -400 149649 56
rect 150066 -400 150122 56
rect 150710 -400 150766 56
rect 151354 -400 151410 56
rect 151906 -400 151962 56
rect 154390 -400 154446 56
rect 155034 -400 155090 56
rect 155678 -400 155734 56
rect 156230 -400 156286 56
rect 158070 -400 158126 56
rect 158714 -400 158770 56
rect 159358 -400 159414 56
rect 159910 -400 159966 56
rect 160580 -400 160632 56
rect 163791 -400 163843 56
rect 253790 -400 253846 56
rect 255630 -400 255686 56
rect 256238 -400 256366 56
rect 257470 -400 257526 56
rect 258035 -400 258249 56
rect 258666 -400 258722 56
rect 259310 -400 259366 56
rect 259954 -400 260010 56
rect 260506 -400 260562 56
rect 262990 -400 263046 56
rect 263634 -400 263690 56
rect 264278 -400 264334 56
rect 264830 -400 264886 56
rect 266670 -400 266726 56
rect 267314 -400 267370 56
rect 267958 -400 268014 56
rect 268510 -400 268566 56
rect 269180 -400 269232 56
rect 273360 -400 273412 56
rect 308590 -400 308646 56
rect 310430 -400 310486 56
rect 311038 -400 311166 56
rect 312270 -400 312326 56
rect 312835 -400 313049 56
rect 313466 -400 313522 56
rect 314110 -400 314166 56
rect 314754 -400 314810 56
rect 315306 -400 315362 56
rect 317790 -400 317846 56
rect 318434 -400 318490 56
rect 319078 -400 319134 56
rect 319630 -400 319686 56
rect 321470 -400 321526 56
rect 322114 -400 322170 56
rect 322758 -400 322814 56
rect 323310 -400 323366 56
rect 323980 -400 324032 56
rect 328165 -400 328217 56
rect 363390 -400 363446 56
rect 365230 -400 365286 56
rect 365838 -400 365966 56
rect 367070 -400 367126 56
rect 367635 -400 367849 56
rect 368266 -400 368322 56
rect 368910 -400 368966 56
rect 369554 -400 369610 56
rect 370106 -400 370162 56
rect 372590 -400 372646 56
rect 373234 -400 373290 56
rect 373878 -400 373934 56
rect 374430 -400 374486 56
rect 376270 -400 376326 56
rect 376914 -400 376970 56
rect 377558 -400 377614 56
rect 378110 -400 378166 56
rect 378780 -400 378832 56
rect 382978 -400 383030 56
rect 418190 -400 418246 56
rect 420030 -400 420086 56
rect 420638 -400 420766 56
rect 421870 -400 421926 56
rect 422435 -400 422649 56
rect 423066 -400 423122 56
rect 423710 -400 423766 56
rect 424354 -400 424410 56
rect 424906 -400 424962 56
rect 427390 -400 427446 56
rect 428034 -400 428090 56
rect 428678 -400 428734 56
rect 429230 -400 429286 56
rect 431070 -400 431126 56
rect 431714 -400 431770 56
rect 432358 -400 432414 56
rect 432910 -400 432966 56
rect 433580 -400 433632 56
rect 437778 -400 437830 56
rect 472990 -400 473046 56
rect 474830 -400 474886 56
rect 475438 -400 475566 56
rect 476670 -400 476726 56
rect 477235 -400 477449 56
rect 477866 -400 477922 56
rect 478510 -400 478566 56
rect 479154 -400 479210 56
rect 479706 -400 479762 56
rect 482190 -400 482246 56
rect 482834 -400 482890 56
rect 483478 -400 483534 56
rect 484030 -400 484086 56
rect 485870 -400 485926 56
rect 486514 -400 486570 56
rect 487158 -400 487214 56
rect 487710 -400 487766 56
rect 488380 -400 488432 56
rect 492635 -400 492687 56
rect 605082 -400 605134 56
rect 605306 -400 605358 56
rect 605530 -400 605582 56
rect 605754 -400 605806 56
rect 605978 -400 606030 56
rect 606202 -400 606254 56
rect 606426 -400 606478 56
rect 606650 -400 606702 56
rect 606874 -400 606926 56
rect 607098 -400 607150 56
rect 607322 -400 607374 56
rect 607546 -400 607598 56
rect 607770 -400 607822 56
rect 607994 -400 608046 56
rect 608218 -400 608270 56
rect 608442 -400 608494 56
rect 608666 -400 608718 56
rect 608890 -400 608942 56
rect 609114 -400 609166 56
rect 609338 -400 609390 56
rect 609562 -400 609614 56
rect 609786 -400 609838 56
rect 610010 -400 610062 56
rect 610234 -400 610286 56
rect 610458 -400 610510 56
rect 610682 -400 610734 56
rect 610906 -400 610958 56
rect 611130 -400 611182 56
rect 611354 -400 611406 56
rect 611578 -400 611630 56
rect 611802 -400 611854 56
rect 612026 -400 612078 56
<< metal3 >>
rect 291362 953266 296142 953726
rect 301342 953266 306122 953726
rect 533562 953266 538342 953726
rect 543542 953266 548322 953726
rect 633266 929006 633726 929068
rect -400 927072 60 927142
rect 633266 927006 633726 927068
rect -400 925232 60 925302
rect 633266 925104 633726 925174
rect -400 924560 60 924688
rect 633266 924552 633726 924622
rect 633266 923908 633726 923978
rect -400 923392 60 923462
rect 633266 923264 633726 923334
rect -400 922677 60 922891
rect -400 922196 60 922266
rect -400 921552 60 921622
rect 633266 921424 633726 921494
rect -400 920908 60 920978
rect 633266 920872 633726 920942
rect -400 920356 60 920426
rect 633266 920228 633726 920298
rect 633266 919584 633726 919654
rect -400 917872 60 917942
rect -400 917228 60 917298
rect 633266 917100 633726 917170
rect -400 916584 60 916654
rect 633266 916548 633726 916618
rect -400 916032 60 916102
rect 633266 915904 633726 915974
rect 633266 915260 633726 915330
rect 633266 914635 633726 914849
rect -400 914192 60 914262
rect 633266 914064 633726 914134
rect -400 913548 60 913618
rect -400 912904 60 912974
rect 633266 912838 633726 912966
rect -400 912352 60 912422
rect 633266 912224 633726 912294
rect 633266 910384 633726 910454
rect -400 906644 60 906704
rect -400 904644 60 904704
rect -400 880014 60 884804
rect -400 875054 60 879716
rect -400 869964 60 874764
rect -400 837742 60 842522
rect 633266 839006 633726 839068
rect 633266 837006 633726 837068
rect 633266 835904 633726 835974
rect 633266 835352 633726 835422
rect 633266 834708 633726 834778
rect 633266 834064 633726 834134
rect -400 827762 60 832542
rect 633266 832224 633726 832294
rect 633266 831672 633726 831742
rect 633266 831028 633726 831098
rect 633266 830384 633726 830454
rect 633266 827900 633726 827970
rect 633266 827348 633726 827418
rect 633266 826704 633726 826774
rect 633266 826060 633726 826130
rect 633266 825435 633726 825649
rect 633266 824864 633726 824934
rect 633266 823638 633726 823766
rect 633266 823024 633726 823094
rect 633266 821184 633726 821254
rect -400 795542 60 800322
rect -400 785562 60 790342
rect 633266 786384 633726 791164
rect 633266 776406 633726 781186
rect -400 757272 60 757342
rect -400 755432 60 755502
rect -400 754760 60 754888
rect -400 753592 60 753662
rect -400 752877 60 753091
rect -400 752396 60 752466
rect -400 751752 60 751822
rect -400 751108 60 751178
rect -400 750556 60 750626
rect 633266 750006 633726 750068
rect -400 748072 60 748142
rect 633266 748006 633726 748068
rect -400 747428 60 747498
rect -400 746784 60 746854
rect 633266 746704 633726 746774
rect -400 746232 60 746302
rect 633266 746152 633726 746222
rect 633266 745508 633726 745578
rect 633266 744864 633726 744934
rect -400 744392 60 744462
rect -400 743748 60 743818
rect -400 743104 60 743174
rect 633266 743024 633726 743094
rect -400 742552 60 742622
rect 633266 742472 633726 742542
rect 633266 741828 633726 741898
rect 633266 741184 633726 741254
rect 633266 738700 633726 738770
rect 633266 738148 633726 738218
rect 633266 737504 633726 737574
rect 633266 736860 633726 736930
rect -400 736644 60 736704
rect 633266 736235 633726 736449
rect 633266 735664 633726 735734
rect -400 734644 60 734704
rect 633266 734438 633726 734566
rect 633266 733824 633726 733894
rect 633266 731984 633726 732054
rect -400 714072 60 714142
rect -400 712232 60 712302
rect -400 711560 60 711688
rect -400 710392 60 710462
rect -400 709677 60 709891
rect -400 709196 60 709266
rect -400 708552 60 708622
rect -400 707908 60 707978
rect -400 707356 60 707426
rect 633266 705006 633726 705068
rect -400 704872 60 704942
rect -400 704228 60 704298
rect -400 703584 60 703654
rect -400 703032 60 703102
rect 633266 703006 633726 703068
rect 633266 701704 633726 701774
rect -400 701192 60 701262
rect 633266 701152 633726 701222
rect -400 700548 60 700618
rect 633266 700508 633726 700578
rect -400 699904 60 699974
rect 633266 699864 633726 699934
rect -400 699352 60 699422
rect 633266 698024 633726 698094
rect 633266 697472 633726 697542
rect 633266 696828 633726 696898
rect 633266 696184 633726 696254
rect -400 693644 60 693704
rect 633266 693700 633726 693770
rect 633266 693148 633726 693218
rect 633266 692504 633726 692574
rect 633266 691860 633726 691930
rect -400 691644 60 691704
rect 633266 691235 633726 691449
rect 633266 690664 633726 690734
rect 633266 689438 633726 689566
rect 633266 688824 633726 688894
rect 633266 686984 633726 687054
rect -400 670872 60 670942
rect -400 669032 60 669102
rect -400 668360 60 668488
rect -400 667192 60 667262
rect -400 666477 60 666691
rect -400 665996 60 666066
rect -400 665352 60 665422
rect -400 664708 60 664778
rect -400 664156 60 664226
rect -400 661672 60 661742
rect -400 661028 60 661098
rect -400 660384 60 660454
rect 633266 660006 633726 660068
rect -400 659832 60 659902
rect -400 657992 60 658062
rect 633266 658006 633726 658068
rect -400 657348 60 657418
rect -400 656704 60 656774
rect 633266 656704 633726 656774
rect -400 656152 60 656222
rect 633266 656152 633726 656222
rect 633266 655508 633726 655578
rect 633266 654864 633726 654934
rect 633266 653024 633726 653094
rect 633266 652472 633726 652542
rect 633266 651828 633726 651898
rect 633266 651184 633726 651254
rect -400 650644 60 650704
rect -400 648644 60 648704
rect 633266 648700 633726 648770
rect 633266 648148 633726 648218
rect 633266 647504 633726 647574
rect 633266 646860 633726 646930
rect 633266 646235 633726 646449
rect 633266 645664 633726 645734
rect 633266 644438 633726 644566
rect 633266 643824 633726 643894
rect 633266 641984 633726 642054
rect -400 627672 60 627742
rect -400 625832 60 625902
rect -400 625160 60 625288
rect -400 623992 60 624062
rect -400 623277 60 623491
rect -400 622796 60 622866
rect -400 622152 60 622222
rect -400 621508 60 621578
rect -400 620956 60 621026
rect -400 618472 60 618542
rect -400 617828 60 617898
rect -400 617184 60 617254
rect -400 616632 60 616702
rect 633266 615006 633726 615068
rect -400 614792 60 614862
rect -400 614148 60 614218
rect -400 613504 60 613574
rect -400 612952 60 613022
rect 633266 613006 633726 613068
rect 633266 611504 633726 611574
rect 633266 610952 633726 611022
rect 633266 610308 633726 610378
rect 633266 609664 633726 609734
rect 633266 607824 633726 607894
rect -400 607644 60 607704
rect 633266 607272 633726 607342
rect 633266 606628 633726 606698
rect 633266 605984 633726 606054
rect -400 605644 60 605704
rect 633266 603500 633726 603570
rect 633266 602948 633726 603018
rect 633266 602304 633726 602374
rect 633266 601660 633726 601730
rect 633266 601035 633726 601249
rect 633266 600464 633726 600534
rect 633266 599238 633726 599366
rect 633266 598624 633726 598694
rect 633266 596784 633726 596854
rect -400 584472 60 584542
rect -400 582632 60 582702
rect -400 581960 60 582088
rect -400 580792 60 580862
rect -400 580077 60 580291
rect -400 579596 60 579666
rect -400 578952 60 579022
rect -400 578308 60 578378
rect -400 577756 60 577826
rect -400 575272 60 575342
rect -400 574628 60 574698
rect -400 573984 60 574054
rect -400 573432 60 573502
rect -400 571592 60 571662
rect -400 570948 60 571018
rect -400 570304 60 570374
rect 633266 570006 633726 570068
rect -400 569752 60 569822
rect 633266 568006 633726 568068
rect 633266 566504 633726 566574
rect 633266 565952 633726 566022
rect 633266 565308 633726 565378
rect -400 564644 60 564704
rect 633266 564664 633726 564734
rect 633266 562824 633726 562894
rect -400 562644 60 562704
rect 633266 562272 633726 562342
rect 633266 561628 633726 561698
rect 633266 560984 633726 561054
rect 633266 558500 633726 558570
rect 633266 557948 633726 558018
rect 633266 557304 633726 557374
rect 633266 556660 633726 556730
rect 633266 556035 633726 556249
rect 633266 555464 633726 555534
rect 633266 554238 633726 554366
rect 633266 553624 633726 553694
rect 633266 551784 633726 551854
rect -400 541272 60 541342
rect -400 539432 60 539502
rect -400 538760 60 538888
rect -400 537592 60 537662
rect -400 536877 60 537091
rect -400 536396 60 536466
rect -400 535752 60 535822
rect -400 535108 60 535178
rect -400 534556 60 534626
rect -400 532072 60 532142
rect -400 531428 60 531498
rect -400 530784 60 530854
rect -400 530232 60 530302
rect -400 528392 60 528462
rect -400 527748 60 527818
rect -400 527104 60 527174
rect -400 526552 60 526622
rect 633266 525006 633726 525068
rect 633266 523005 633726 523067
rect -400 521644 60 521704
rect 633266 521304 633726 521374
rect 633266 520752 633726 520822
rect 633266 520108 633726 520178
rect -400 519644 60 519704
rect 633266 519464 633726 519534
rect 633266 517624 633726 517694
rect 633266 517072 633726 517142
rect 633266 516428 633726 516498
rect 633266 515784 633726 515854
rect 633266 513300 633726 513370
rect 633266 512748 633726 512818
rect 633266 512104 633726 512174
rect 633266 511460 633726 511530
rect 633266 510835 633726 511049
rect 633266 510264 633726 510334
rect 633266 509038 633726 509166
rect 633266 508424 633726 508494
rect 633266 506584 633726 506654
rect -400 498072 60 498142
rect -400 496232 60 496302
rect -400 495560 60 495688
rect -400 494392 60 494462
rect -400 493677 60 493891
rect -400 493196 60 493266
rect -400 492552 60 492622
rect -400 491908 60 491978
rect -400 491356 60 491426
rect -400 488872 60 488942
rect -400 488228 60 488298
rect -400 487584 60 487654
rect -400 487032 60 487102
rect -400 485192 60 485262
rect -400 484548 60 484618
rect -400 483904 60 483974
rect -400 483352 60 483422
rect -400 478644 60 478704
rect -400 476644 60 476704
rect 633266 471784 633726 476564
rect 633266 461804 633726 466584
rect -400 450940 60 455720
rect -400 440962 60 445742
rect 633266 427762 633726 432562
rect 633266 422810 633726 427472
rect 633266 417722 633726 422512
rect -400 408814 60 413604
rect -400 403862 60 408514
rect -400 398762 60 403562
rect 633266 383584 633726 388364
rect 633266 373606 633726 378386
rect -400 370472 60 370542
rect -400 368632 60 368702
rect -400 367960 60 368088
rect -400 366792 60 366862
rect -400 366077 60 366291
rect -400 365596 60 365666
rect -400 364952 60 365022
rect -400 364308 60 364378
rect -400 363756 60 363826
rect -400 361272 60 361342
rect -400 360628 60 360698
rect -400 359984 60 360054
rect -400 359432 60 359502
rect -400 357592 60 357662
rect -400 356948 60 357018
rect -400 356304 60 356374
rect -400 355752 60 355822
rect -400 349644 60 349704
rect 633266 348006 633726 348068
rect -400 347644 60 347704
rect 633266 346005 633726 346067
rect 633266 344104 633726 344174
rect 633266 343552 633726 343622
rect 633266 342908 633726 342978
rect 633266 342264 633726 342334
rect 633266 340424 633726 340494
rect 633266 339872 633726 339942
rect 633266 339228 633726 339298
rect 633266 338584 633726 338654
rect 633266 336100 633726 336170
rect 633266 335548 633726 335618
rect 633266 334904 633726 334974
rect 633266 334260 633726 334330
rect 633266 333635 633726 333849
rect 633266 333064 633726 333134
rect 633266 331838 633726 331966
rect 633266 331224 633726 331294
rect 633266 329384 633726 329454
rect -400 327272 60 327342
rect -400 325432 60 325502
rect -400 324760 60 324888
rect -400 323592 60 323662
rect -400 322877 60 323091
rect -400 322396 60 322466
rect -400 321752 60 321822
rect -400 321108 60 321178
rect -400 320556 60 320626
rect -400 318072 60 318142
rect -400 317428 60 317498
rect -400 316784 60 316854
rect -400 316232 60 316302
rect -400 314392 60 314462
rect -400 313748 60 313818
rect -400 313104 60 313174
rect -400 312552 60 312622
rect -400 306644 60 306704
rect -400 304644 60 304704
rect 633266 303006 633726 303068
rect 633266 301005 633726 301067
rect 633266 298904 633726 298974
rect 633266 298352 633726 298422
rect 633266 297708 633726 297778
rect 633266 297064 633726 297134
rect 633266 295224 633726 295294
rect 633266 294672 633726 294742
rect 633266 294028 633726 294098
rect 633266 293384 633726 293454
rect 633266 290900 633726 290970
rect 633266 290348 633726 290418
rect 633266 289704 633726 289774
rect 633266 289060 633726 289130
rect 633266 288435 633726 288649
rect 633266 287864 633726 287934
rect 633266 286638 633726 286766
rect 633266 286024 633726 286094
rect 633266 284184 633726 284254
rect -400 284072 60 284142
rect -400 282232 60 282302
rect -400 281560 60 281688
rect -400 280392 60 280462
rect -400 279677 60 279891
rect -400 279196 60 279266
rect -400 278552 60 278622
rect -400 277908 60 277978
rect -400 277356 60 277426
rect -400 274872 60 274942
rect -400 274228 60 274298
rect -400 273584 60 273654
rect -400 273032 60 273102
rect -400 271192 60 271262
rect -400 270548 60 270618
rect -400 269904 60 269974
rect -400 269352 60 269422
rect -400 263644 60 263704
rect -400 261644 60 261704
rect 633266 258006 633726 258068
rect 633266 256005 633726 256067
rect 633266 253904 633726 253974
rect 633266 253352 633726 253422
rect 633266 252708 633726 252778
rect 633266 252064 633726 252134
rect 633266 250224 633726 250294
rect 633266 249672 633726 249742
rect 633266 249028 633726 249098
rect 633266 248384 633726 248454
rect 633266 245900 633726 245970
rect 633266 245348 633726 245418
rect 633266 244704 633726 244774
rect 633266 244060 633726 244130
rect 633266 243435 633726 243649
rect 633266 242864 633726 242934
rect 633266 241638 633726 241766
rect 633266 241024 633726 241094
rect -400 240872 60 240942
rect 633266 239184 633726 239254
rect -400 239032 60 239102
rect -400 238360 60 238488
rect -400 237192 60 237262
rect -400 236477 60 236691
rect -400 235996 60 236066
rect -400 235352 60 235422
rect -400 234708 60 234778
rect -400 234156 60 234226
rect -400 231672 60 231742
rect -400 231028 60 231098
rect -400 230384 60 230454
rect -400 229832 60 229902
rect -400 227992 60 228062
rect -400 227348 60 227418
rect -400 226704 60 226774
rect -400 226152 60 226222
rect -400 220644 60 220704
rect -400 218644 60 218704
rect 633266 213006 633726 213068
rect 633266 211005 633726 211067
rect 633266 208904 633726 208974
rect 633266 208352 633726 208422
rect 633266 207708 633726 207778
rect 633266 207064 633726 207134
rect 633266 205224 633726 205294
rect 633266 204672 633726 204742
rect 633266 204028 633726 204098
rect 633266 203384 633726 203454
rect 633266 200900 633726 200970
rect 633266 200348 633726 200418
rect 633266 199704 633726 199774
rect 633266 199060 633726 199130
rect 633266 198435 633726 198649
rect 633266 197864 633726 197934
rect -400 197672 60 197742
rect 633266 196638 633726 196766
rect 633266 196024 633726 196094
rect -400 195832 60 195902
rect -400 195160 60 195288
rect 633266 194184 633726 194254
rect -400 193992 60 194062
rect -400 193277 60 193491
rect -400 192796 60 192866
rect -400 192152 60 192222
rect -400 191508 60 191578
rect -400 190956 60 191026
rect -400 188472 60 188542
rect -400 187828 60 187898
rect -400 187184 60 187254
rect -400 186632 60 186702
rect -400 184792 60 184862
rect -400 184148 60 184218
rect -400 183504 60 183574
rect -400 182952 60 183022
rect -400 177644 60 177704
rect -400 175644 60 175704
rect 633266 168006 633726 168068
rect 633266 166005 633726 166067
rect 633266 163704 633726 163774
rect 633266 163152 633726 163222
rect 633266 162508 633726 162578
rect 633266 161864 633726 161934
rect 633266 160024 633726 160094
rect 633266 159472 633726 159542
rect 633266 158828 633726 158898
rect 633266 158184 633726 158254
rect 633266 155700 633726 155770
rect 633266 155148 633726 155218
rect -400 154472 60 154542
rect 633266 154504 633726 154574
rect 633266 153860 633726 153930
rect 633266 153235 633726 153449
rect -400 152632 60 152702
rect 633266 152664 633726 152734
rect -400 151960 60 152088
rect 633266 151438 633726 151566
rect -400 150792 60 150862
rect 633266 150824 633726 150894
rect -400 150077 60 150291
rect -400 149596 60 149666
rect -400 148952 60 149022
rect 633266 148984 633726 149054
rect -400 148308 60 148378
rect -400 147756 60 147826
rect -400 145272 60 145342
rect -400 144628 60 144698
rect -400 143984 60 144054
rect -400 143432 60 143502
rect -400 141592 60 141662
rect -400 140948 60 141018
rect -400 140304 60 140374
rect -400 139752 60 139822
rect -400 134644 60 134704
rect -400 132644 60 132704
rect 633266 123006 633726 123068
rect 633266 121005 633726 121067
rect 633266 118704 633726 118774
rect 633266 118152 633726 118222
rect 633266 117508 633726 117578
rect 633266 116864 633726 116934
rect 633266 115024 633726 115094
rect 633266 114472 633726 114542
rect 633266 113828 633726 113898
rect 633266 113184 633726 113254
rect 633266 110700 633726 110770
rect 633266 110148 633726 110218
rect 633266 109504 633726 109574
rect 633266 108860 633726 108930
rect 633266 108235 633726 108449
rect 633266 107664 633726 107734
rect 633266 106438 633726 106566
rect 633266 105824 633726 105894
rect 633266 103984 633726 104054
rect -400 78140 60 82920
rect 633266 78006 633726 78068
rect 633266 76005 633726 76067
rect 633266 73504 633726 73574
rect 633266 72952 633726 73022
rect -400 68162 60 72942
rect 633266 72308 633726 72378
rect 633266 71664 633726 71734
rect 633266 69824 633726 69894
rect 633266 69272 633726 69342
rect 633266 68628 633726 68698
rect 633266 67984 633726 68054
rect 633266 65500 633726 65570
rect 633266 64948 633726 65018
rect 633266 64304 633726 64374
rect 633266 63660 633726 63730
rect 633266 63035 633726 63249
rect 633266 62464 633726 62534
rect 633266 61238 633726 61366
rect 633266 60624 633726 60694
rect 633266 58784 633726 58854
rect -400 53595 60 53665
rect -400 53372 60 53442
rect -400 53147 60 53217
rect -400 36014 60 40804
rect -400 25962 60 30762
rect 36806 -400 41586 60
rect 46784 -400 51564 60
rect 199284 -400 203914 60
rect 209164 -400 213964 60
rect 527006 -400 531786 60
rect 536984 -400 541764 60
rect 580806 -400 585586 60
rect 590784 -400 595564 60
<< comment >>
rect -400 953326 633726 953726
rect -400 0 0 953326
rect 633326 58370 633726 953326
rect 633326 0 633726 58369
rect -400 -400 633726 0
<< labels >>
flabel metal2 485870 -400 485926 56 0 FreeSans 400 270 0 0 gpio_vtrip_sel[43]
port 290 nsew
flabel metal2 s 594004 953270 594060 953726 0 FreeSans 400 90 0 0 gpio_analog_en[15]
port 450 nsew
flabel metal2 s 592716 953270 592772 953726 0 FreeSans 400 90 0 0 gpio_analog_pol[15]
port 538 nsew
flabel metal2 s 589680 953270 589736 953726 0 FreeSans 400 90 0 0 gpio_analog_sel[15]
port 494 nsew
flabel metal2 s 593360 953270 593416 953726 0 FreeSans 400 90 0 0 gpio_dm0[15]
port 582 nsew
flabel metal2 s 595200 953270 595256 953726 0 FreeSans 400 90 0 0 gpio_dm1[15]
port 626 nsew
flabel metal2 s 589036 953270 589092 953726 0 FreeSans 400 90 0 0 gpio_dm2[15]
port 670 nsew
flabel metal2 s 588392 953270 588448 953726 0 FreeSans 400 90 0 0 gpio_holdover[15]
port 406 nsew
flabel metal2 s 585356 953270 585412 953726 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[15]
port 274 nsew
flabel metal2 s 592164 953270 592220 953726 0 FreeSans 400 90 0 0 gpio_inp_dis[15]
port 230 nsew
flabel metal2 s 584712 953270 584768 953726 0 FreeSans 400 90 0 0 gpio_oeb[15]
port 186 nsew
flabel metal2 s 587840 953270 587896 953726 0 FreeSans 400 90 0 0 gpio_out[15]
port 142 nsew
flabel metal2 s 597040 953270 597096 953726 0 FreeSans 400 90 0 0 gpio_slow_sel[15]
port 362 nsew
flabel metal2 s 586000 953270 586056 953726 0 FreeSans 400 90 0 0 gpio_vtrip_sel[15]
port 318 nsew
flabel metal2 s 598880 953270 598936 953726 0 FreeSans 400 90 0 0 gpio_in[15]
port 714 nsew
flabel metal2 s 492204 953270 492260 953726 0 FreeSans 400 90 0 0 gpio_analog_en[16]
port 449 nsew
flabel metal2 s 490916 953270 490972 953726 0 FreeSans 400 90 0 0 gpio_analog_pol[16]
port 537 nsew
flabel metal2 s 487880 953270 487936 953726 0 FreeSans 400 90 0 0 gpio_analog_sel[16]
port 493 nsew
flabel metal2 s 491560 953270 491616 953726 0 FreeSans 400 90 0 0 gpio_dm0[16]
port 581 nsew
flabel metal2 s 493400 953270 493456 953726 0 FreeSans 400 90 0 0 gpio_dm1[16]
port 625 nsew
flabel metal2 s 487236 953270 487292 953726 0 FreeSans 400 90 0 0 gpio_dm2[16]
port 669 nsew
flabel metal2 s 486592 953270 486648 953726 0 FreeSans 400 90 0 0 gpio_holdover[16]
port 405 nsew
flabel metal2 s 483556 953270 483612 953726 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[16]
port 273 nsew
flabel metal2 s 490364 953270 490420 953726 0 FreeSans 400 90 0 0 gpio_inp_dis[16]
port 229 nsew
flabel metal2 s 482912 953270 482968 953726 0 FreeSans 400 90 0 0 gpio_oeb[16]
port 185 nsew
flabel metal2 s 486040 953270 486096 953726 0 FreeSans 400 90 0 0 gpio_out[16]
port 141 nsew
flabel metal2 s 495240 953270 495296 953726 0 FreeSans 400 90 0 0 gpio_slow_sel[16]
port 361 nsew
flabel metal2 s 484200 953270 484256 953726 0 FreeSans 400 90 0 0 gpio_vtrip_sel[16]
port 317 nsew
flabel metal2 s 497080 953270 497136 953726 0 FreeSans 400 90 0 0 gpio_in[16]
port 713 nsew
flabel metal2 s 442000 953270 442056 953726 0 FreeSans 400 90 0 0 gpio_dm1[17]
port 624 nsew
flabel metal2 s 435836 953270 435892 953726 0 FreeSans 400 90 0 0 gpio_dm2[17]
port 668 nsew
flabel metal2 s 435192 953270 435248 953726 0 FreeSans 400 90 0 0 gpio_holdover[17]
port 404 nsew
flabel metal2 s 432156 953270 432212 953726 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[17]
port 272 nsew
flabel metal2 s 438964 953270 439020 953726 0 FreeSans 400 90 0 0 gpio_inp_dis[17]
port 228 nsew
flabel metal2 s 431512 953270 431568 953726 0 FreeSans 400 90 0 0 gpio_oeb[17]
port 184 nsew
flabel metal2 s 434640 953270 434696 953726 0 FreeSans 400 90 0 0 gpio_out[17]
port 140 nsew
flabel metal2 s 443840 953270 443896 953726 0 FreeSans 400 90 0 0 gpio_slow_sel[17]
port 360 nsew
flabel metal2 s 432800 953270 432856 953726 0 FreeSans 400 90 0 0 gpio_vtrip_sel[17]
port 316 nsew
flabel metal2 s 445680 953270 445736 953726 0 FreeSans 400 90 0 0 gpio_in[17]
port 712 nsew
flabel metal2 s 351804 953270 351860 953726 0 FreeSans 400 90 0 0 gpio_analog_en[18]
port 447 nsew
flabel metal2 s 350516 953270 350572 953726 0 FreeSans 400 90 0 0 gpio_analog_pol[18]
port 535 nsew
flabel metal2 s 347480 953270 347536 953726 0 FreeSans 400 90 0 0 gpio_analog_sel[18]
port 491 nsew
flabel metal2 s 351160 953270 351216 953726 0 FreeSans 400 90 0 0 gpio_dm0[18]
port 579 nsew
flabel metal2 s 353000 953270 353056 953726 0 FreeSans 400 90 0 0 gpio_dm1[18]
port 623 nsew
flabel metal2 s 346836 953270 346892 953726 0 FreeSans 400 90 0 0 gpio_dm2[18]
port 667 nsew
flabel metal2 s 346192 953270 346248 953726 0 FreeSans 400 90 0 0 gpio_holdover[18]
port 403 nsew
flabel metal2 s 343156 953270 343212 953726 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[18]
port 271 nsew
flabel metal2 s 349964 953270 350020 953726 0 FreeSans 400 90 0 0 gpio_inp_dis[18]
port 227 nsew
flabel metal2 s 342512 953270 342568 953726 0 FreeSans 400 90 0 0 gpio_oeb[18]
port 183 nsew
flabel metal2 s 345640 953270 345696 953726 0 FreeSans 400 90 0 0 gpio_out[18]
port 139 nsew
flabel metal2 s 354840 953270 354896 953726 0 FreeSans 400 90 0 0 gpio_slow_sel[18]
port 359 nsew
flabel metal2 s 343800 953270 343856 953726 0 FreeSans 400 90 0 0 gpio_vtrip_sel[18]
port 315 nsew
flabel metal2 s 356680 953270 356736 953726 0 FreeSans 400 90 0 0 gpio_in[18]
port 711 nsew
flabel metal2 s 440804 953270 440860 953726 0 FreeSans 400 90 0 0 gpio_analog_en[17]
port 448 nsew
flabel metal2 s 439516 953270 439572 953726 0 FreeSans 400 90 0 0 gpio_analog_pol[17]
port 536 nsew
flabel metal2 s 436480 953270 436536 953726 0 FreeSans 400 90 0 0 gpio_analog_sel[17]
port 492 nsew
flabel metal2 s 440160 953270 440216 953726 0 FreeSans 400 90 0 0 gpio_dm0[17]
port 580 nsew
flabel metal2 s 253040 953270 253096 953726 0 FreeSans 400 90 0 0 gpio_slow_sel[19]
port 358 nsew
flabel metal2 s 242000 953270 242056 953726 0 FreeSans 400 90 0 0 gpio_vtrip_sel[19]
port 314 nsew
flabel metal2 s 254880 953270 254936 953726 0 FreeSans 400 90 0 0 gpio_in[19]
port 710 nsew
flabel metal2 s 198404 953270 198460 953726 0 FreeSans 400 90 0 0 gpio_analog_en[20]
port 445 nsew
flabel metal2 s 197116 953270 197172 953726 0 FreeSans 400 90 0 0 gpio_analog_pol[20]
port 533 nsew
flabel metal2 s 194080 953270 194136 953726 0 FreeSans 400 90 0 0 gpio_analog_sel[20]
port 489 nsew
flabel metal2 s 197760 953270 197816 953726 0 FreeSans 400 90 0 0 gpio_dm0[20]
port 577 nsew
flabel metal2 s 199600 953270 199656 953726 0 FreeSans 400 90 0 0 gpio_dm1[20]
port 621 nsew
flabel metal2 s 193436 953270 193492 953726 0 FreeSans 400 90 0 0 gpio_dm2[20]
port 665 nsew
flabel metal2 s 192792 953270 192848 953726 0 FreeSans 400 90 0 0 gpio_holdover[20]
port 401 nsew
flabel metal2 s 189756 953270 189812 953726 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[20]
port 269 nsew
flabel metal2 s 196564 953270 196620 953726 0 FreeSans 400 90 0 0 gpio_inp_dis[20]
port 225 nsew
flabel metal2 s 189112 953270 189168 953726 0 FreeSans 400 90 0 0 gpio_oeb[20]
port 181 nsew
flabel metal2 s 192240 953270 192296 953726 0 FreeSans 400 90 0 0 gpio_out[20]
port 137 nsew
flabel metal2 s 201440 953270 201496 953726 0 FreeSans 400 90 0 0 gpio_slow_sel[20]
port 357 nsew
flabel metal2 s 190400 953270 190456 953726 0 FreeSans 400 90 0 0 gpio_vtrip_sel[20]
port 313 nsew
flabel metal2 s 203280 953270 203336 953726 0 FreeSans 400 90 0 0 gpio_in[20]
port 709 nsew
flabel metal2 s 250004 953270 250060 953726 0 FreeSans 400 90 0 0 gpio_analog_en[19]
port 446 nsew
flabel metal2 s 248716 953270 248772 953726 0 FreeSans 400 90 0 0 gpio_analog_pol[19]
port 534 nsew
flabel metal2 s 245680 953270 245736 953726 0 FreeSans 400 90 0 0 gpio_analog_sel[19]
port 490 nsew
flabel metal2 s 249360 953270 249416 953726 0 FreeSans 400 90 0 0 gpio_dm0[19]
port 578 nsew
flabel metal2 s 251200 953270 251256 953726 0 FreeSans 400 90 0 0 gpio_dm1[19]
port 622 nsew
flabel metal2 s 245036 953270 245092 953726 0 FreeSans 400 90 0 0 gpio_dm2[19]
port 666 nsew
flabel metal2 s 244392 953270 244448 953726 0 FreeSans 400 90 0 0 gpio_holdover[19]
port 402 nsew
flabel metal2 s 241356 953270 241412 953726 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[19]
port 270 nsew
flabel metal2 s 248164 953270 248220 953726 0 FreeSans 400 90 0 0 gpio_inp_dis[19]
port 226 nsew
flabel metal2 s 240712 953270 240768 953726 0 FreeSans 400 90 0 0 gpio_oeb[19]
port 182 nsew
flabel metal2 s 243840 953270 243896 953726 0 FreeSans 400 90 0 0 gpio_out[19]
port 138 nsew
flabel metal2 s 151880 953270 151936 953726 0 FreeSans 400 90 0 0 gpio_in[21]
port 708 nsew
flabel metal2 s 95604 953270 95660 953726 0 FreeSans 400 90 0 0 gpio_analog_en[22]
port 443 nsew
flabel metal2 s 94316 953270 94372 953726 0 FreeSans 400 90 0 0 gpio_analog_pol[22]
port 531 nsew
flabel metal2 s 91280 953270 91336 953726 0 FreeSans 400 90 0 0 gpio_analog_sel[22]
port 487 nsew
flabel metal2 s 94960 953270 95016 953726 0 FreeSans 400 90 0 0 gpio_dm0[22]
port 575 nsew
flabel metal2 s 96800 953270 96856 953726 0 FreeSans 400 90 0 0 gpio_dm1[22]
port 619 nsew
flabel metal2 s 90636 953270 90692 953726 0 FreeSans 400 90 0 0 gpio_dm2[22]
port 663 nsew
flabel metal2 s 89992 953270 90048 953726 0 FreeSans 400 90 0 0 gpio_holdover[22]
port 399 nsew
flabel metal2 s 86956 953270 87012 953726 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[22]
port 267 nsew
flabel metal2 s 93764 953270 93820 953726 0 FreeSans 400 90 0 0 gpio_inp_dis[22]
port 223 nsew
flabel metal2 s 86312 953270 86368 953726 0 FreeSans 400 90 0 0 gpio_oeb[22]
port 179 nsew
flabel metal2 s 89440 953270 89496 953726 0 FreeSans 400 90 0 0 gpio_out[22]
port 135 nsew
flabel metal2 s 98640 953270 98696 953726 0 FreeSans 400 90 0 0 gpio_slow_sel[22]
port 355 nsew
flabel metal2 s 87600 953270 87656 953726 0 FreeSans 400 90 0 0 gpio_vtrip_sel[22]
port 311 nsew
flabel metal2 s 100480 953270 100536 953726 0 FreeSans 400 90 0 0 gpio_in[22]
port 707 nsew
flabel metal2 s 44204 953270 44260 953726 0 FreeSans 400 90 0 0 gpio_analog_en[23]
port 442 nsew
flabel metal2 s 42916 953270 42972 953726 0 FreeSans 400 90 0 0 gpio_analog_pol[23]
port 530 nsew
flabel metal2 s 39880 953270 39936 953726 0 FreeSans 400 90 0 0 gpio_analog_sel[23]
port 486 nsew
flabel metal2 s 43560 953270 43616 953726 0 FreeSans 400 90 0 0 gpio_dm0[23]
port 574 nsew
flabel metal2 s 45400 953270 45456 953726 0 FreeSans 400 90 0 0 gpio_dm1[23]
port 618 nsew
flabel metal2 s 39236 953270 39292 953726 0 FreeSans 400 90 0 0 gpio_dm2[23]
port 662 nsew
flabel metal2 s 38592 953270 38648 953726 0 FreeSans 400 90 0 0 gpio_holdover[23]
port 398 nsew
flabel metal2 s 35556 953270 35612 953726 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[23]
port 266 nsew
flabel metal2 s 42364 953270 42420 953726 0 FreeSans 400 90 0 0 gpio_inp_dis[23]
port 222 nsew
flabel metal2 s 34912 953270 34968 953726 0 FreeSans 400 90 0 0 gpio_oeb[23]
port 178 nsew
flabel metal2 s 38040 953270 38096 953726 0 FreeSans 400 90 0 0 gpio_out[23]
port 134 nsew
flabel metal2 s 47240 953270 47296 953726 0 FreeSans 400 90 0 0 gpio_slow_sel[23]
port 354 nsew
flabel metal2 s 36200 953270 36256 953726 0 FreeSans 400 90 0 0 gpio_vtrip_sel[23]
port 310 nsew
flabel metal2 s 49080 953270 49136 953726 0 FreeSans 400 90 0 0 gpio_in[23]
port 706 nsew
flabel metal2 s 147004 953270 147060 953726 0 FreeSans 400 90 0 0 gpio_analog_en[21]
port 444 nsew
flabel metal2 s 145716 953270 145772 953726 0 FreeSans 400 90 0 0 gpio_analog_pol[21]
port 532 nsew
flabel metal2 s 142680 953270 142736 953726 0 FreeSans 400 90 0 0 gpio_analog_sel[21]
port 488 nsew
flabel metal2 s 146360 953270 146416 953726 0 FreeSans 400 90 0 0 gpio_dm0[21]
port 576 nsew
flabel metal2 s 148200 953270 148256 953726 0 FreeSans 400 90 0 0 gpio_dm1[21]
port 620 nsew
flabel metal2 s 142036 953270 142092 953726 0 FreeSans 400 90 0 0 gpio_dm2[21]
port 664 nsew
flabel metal2 s 141392 953270 141448 953726 0 FreeSans 400 90 0 0 gpio_holdover[21]
port 400 nsew
flabel metal2 s 138356 953270 138412 953726 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[21]
port 268 nsew
flabel metal2 s 145164 953270 145220 953726 0 FreeSans 400 90 0 0 gpio_inp_dis[21]
port 224 nsew
flabel metal2 s 137712 953270 137768 953726 0 FreeSans 400 90 0 0 gpio_oeb[21]
port 180 nsew
flabel metal2 s 140840 953270 140896 953726 0 FreeSans 400 90 0 0 gpio_out[21]
port 136 nsew
flabel metal2 s 150040 953270 150096 953726 0 FreeSans 400 90 0 0 gpio_slow_sel[21]
port 356 nsew
flabel metal2 s 139000 953270 139056 953726 0 FreeSans 400 90 0 0 gpio_vtrip_sel[21]
port 312 nsew
flabel metal2 145190 -400 145246 56 0 FreeSans 400 270 0 0 gpio_in[38]
port 691 nsew
flabel metal2 147030 -400 147086 56 0 FreeSans 400 270 0 0 gpio_slow_sel[38]
port 339 nsew
flabel metal2 148870 -400 148926 56 0 FreeSans 400 270 0 0 gpio_dm1[38]
port 559 nsew
flabel metal2 150710 -400 150766 56 0 FreeSans 400 270 0 0 gpio_dm0[38]
port 603 nsew
flabel metal2 151354 -400 151410 56 0 FreeSans 400 270 0 0 gpio_analog_pol[38]
port 515 nsew
flabel metal2 150066 -400 150122 56 0 FreeSans 400 270 0 0 gpio_analog_en[38]
port 427 nsew
flabel metal2 151906 -400 151962 56 0 FreeSans 400 270 0 0 gpio_inp_dis[38]
port 207 nsew
flabel metal2 154390 -400 154446 56 0 FreeSans 400 270 0 0 gpio_analog_sel[38]
port 471 nsew
flabel metal2 155034 -400 155090 56 0 FreeSans 400 270 0 0 gpio_dm2[38]
port 647 nsew
flabel metal2 155678 -400 155734 56 0 FreeSans 400 270 0 0 gpio_holdover[38]
port 383 nsew
flabel metal2 156230 -400 156286 56 0 FreeSans 400 270 0 0 gpio_out[38]
port 119 nsew
flabel metal2 158070 -400 158126 56 0 FreeSans 400 270 0 0 gpio_vtrip_sel[38]
port 295 nsew
flabel metal2 158714 -400 158770 56 0 FreeSans 400 270 0 0 gpio_ib_mode_sel[38]
port 251 nsew
flabel metal2 159358 -400 159414 56 0 FreeSans 400 270 0 0 gpio_oeb[38]
port 163 nsew
flabel metal2 253790 -400 253846 56 0 FreeSans 400 270 0 0 gpio_in[39]
port 690 nsew
flabel metal2 255630 -400 255686 56 0 FreeSans 400 270 0 0 gpio_slow_sel[39]
port 338 nsew
flabel metal2 257470 -400 257526 56 0 FreeSans 400 270 0 0 gpio_dm1[39]
port 602 nsew
flabel metal2 259310 -400 259366 56 0 FreeSans 400 270 0 0 gpio_dm0[39]
port 558 nsew
flabel metal2 259954 -400 260010 56 0 FreeSans 400 270 0 0 gpio_analog_pol[39]
port 514 nsew
flabel metal2 258666 -400 258722 56 0 FreeSans 400 270 0 0 gpio_analog_en[39]
port 426 nsew
flabel metal2 260506 -400 260562 56 0 FreeSans 400 270 0 0 gpio_inp_dis[39]
port 206 nsew
flabel metal2 262990 -400 263046 56 0 FreeSans 400 270 0 0 gpio_analog_sel[39]
port 470 nsew
flabel metal2 263634 -400 263690 56 0 FreeSans 400 270 0 0 gpio_dm2[39]
port 646 nsew
flabel metal2 264278 -400 264334 56 0 FreeSans 400 270 0 0 gpio_holdover[39]
port 382 nsew
flabel metal2 264830 -400 264886 56 0 FreeSans 400 270 0 0 gpio_out[39]
port 118 nsew
flabel metal2 266670 -400 266726 56 0 FreeSans 400 270 0 0 gpio_vtrip_sel[39]
port 294 nsew
flabel metal2 267314 -400 267370 56 0 FreeSans 400 270 0 0 gpio_ib_mode_sel[39]
port 250 nsew
flabel metal2 267958 -400 268014 56 0 FreeSans 400 270 0 0 gpio_oeb[39]
port 162 nsew
flabel metal2 308590 -400 308646 56 0 FreeSans 400 270 0 0 gpio_in[40]
port 689 nsew
flabel metal2 310430 -400 310486 56 0 FreeSans 400 270 0 0 gpio_slow_sel[40]
port 337 nsew
flabel metal2 312270 -400 312326 56 0 FreeSans 400 270 0 0 gpio_dm1[40]
port 601 nsew
flabel metal2 314110 -400 314166 56 0 FreeSans 400 270 0 0 gpio_dm0[40]
port 557 nsew
flabel metal2 314754 -400 314810 56 0 FreeSans 400 270 0 0 gpio_analog_pol[40]
port 513 nsew
flabel metal2 313466 -400 313522 56 0 FreeSans 400 270 0 0 gpio_analog_en[40]
port 425 nsew
flabel metal2 315306 -400 315362 56 0 FreeSans 400 270 0 0 gpio_inp_dis[40]
port 205 nsew
flabel metal2 317790 -400 317846 56 0 FreeSans 400 270 0 0 gpio_analog_sel[40]
port 469 nsew
flabel metal2 318434 -400 318490 56 0 FreeSans 400 270 0 0 gpio_dm2[40]
port 645 nsew
flabel metal2 319078 -400 319134 56 0 FreeSans 400 270 0 0 gpio_holdover[40]
port 381 nsew
flabel metal2 319630 -400 319686 56 0 FreeSans 400 270 0 0 gpio_out[40]
port 117 nsew
flabel metal2 321470 -400 321526 56 0 FreeSans 400 270 0 0 gpio_vtrip_sel[40]
port 293 nsew
flabel metal2 322114 -400 322170 56 0 FreeSans 400 270 0 0 gpio_ib_mode_sel[40]
port 249 nsew
flabel metal2 322758 -400 322814 56 0 FreeSans 400 270 0 0 gpio_oeb[40]
port 161 nsew
flabel metal2 363390 -400 363446 56 0 FreeSans 400 270 0 0 gpio_in[41]
port 688 nsew
flabel metal2 365230 -400 365286 56 0 FreeSans 400 270 0 0 gpio_slow_sel[41]
port 336 nsew
flabel metal2 367070 -400 367126 56 0 FreeSans 400 270 0 0 gpio_dm1[41]
port 600 nsew
flabel metal2 368910 -400 368966 56 0 FreeSans 400 270 0 0 gpio_dm0[41]
port 556 nsew
flabel metal2 369554 -400 369610 56 0 FreeSans 400 270 0 0 gpio_analog_pol[41]
port 512 nsew
flabel metal2 368266 -400 368322 56 0 FreeSans 400 270 0 0 gpio_analog_en[41]
port 424 nsew
flabel metal2 370106 -400 370162 56 0 FreeSans 400 270 0 0 gpio_inp_dis[41]
port 204 nsew
flabel metal2 372590 -400 372646 56 0 FreeSans 400 270 0 0 gpio_analog_sel[41]
port 468 nsew
flabel metal2 373234 -400 373290 56 0 FreeSans 400 270 0 0 gpio_dm2[41]
port 644 nsew
flabel metal2 373878 -400 373934 56 0 FreeSans 400 270 0 0 gpio_holdover[41]
port 380 nsew
flabel metal2 374430 -400 374486 56 0 FreeSans 400 270 0 0 gpio_out[41]
port 116 nsew
flabel metal2 376270 -400 376326 56 0 FreeSans 400 270 0 0 gpio_vtrip_sel[41]
port 292 nsew
flabel metal2 376914 -400 376970 56 0 FreeSans 400 270 0 0 gpio_ib_mode_sel[41]
port 248 nsew
flabel metal2 377558 -400 377614 56 0 FreeSans 400 270 0 0 gpio_oeb[41]
port 160 nsew
flabel metal2 418190 -400 418246 56 0 FreeSans 400 270 0 0 gpio_in[42]
port 687 nsew
flabel metal2 420030 -400 420086 56 0 FreeSans 400 270 0 0 gpio_slow_sel[42]
port 335 nsew
flabel metal2 421870 -400 421926 56 0 FreeSans 400 270 0 0 gpio_dm1[42]
port 599 nsew
flabel metal2 423710 -400 423766 56 0 FreeSans 400 270 0 0 gpio_dm0[42]
port 555 nsew
flabel metal2 424354 -400 424410 56 0 FreeSans 400 270 0 0 gpio_analog_pol[42]
port 511 nsew
flabel metal2 423066 -400 423122 56 0 FreeSans 400 270 0 0 gpio_analog_en[42]
port 423 nsew
flabel metal2 424906 -400 424962 56 0 FreeSans 400 270 0 0 gpio_inp_dis[42]
port 203 nsew
flabel metal2 427390 -400 427446 56 0 FreeSans 400 270 0 0 gpio_analog_sel[42]
port 467 nsew
flabel metal2 428034 -400 428090 56 0 FreeSans 400 270 0 0 gpio_dm2[42]
port 643 nsew
flabel metal2 428678 -400 428734 56 0 FreeSans 400 270 0 0 gpio_holdover[42]
port 379 nsew
flabel metal2 429230 -400 429286 56 0 FreeSans 400 270 0 0 gpio_out[42]
port 115 nsew
flabel metal2 431070 -400 431126 56 0 FreeSans 400 270 0 0 gpio_vtrip_sel[42]
port 291 nsew
flabel metal2 431714 -400 431770 56 0 FreeSans 400 270 0 0 gpio_ib_mode_sel[42]
port 247 nsew
flabel metal2 432358 -400 432414 56 0 FreeSans 400 270 0 0 gpio_oeb[42]
port 159 nsew
flabel metal2 472990 -400 473046 56 0 FreeSans 400 270 0 0 gpio_in[43]
port 686 nsew
flabel metal2 474830 -400 474886 56 0 FreeSans 400 270 0 0 gpio_slow_sel[43]
port 334 nsew
flabel metal2 476670 -400 476726 56 0 FreeSans 400 270 0 0 gpio_dm1[43]
port 598 nsew
flabel metal2 478510 -400 478566 56 0 FreeSans 400 270 0 0 gpio_dm0[43]
port 554 nsew
flabel metal2 479154 -400 479210 56 0 FreeSans 400 270 0 0 gpio_analog_pol[43]
port 510 nsew
flabel metal2 477866 -400 477922 56 0 FreeSans 400 270 0 0 gpio_analog_en[43]
port 422 nsew
flabel metal2 479706 -400 479762 56 0 FreeSans 400 270 0 0 gpio_inp_dis[43]
port 202 nsew
flabel metal2 482190 -400 482246 56 0 FreeSans 400 270 0 0 gpio_analog_sel[43]
port 466 nsew
flabel metal2 482834 -400 482890 56 0 FreeSans 400 270 0 0 gpio_dm2[43]
port 642 nsew
flabel metal2 483478 -400 483534 56 0 FreeSans 400 270 0 0 gpio_holdover[43]
port 378 nsew
flabel metal2 484030 -400 484086 56 0 FreeSans 400 270 0 0 gpio_out[43]
port 114 nsew
flabel metal2 486514 -400 486570 56 0 FreeSans 400 270 0 0 gpio_ib_mode_sel[43]
port 246 nsew
flabel metal2 487158 -400 487214 56 0 FreeSans 400 270 0 0 gpio_oeb[43]
port 158 nsew
flabel metal2 s 584160 953270 584216 953726 0 FreeSans 400 90 0 0 gpio_in_h[15]
port 758 nsew
flabel metal2 s 482360 953270 482416 953726 0 FreeSans 400 90 0 0 gpio_in_h[16]
port 757 nsew
flabel metal2 s 430960 953270 431016 953726 0 FreeSans 400 90 0 0 gpio_in_h[17]
port 756 nsew
flabel metal2 s 341960 953270 342016 953726 0 FreeSans 400 90 0 0 gpio_in_h[18]
port 755 nsew
flabel metal2 s 240160 953270 240216 953726 0 FreeSans 400 90 0 0 gpio_in_h[19]
port 754 nsew
flabel metal2 s 188560 953270 188616 953726 0 FreeSans 400 90 0 0 gpio_in_h[20]
port 753 nsew
flabel metal2 s 137160 953270 137216 953726 0 FreeSans 400 90 0 0 gpio_in_h[21]
port 752 nsew
flabel metal2 s 85760 953270 85816 953726 0 FreeSans 400 90 0 0 gpio_in_h[22]
port 751 nsew
flabel metal2 s 34360 953270 34416 953726 0 FreeSans 400 90 0 0 gpio_in_h[23]
port 750 nsew
flabel metal2 s 159910 -400 159966 56 0 FreeSans 400 90 0 0 gpio_in_h[38]
port 735 nsew
flabel metal2 s 268510 -400 268566 56 0 FreeSans 400 90 0 0 gpio_in_h[39]
port 734 nsew
flabel metal2 s 323310 -400 323366 56 0 FreeSans 400 90 0 0 gpio_in_h[40]
port 733 nsew
flabel metal2 s 378110 -400 378166 56 0 FreeSans 400 90 0 0 gpio_in_h[41]
port 732 nsew
flabel metal2 s 432910 -400 432966 56 0 FreeSans 400 90 0 0 gpio_in_h[42]
port 731 nsew
flabel metal2 s 487710 -400 487766 56 0 FreeSans 400 90 0 0 gpio_in_h[43]
port 730 nsew
flabel metal3 633266 422810 633726 427472 0 FreeSans 3200 90 0 0 vccd1
port 28 nsew
flabel metal3 s 633266 786384 633726 791164 0 FreeSans 3200 90 0 0 vdda1
port 24 nsew
flabel metal3 s 633266 471784 633726 476564 0 FreeSans 3200 90 0 0 vdda1
port 24 nsew
flabel metal3 s 633266 383584 633726 388364 0 FreeSans 3200 90 0 0 vssa1
port 26 nsew
flabel metal3 s 533562 953266 538342 953726 0 FreeSans 3200 0 0 0 vssa1
port 26 nsew
flabel metal3 291362 953266 296142 953726 0 FreeSans 3200 0 0 0 vssio
port 19 nsew
flabel metal3 -400 880014 60 884804 0 FreeSans 3200 90 0 0 vccd2
port 29 nsew
flabel metal3 -400 827762 60 832542 0 FreeSans 3200 90 0 0 vddio
port 18 nsew
flabel metal3 -400 785562 60 790342 0 FreeSans 3200 90 0 0 vssa2
port 27 nsew
flabel metal3 -400 440962 60 445742 0 FreeSans 3200 90 0 0 vdda2
port 25 nsew
flabel metal3 -400 68162 60 72942 0 FreeSans 3200 90 0 0 vddio
port 18 nsew
flabel metal3 536984 -400 541764 60 0 FreeSans 3200 0 0 0 vssio
port 19 nsew
flabel metal3 590784 -400 595564 60 0 FreeSans 3200 0 0 0 vdda
port 22 nsew
flabel comment s 107715 141850 108715 141850 0 FreeSans 1120000 60 0 0 example
flabel metal3 s 633266 556035 633726 556249 0 FreeSans 400 0 0 0 analog_noesd_io[8]
port 941 nsew
flabel metal3 -400 906644 60 906704 0 FreeSans 400 0 0 0 gpio_loopback_one[24]
port 837 nsew
flabel metal3 -400 736644 60 736704 0 FreeSans 400 0 0 0 gpio_loopback_one[25]
port 836 nsew
flabel metal3 -400 693644 60 693704 0 FreeSans 400 0 0 0 gpio_loopback_one[26]
port 835 nsew
flabel metal3 -400 650644 60 650704 0 FreeSans 400 0 0 0 gpio_loopback_one[27]
port 834 nsew
flabel metal3 -400 607644 60 607704 0 FreeSans 400 0 0 0 gpio_loopback_one[28]
port 833 nsew
flabel metal3 -400 564644 60 564704 0 FreeSans 400 0 0 0 gpio_loopback_one[29]
port 832 nsew
flabel metal3 -400 521644 60 521704 0 FreeSans 400 0 0 0 gpio_loopback_one[30]
port 831 nsew
flabel metal3 -400 478644 60 478704 0 FreeSans 400 0 0 0 gpio_loopback_one[31]
port 830 nsew
flabel metal3 -400 349644 60 349704 0 FreeSans 400 0 0 0 gpio_loopback_one[32]
port 829 nsew
flabel metal3 -400 306644 60 306704 0 FreeSans 400 0 0 0 gpio_loopback_one[33]
port 828 nsew
flabel metal3 -400 263644 60 263704 0 FreeSans 400 0 0 0 gpio_loopback_one[34]
port 827 nsew
flabel metal3 -400 220644 60 220704 0 FreeSans 400 0 0 0 gpio_loopback_one[35]
port 826 nsew
flabel metal3 -400 177644 60 177704 0 FreeSans 400 0 0 0 gpio_loopback_one[36]
port 825 nsew
flabel metal3 -400 134644 60 134704 0 FreeSans 400 0 0 0 gpio_loopback_one[37]
port 824 nsew
flabel metal2 s 488380 -400 488432 56 0 FreeSans 400 90 0 0 gpio_loopback_one[43]
port 818 nsew
flabel metal2 s 492635 -400 492687 56 0 FreeSans 400 90 0 0 gpio_loopback_zero[43]
port 774 nsew
flabel metal2 s 433580 -400 433632 56 0 FreeSans 400 90 0 0 gpio_loopback_one[42]
port 819 nsew
flabel metal2 s 437778 -400 437830 56 0 FreeSans 400 90 0 0 gpio_loopback_zero[42]
port 775 nsew
flabel metal2 s 378780 -400 378832 56 0 FreeSans 400 90 0 0 gpio_loopback_one[41]
port 820 nsew
flabel metal2 s 382978 -400 383030 56 0 FreeSans 400 90 0 0 gpio_loopback_zero[41]
port 776 nsew
flabel metal2 s 323980 -400 324032 56 0 FreeSans 400 90 0 0 gpio_loopback_one[40]
port 821 nsew
flabel metal2 s 328165 -400 328217 56 0 FreeSans 400 90 0 0 gpio_loopback_zero[40]
port 777 nsew
flabel metal2 s 269180 -400 269232 56 0 FreeSans 400 90 0 0 gpio_loopback_one[39]
port 822 nsew
flabel metal2 s 273360 -400 273412 56 0 FreeSans 400 90 0 0 gpio_loopback_zero[39]
port 778 nsew
flabel metal2 s 160580 -400 160632 56 0 FreeSans 400 90 0 0 gpio_loopback_one[38]
port 823 nsew
flabel metal2 s 163791 -400 163843 56 0 FreeSans 400 90 0 0 gpio_loopback_zero[38]
port 779 nsew
flabel metal2 s 110164 -400 110220 56 0 FreeSans 400 90 0 0 resetb_l
port 37 nsew
flabel metal2 s 99576 -400 99632 56 0 FreeSans 400 90 0 0 resetb_h
port 36 nsew
flabel metal3 -400 53372 60 53442 0 FreeSans 400 0 0 0 por_l
port 35 nsew
flabel metal3 -400 53595 60 53665 0 FreeSans 400 0 0 0 porb_l
port 34 nsew
flabel metal2 s 605082 -400 605134 56 0 FreeSans 400 90 0 0 mask_rev[0]
port 69 nsew
flabel metal3 -400 53147 60 53217 0 FreeSans 400 0 0 0 porb_h
port 33 nsew
flabel metal2 578298 953270 578358 953726 0 FreeSans 400 90 0 0 gpio_loopback_one[15]
port 846 nsew
flabel metal2 478898 953270 478958 953726 0 FreeSans 400 90 0 0 gpio_loopback_one[16]
port 845 nsew
flabel metal2 427698 953270 427758 953726 0 FreeSans 400 90 0 0 gpio_loopback_one[17]
port 844 nsew
flabel metal2 338698 953270 338758 953726 0 FreeSans 400 90 0 0 gpio_loopback_one[18]
port 843 nsew
flabel metal2 234298 953270 234358 953726 0 FreeSans 400 90 0 0 gpio_loopback_one[19]
port 842 nsew
flabel metal2 183098 953270 183158 953726 0 FreeSans 400 90 0 0 gpio_loopback_one[20]
port 841 nsew
flabel metal2 131898 953270 131958 953726 0 FreeSans 400 90 0 0 gpio_loopback_one[21]
port 840 nsew
flabel metal2 80698 953270 80758 953726 0 FreeSans 400 90 0 0 gpio_loopback_one[22]
port 839 nsew
flabel metal2 29498 953270 29558 953726 0 FreeSans 400 90 0 0 gpio_loopback_one[23]
port 838 nsew
flabel metal3 633266 523005 633726 523067 0 FreeSans 400 0 0 0 gpio_loopback_one[7]
port 854 nsew
flabel metal3 633266 346005 633726 346067 0 FreeSans 400 0 0 0 gpio_loopback_one[6]
port 855 nsew
flabel metal3 633266 301005 633726 301067 0 FreeSans 400 0 0 0 gpio_loopback_one[5]
port 856 nsew
flabel metal3 633266 256005 633726 256067 0 FreeSans 400 0 0 0 gpio_loopback_one[4]
port 857 nsew
flabel metal3 633266 211005 633726 211067 0 FreeSans 400 0 0 0 gpio_loopback_one[3]
port 858 nsew
flabel metal3 633266 166005 633726 166067 0 FreeSans 400 0 0 0 gpio_loopback_one[2]
port 859 nsew
flabel metal3 633266 121005 633726 121067 0 FreeSans 400 0 0 0 gpio_loopback_one[1]
port 860 nsew
flabel metal3 633266 76005 633726 76067 0 FreeSans 400 0 0 0 gpio_loopback_one[0]
port 861 nsew
flabel metal2 s 605978 -400 606030 56 0 FreeSans 400 90 0 0 mask_rev[4]
port 65 nsew
flabel metal2 s 606202 -400 606254 56 0 FreeSans 400 90 0 0 mask_rev[5]
port 64 nsew
flabel metal2 s 606426 -400 606478 56 0 FreeSans 400 90 0 0 mask_rev[6]
port 63 nsew
flabel metal2 s 606650 -400 606702 56 0 FreeSans 400 90 0 0 mask_rev[7]
port 62 nsew
flabel metal2 s 606874 -400 606926 56 0 FreeSans 400 90 0 0 mask_rev[8]
port 61 nsew
flabel metal2 s 607098 -400 607150 56 0 FreeSans 400 90 0 0 mask_rev[9]
port 60 nsew
flabel metal2 s 607322 -400 607374 56 0 FreeSans 400 90 0 0 mask_rev[10]
port 59 nsew
flabel metal2 s 607546 -400 607598 56 0 FreeSans 400 90 0 0 mask_rev[11]
port 58 nsew
flabel metal2 s 607770 -400 607822 56 0 FreeSans 400 90 0 0 mask_rev[12]
port 57 nsew
flabel metal2 s 607994 -400 608046 56 0 FreeSans 400 90 0 0 mask_rev[13]
port 60 nsew
flabel metal2 s 608218 -400 608270 56 0 FreeSans 400 90 0 0 mask_rev[14]
port 55 nsew
flabel metal2 s 608442 -400 608494 56 0 FreeSans 400 90 0 0 mask_rev[15]
port 54 nsew
flabel metal2 s 608666 -400 608718 56 0 FreeSans 400 90 0 0 mask_rev[16]
port 53 nsew
flabel metal2 s 608890 -400 608942 56 0 FreeSans 400 90 0 0 mask_rev[17]
port 52 nsew
flabel metal2 s 609114 -400 609166 56 0 FreeSans 400 90 0 0 mask_rev[18]
port 51 nsew
flabel metal2 s 609338 -400 609390 56 0 FreeSans 400 90 0 0 mask_rev[19]
port 50 nsew
flabel metal2 s 609562 -400 609614 56 0 FreeSans 400 90 0 0 mask_rev[20]
port 49 nsew
flabel metal2 s 609786 -400 609838 56 0 FreeSans 400 90 0 0 mask_rev[21]
port 48 nsew
flabel metal2 s 610010 -400 610062 56 0 FreeSans 400 90 0 0 mask_rev[22]
port 47 nsew
flabel metal2 s 610234 -400 610286 56 0 FreeSans 400 90 0 0 mask_rev[23]
port 46 nsew
flabel metal2 s 610458 -400 610510 56 0 FreeSans 400 90 0 0 mask_rev[24]
port 45 nsew
flabel metal2 s 610682 -400 610734 56 0 FreeSans 400 90 0 0 mask_rev[25]
port 44 nsew
flabel metal2 s 610906 -400 610958 56 0 FreeSans 400 90 0 0 mask_rev[26]
port 43 nsew
flabel metal2 s 611130 -400 611182 56 0 FreeSans 400 90 0 0 mask_rev[27]
port 42 nsew
flabel metal2 s 611354 -400 611406 56 0 FreeSans 400 90 0 0 mask_rev[28]
port 41 nsew
flabel metal2 s 611578 -400 611630 56 0 FreeSans 400 90 0 0 mask_rev[29]
port 40 nsew
flabel metal2 s 611802 -400 611854 56 0 FreeSans 400 90 0 0 mask_rev[30]
port 39 nsew
flabel metal2 s 612026 -400 612078 56 0 FreeSans 400 90 0 0 mask_rev[31]
port 38 nsew
flabel metal2 s 605754 -400 605806 56 0 FreeSans 400 90 0 0 mask_rev[3]
port 66 nsew
flabel metal2 s 605530 -400 605582 56 0 FreeSans 400 90 0 0 mask_rev[2]
port 67 nsew
flabel metal2 s 605306 -400 605358 56 0 FreeSans 400 90 0 0 mask_rev[1]
port 68 nsew
flabel metal3 -400 734644 60 734704 0 FreeSans 400 0 0 0 gpio_loopback_zero[25]
port 792 nsew
flabel metal3 -400 648644 60 648704 0 FreeSans 400 0 0 0 gpio_loopback_zero[27]
port 790 nsew
flabel metal3 -400 562644 60 562704 0 FreeSans 400 0 0 0 gpio_loopback_zero[29]
port 788 nsew
flabel metal3 -400 476644 60 476704 0 FreeSans 400 0 0 0 gpio_loopback_zero[31]
port 786 nsew
flabel metal3 -400 304644 60 304704 0 FreeSans 400 0 0 0 gpio_loopback_zero[33]
port 784 nsew
flabel metal3 -400 218644 60 218704 0 FreeSans 400 0 0 0 gpio_loopback_zero[35]
port 782 nsew
flabel metal3 -400 132644 60 132704 0 FreeSans 400 0 0 0 gpio_loopback_zero[37]
port 780 nsew
flabel metal3 -400 904644 60 904704 0 FreeSans 400 0 0 0 gpio_loopback_zero[24]
port 793 nsew
flabel metal3 -400 691644 60 691704 0 FreeSans 400 0 0 0 gpio_loopback_zero[26]
port 791 nsew
flabel metal3 -400 605644 60 605704 0 FreeSans 400 0 0 0 gpio_loopback_zero[28]
port 789 nsew
flabel metal3 -400 519644 60 519704 0 FreeSans 400 0 0 0 gpio_loopback_zero[30]
port 787 nsew
flabel metal3 -400 347644 60 347704 0 FreeSans 400 0 0 0 gpio_loopback_zero[32]
port 785 nsew
flabel metal3 -400 261644 60 261704 0 FreeSans 400 0 0 0 gpio_loopback_zero[34]
port 783 nsew
flabel metal3 -400 175644 60 175704 0 FreeSans 400 0 0 0 gpio_loopback_zero[36]
port 781 nsew
flabel metal2 147030 -400 147086 56 0 FreeSans 400 270 0 0 gpio_slow_sel[38]
port 339 nsew
flabel metal2 145190 -400 145246 56 0 FreeSans 400 270 0 0 gpio_in[38]
port 691 nsew
flabel metal3 46784 -400 51564 60 0 FreeSans 3200 0 0 0 vssa
port 23 nsew
flabel metal3 633266 61238 633726 61366 0 FreeSans 400 0 0 0 analog_io[0]
port 905 nsew
flabel metal3 633266 63035 633726 63249 0 FreeSans 400 0 0 0 analog_noesd_io[0]
port 949 nsew
flabel metal3 633266 108235 633726 108449 0 FreeSans 400 0 0 0 analog_noesd_io[1]
port 948 nsew
flabel metal3 633266 106438 633726 106566 0 FreeSans 400 0 0 0 analog_io[1]
port 904 nsew
flabel metal3 633266 151438 633726 151566 0 FreeSans 400 0 0 0 analog_io[2]
port 903 nsew
flabel metal3 633266 153235 633726 153449 0 FreeSans 400 0 0 0 analog_noesd_io[2]
port 947 nsew
flabel metal3 633266 196638 633726 196766 0 FreeSans 400 0 0 0 analog_io[3]
port 902 nsew
flabel metal3 633266 198435 633726 198649 0 FreeSans 400 0 0 0 analog_noesd_io[3]
port 946 nsew
flabel metal3 633266 241638 633726 241766 0 FreeSans 400 0 0 0 analog_io[4]
port 901 nsew
flabel metal3 633266 243435 633726 243649 0 FreeSans 400 0 0 0 analog_noesd_io[4]
port 945 nsew
flabel metal3 633266 286638 633726 286766 0 FreeSans 400 0 0 0 analog_io[5]
port 900 nsew
flabel metal3 633266 288435 633726 288649 0 FreeSans 400 0 0 0 analog_noesd_io[5]
port 944 nsew
flabel metal3 633266 331838 633726 331966 0 FreeSans 400 0 0 0 analog_io[6]
port 899 nsew
flabel metal3 633266 333635 633726 333849 0 FreeSans 400 0 0 0 analog_noesd_io[6]
port 943 nsew
flabel metal3 s 633266 509038 633726 509166 0 FreeSans 400 0 0 0 analog_io[7]
port 898 nsew
flabel metal3 s 633266 510835 633726 511049 0 FreeSans 400 0 0 0 analog_noesd_io[7]
port 942 nsew
flabel metal3 s 633266 554238 633726 554366 0 FreeSans 400 0 0 0 analog_io[8]
port 897 nsew
flabel metal3 s 633266 599238 633726 599366 0 FreeSans 400 0 0 0 analog_io[9]
port 896 nsew
flabel metal3 s 633266 601035 633726 601249 0 FreeSans 400 0 0 0 analog_noesd_io[9]
port 940 nsew
flabel metal3 s 633266 644438 633726 644566 0 FreeSans 400 0 0 0 analog_io[10]
port 895 nsew
flabel metal3 s 633266 646235 633726 646449 0 FreeSans 400 0 0 0 analog_noesd_io[10]
port 939 nsew
flabel metal3 s 633266 689438 633726 689566 0 FreeSans 400 0 0 0 analog_io[11]
port 894 nsew
flabel metal3 s 633266 691235 633726 691449 0 FreeSans 400 0 0 0 analog_noesd_io[11]
port 938 nsew
flabel metal3 s 633266 734438 633726 734566 0 FreeSans 400 0 0 0 analog_io[12]
port 893 nsew
flabel metal3 s 633266 823638 633726 823766 0 FreeSans 400 0 0 0 analog_io[13]
port 892 nsew
flabel metal3 s 633266 912838 633726 912966 0 FreeSans 400 0 0 0 analog_io[14]
port 891 nsew
flabel metal3 s 633266 736235 633726 736449 0 FreeSans 400 0 0 0 analog_noesd_io[12]
port 937 nsew
flabel metal3 s 633266 825435 633726 825649 0 FreeSans 400 0 0 0 analog_noesd_io[13]
port 936 nsew
flabel metal3 s 633266 914635 633726 914849 0 FreeSans 400 0 0 0 analog_noesd_io[14]
port 935 nsew
flabel metal2 s 596360 953270 596488 953726 0 FreeSans 400 90 0 0 analog_io[15]
port 890 nsew
flabel metal2 s 494560 953270 494688 953726 0 FreeSans 400 90 0 0 analog_io[16]
port 889 nsew
flabel metal2 s 443160 953270 443288 953726 0 FreeSans 400 90 0 0 analog_io[17]
port 888 nsew
flabel metal2 s 354160 953270 354288 953726 0 FreeSans 400 90 0 0 analog_io[18]
port 887 nsew
flabel metal2 s 252360 953270 252488 953726 0 FreeSans 400 90 0 0 analog_io[19]
port 886 nsew
flabel metal2 s 200760 953270 200888 953726 0 FreeSans 400 90 0 0 analog_io[20]
port 885 nsew
flabel metal2 s 149360 953270 149488 953726 0 FreeSans 400 90 0 0 analog_io[21]
port 884 nsew
flabel metal2 s 97960 953270 98088 953726 0 FreeSans 400 90 0 0 analog_io[22]
port 883 nsew
flabel metal2 s 46560 953270 46688 953726 0 FreeSans 400 90 0 0 analog_io[23]
port 882 nsew
flabel metal2 s 594477 953270 594691 953726 0 FreeSans 400 90 0 0 analog_noesd_io[15]
port 934 nsew
flabel metal2 s 492677 953270 492891 953726 0 FreeSans 400 90 0 0 analog_noesd_io[16]
port 933 nsew
flabel metal2 s 441277 953270 441491 953726 0 FreeSans 400 90 0 0 analog_noesd_io[17]
port 932 nsew
flabel metal2 s 352277 953270 352491 953726 0 FreeSans 400 90 0 0 analog_noesd_io[18]
port 931 nsew
flabel metal2 s 250477 953270 250691 953726 0 FreeSans 400 90 0 0 analog_noesd_io[19]
port 930 nsew
flabel metal2 s 198877 953270 199091 953726 0 FreeSans 400 90 0 0 analog_noesd_io[20]
port 929 nsew
flabel metal2 s 147477 953270 147691 953726 0 FreeSans 400 90 0 0 analog_noesd_io[21]
port 928 nsew
flabel metal2 s 96077 953270 96291 953726 0 FreeSans 400 90 0 0 analog_noesd_io[22]
port 927 nsew
flabel metal2 s 44677 953270 44891 953726 0 FreeSans 400 90 0 0 analog_noesd_io[23]
port 926 nsew
flabel metal3 s -400 754760 60 754888 0 FreeSans 400 0 0 0 analog_io[25]
port 880 nsew
flabel metal3 s -400 711560 60 711688 0 FreeSans 400 0 0 0 analog_io[26]
port 879 nsew
flabel metal3 s -400 668360 60 668488 0 FreeSans 400 0 0 0 analog_io[27]
port 878 nsew
flabel metal3 s -400 625160 60 625288 0 FreeSans 400 0 0 0 analog_io[28]
port 877 nsew
flabel metal3 s -400 581960 60 582088 0 FreeSans 400 0 0 0 analog_io[29]
port 876 nsew
flabel metal3 s -400 538760 60 538888 0 FreeSans 400 0 0 0 analog_io[30]
port 875 nsew
flabel metal3 s -400 495560 60 495688 0 FreeSans 400 0 0 0 analog_io[31]
port 874 nsew
flabel metal3 s -400 367960 60 368088 0 FreeSans 400 0 0 0 analog_io[32]
port 873 nsew
flabel metal3 s -400 324760 60 324888 0 FreeSans 400 0 0 0 analog_io[33]
port 872 nsew
flabel metal3 s -400 281560 60 281688 0 FreeSans 400 0 0 0 analog_io[34]
port 871 nsew
flabel metal3 s -400 238360 60 238488 0 FreeSans 400 0 0 0 analog_io[35]
port 870 nsew
flabel metal3 s -400 195160 60 195288 0 FreeSans 400 0 0 0 analog_io[36]
port 869 nsew
flabel metal3 s -400 151960 60 152088 0 FreeSans 400 0 0 0 analog_io[37]
port 868 nsew
flabel metal3 s -400 752877 60 753091 0 FreeSans 400 0 0 0 analog_noesd_io[25]
port 924 nsew
flabel metal3 s -400 709677 60 709891 0 FreeSans 400 0 0 0 analog_noesd_io[26]
port 923 nsew
flabel metal3 s -400 666477 60 666691 0 FreeSans 400 0 0 0 analog_noesd_io[27]
port 922 nsew
flabel metal3 s -400 623277 60 623491 0 FreeSans 400 0 0 0 analog_noesd_io[28]
port 921 nsew
flabel metal3 s -400 580077 60 580291 0 FreeSans 400 0 0 0 analog_noesd_io[29]
port 920 nsew
flabel metal3 s -400 536877 60 537091 0 FreeSans 400 0 0 0 analog_noesd_io[30]
port 919 nsew
flabel metal3 s -400 366077 60 366291 0 FreeSans 400 0 0 0 analog_noesd_io[32]
port 917 nsew
flabel metal3 s -400 322877 60 323091 0 FreeSans 400 0 0 0 analog_noesd_io[33]
port 916 nsew
flabel metal3 s -400 279677 60 279891 0 FreeSans 400 0 0 0 analog_noesd_io[34]
port 915 nsew
flabel metal3 s -400 236477 60 236691 0 FreeSans 400 0 0 0 analog_noesd_io[35]
port 914 nsew
flabel metal3 s -400 193277 60 193491 0 FreeSans 400 0 0 0 analog_noesd_io[36]
port 913 nsew
flabel metal3 s -400 150077 60 150291 0 FreeSans 400 0 0 0 analog_noesd_io[37]
port 912 nsew
flabel metal2 s 256238 -400 256366 56 0 FreeSans 400 90 0 0 analog_io[39]
port 866 nsew
flabel metal2 s 311038 -400 311166 56 0 FreeSans 400 90 0 0 analog_io[40]
port 865 nsew
flabel metal2 s 365838 -400 365966 56 0 FreeSans 400 90 0 0 analog_io[41]
port 864 nsew
flabel metal2 s 420638 -400 420766 56 0 FreeSans 400 90 0 0 analog_io[42]
port 863 nsew
flabel metal2 s 475438 -400 475566 56 0 FreeSans 400 90 0 0 analog_io[43]
port 862 nsew
flabel metal2 s 258035 -400 258249 56 0 FreeSans 400 90 0 0 analog_noesd_io[39]
port 910 nsew
flabel metal2 s 312835 -400 313049 56 0 FreeSans 400 90 0 0 analog_noesd_io[40]
port 909 nsew
flabel metal2 s 367635 -400 367849 56 0 FreeSans 400 90 0 0 analog_noesd_io[41]
port 908 nsew
flabel metal2 s 422435 -400 422649 56 0 FreeSans 400 90 0 0 analog_noesd_io[42]
port 907 nsew
flabel metal2 s 477235 -400 477449 56 0 FreeSans 400 90 0 0 analog_noesd_io[43]
port 906 nsew
flabel metal2 s 149435 -400 149649 56 0 FreeSans 400 90 0 0 analog_noesd_io[38]
port 911 nsew
flabel metal2 s 147638 -400 147766 56 0 FreeSans 400 90 0 0 analog_io[38]
port 867 nsew
flabel metal2 148870 -400 148926 56 0 FreeSans 400 270 0 0 gpio_dm1[38]
port 603 nsew
flabel metal2 150710 -400 150766 56 0 FreeSans 400 270 0 0 gpio_dm0[38]
port 559 nsew
flabel metal3 s -400 493677 60 493891 0 FreeSans 400 0 0 0 analog_noesd_io[31]
port 918 nsew
flabel metal3 s 633266 373606 633726 378386 0 FreeSans 3200 90 0 0 vssa1
port 26 nsew
flabel metal3 633266 417722 633726 422512 0 FreeSans 3200 90 0 0 vssd1
port 30 nsew
flabel metal3 633266 427762 633726 432562 0 FreeSans 3200 90 0 0 vssd1
port 30 nsew
flabel metal3 s 633266 461804 633726 466584 0 FreeSans 3200 90 0 0 vdda1
port 24 nsew
flabel metal3 633266 568006 633726 568068 0 FreeSans 400 0 0 0 gpio_loopback_one[8]
port 853 nsew
flabel metal3 633266 613006 633726 613068 0 FreeSans 400 0 0 0 gpio_loopback_one[9]
port 852 nsew
flabel metal3 633266 658006 633726 658068 0 FreeSans 400 0 0 0 gpio_loopback_one[10]
port 851 nsew
flabel metal3 633266 703006 633726 703068 0 FreeSans 400 0 0 0 gpio_loopback_one[11]
port 850 nsew
flabel metal3 633266 748006 633726 748068 0 FreeSans 400 0 0 0 gpio_loopback_one[12]
port 849 nsew
flabel metal3 s 633266 776406 633726 781186 0 FreeSans 3200 90 0 0 vdda1
port 24 nsew
flabel metal3 633266 837006 633726 837068 0 FreeSans 400 0 0 0 gpio_loopback_one[13]
port 848 nsew
flabel metal3 633266 927006 633726 927068 0 FreeSans 400 0 0 0 gpio_loopback_one[14]
port 847 nsew
flabel metal3 s 543542 953266 548322 953726 0 FreeSans 3200 0 0 0 vssa1
port 26 nsew
flabel metal3 301342 953266 306122 953726 0 FreeSans 3200 0 0 0 vssio
port 19 nsew
flabel metal3 -400 875054 60 879716 0 FreeSans 3200 90 0 0 vssd2
port 31 nsew
flabel metal3 -400 869964 60 874764 0 FreeSans 3200 90 0 0 vccd2
port 29 nsew
flabel metal3 -400 837742 60 842522 0 FreeSans 3200 90 0 0 vddio
port 18 nsew
flabel metal3 -400 795542 60 800322 0 FreeSans 3200 90 0 0 vssa2
port 27 nsew
flabel metal3 s -400 757272 60 757342 0 FreeSans 400 0 0 0 gpio_in[25]
port 704 nsew
flabel metal3 s -400 755432 60 755502 0 FreeSans 400 0 0 0 gpio_slow_sel[25]
port 352 nsew
flabel metal3 s -400 753592 60 753662 0 FreeSans 400 0 0 0 gpio_dm1[25]
port 616 nsew
flabel metal3 s -400 752396 60 752466 0 FreeSans 400 0 0 0 gpio_analog_en[25]
port 440 nsew
flabel metal3 s -400 751752 60 751822 0 FreeSans 400 0 0 0 gpio_dm0[25]
port 572 nsew
flabel metal3 s -400 751108 60 751178 0 FreeSans 400 0 0 0 gpio_analog_pol[25]
port 528 nsew
flabel metal3 s -400 750556 60 750626 0 FreeSans 400 0 0 0 gpio_inp_dis[25]
port 220 nsew
flabel metal3 s -400 748072 60 748142 0 FreeSans 400 0 0 0 gpio_analog_sel[25]
port 484 nsew
flabel metal3 s -400 747428 60 747498 0 FreeSans 400 0 0 0 gpio_dm2[25]
port 660 nsew
flabel metal3 s -400 746784 60 746854 0 FreeSans 400 0 0 0 gpio_holdover[25]
port 396 nsew
flabel metal3 s -400 746232 60 746302 0 FreeSans 400 0 0 0 gpio_out[25]
port 132 nsew
flabel metal3 s -400 744392 60 744462 0 FreeSans 400 0 0 0 gpio_vtrip_sel[25]
port 308 nsew
flabel metal3 s -400 743748 60 743818 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[25]
port 264 nsew
flabel metal3 s -400 743104 60 743174 0 FreeSans 400 0 0 0 gpio_oeb[25]
port 176 nsew
flabel metal3 s -400 742552 60 742622 0 FreeSans 400 0 0 0 gpio_in_h[25]
port 748 nsew
flabel metal3 s -400 714072 60 714142 0 FreeSans 400 0 0 0 gpio_in[26]
port 703 nsew
flabel metal3 s -400 712232 60 712302 0 FreeSans 400 0 0 0 gpio_slow_sel[26]
port 351 nsew
flabel metal3 s -400 710392 60 710462 0 FreeSans 400 0 0 0 gpio_dm1[26]
port 615 nsew
flabel metal3 s -400 709196 60 709266 0 FreeSans 400 0 0 0 gpio_analog_en[26]
port 439 nsew
flabel metal3 s -400 708552 60 708622 0 FreeSans 400 0 0 0 gpio_dm0[26]
port 571 nsew
flabel metal3 s -400 707908 60 707978 0 FreeSans 400 0 0 0 gpio_analog_pol[26]
port 527 nsew
flabel metal3 s -400 707356 60 707426 0 FreeSans 400 0 0 0 gpio_inp_dis[26]
port 219 nsew
flabel metal3 s -400 704872 60 704942 0 FreeSans 400 0 0 0 gpio_analog_sel[26]
port 483 nsew
flabel metal3 s -400 704228 60 704298 0 FreeSans 400 0 0 0 gpio_dm2[26]
port 659 nsew
flabel metal3 s -400 703584 60 703654 0 FreeSans 400 0 0 0 gpio_holdover[26]
port 395 nsew
flabel metal3 s -400 703032 60 703102 0 FreeSans 400 0 0 0 gpio_out[26]
port 131 nsew
flabel metal3 s -400 701192 60 701262 0 FreeSans 400 0 0 0 gpio_vtrip_sel[26]
port 307 nsew
flabel metal3 s -400 700548 60 700618 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[26]
port 263 nsew
flabel metal3 s -400 699904 60 699974 0 FreeSans 400 0 0 0 gpio_oeb[26]
port 175 nsew
flabel metal3 s -400 699352 60 699422 0 FreeSans 400 0 0 0 gpio_in_h[26]
port 747 nsew
flabel metal3 s -400 141592 60 141662 0 FreeSans 400 0 0 0 gpio_vtrip_sel[37]
port 296 nsew
flabel metal3 s -400 149596 60 149666 0 FreeSans 400 0 0 0 gpio_analog_en[37]
port 428 nsew
flabel metal3 s -400 148308 60 148378 0 FreeSans 400 0 0 0 gpio_analog_pol[37]
port 516 nsew
flabel metal3 s -400 145272 60 145342 0 FreeSans 400 0 0 0 gpio_analog_sel[37]
port 472 nsew
flabel metal3 s -400 148952 60 149022 0 FreeSans 400 0 0 0 gpio_dm0[37]
port 560 nsew
flabel metal3 s -400 144628 60 144698 0 FreeSans 400 0 0 0 gpio_dm2[37]
port 648 nsew
flabel metal3 s -400 143984 60 144054 0 FreeSans 400 0 0 0 gpio_holdover[37]
port 384 nsew
flabel metal3 s -400 140948 60 141018 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[37]
port 252 nsew
flabel metal3 s -400 140304 60 140374 0 FreeSans 400 0 0 0 gpio_oeb[37]
port 164 nsew
flabel metal3 s -400 143432 60 143502 0 FreeSans 400 0 0 0 gpio_out[37]
port 120 nsew
flabel metal3 s -400 147756 60 147826 0 FreeSans 400 0 0 0 gpio_inp_dis[37]
port 208 nsew
flabel metal3 s -400 139752 60 139822 0 FreeSans 400 0 0 0 gpio_in_h[37]
port 736 nsew
flabel metal3 s -400 150792 60 150862 0 FreeSans 400 0 0 0 gpio_dm1[37]
port 604 nsew
flabel metal3 s -400 152632 60 152702 0 FreeSans 400 0 0 0 gpio_slow_sel[37]
port 340 nsew
flabel metal3 s -400 154472 60 154542 0 FreeSans 400 0 0 0 gpio_in[37]
port 692 nsew
flabel metal3 s -400 187828 60 187898 0 FreeSans 400 0 0 0 gpio_dm2[36]
port 649 nsew
flabel metal3 s -400 187184 60 187254 0 FreeSans 400 0 0 0 gpio_holdover[36]
port 385 nsew
flabel metal3 s -400 184148 60 184218 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[36]
port 253 nsew
flabel metal3 s -400 190956 60 191026 0 FreeSans 400 0 0 0 gpio_inp_dis[36]
port 209 nsew
flabel metal3 s -400 183504 60 183574 0 FreeSans 400 0 0 0 gpio_oeb[36]
port 165 nsew
flabel metal3 s -400 186632 60 186702 0 FreeSans 400 0 0 0 gpio_out[36]
port 121 nsew
flabel metal3 s -400 184792 60 184862 0 FreeSans 400 0 0 0 gpio_vtrip_sel[36]
port 297 nsew
flabel metal3 s -400 192796 60 192866 0 FreeSans 400 0 0 0 gpio_analog_en[36]
port 429 nsew
flabel metal3 s -400 191508 60 191578 0 FreeSans 400 0 0 0 gpio_analog_pol[36]
port 517 nsew
flabel metal3 s -400 188472 60 188542 0 FreeSans 400 0 0 0 gpio_analog_sel[36]
port 473 nsew
flabel metal3 s -400 192152 60 192222 0 FreeSans 400 0 0 0 gpio_dm0[36]
port 561 nsew
flabel metal3 s -400 182952 60 183022 0 FreeSans 400 0 0 0 gpio_in_h[36]
port 737 nsew
flabel metal3 s -400 193992 60 194062 0 FreeSans 400 0 0 0 gpio_dm1[36]
port 605 nsew
flabel metal3 s -400 195832 60 195902 0 FreeSans 400 0 0 0 gpio_slow_sel[36]
port 341 nsew
flabel metal3 s -400 197672 60 197742 0 FreeSans 400 0 0 0 gpio_in[36]
port 693 nsew
flabel metal3 s -400 235996 60 236066 0 FreeSans 400 0 0 0 gpio_analog_en[35]
port 430 nsew
flabel metal3 s -400 234708 60 234778 0 FreeSans 400 0 0 0 gpio_analog_pol[35]
port 518 nsew
flabel metal3 s -400 231672 60 231742 0 FreeSans 400 0 0 0 gpio_analog_sel[35]
port 474 nsew
flabel metal3 s -400 235352 60 235422 0 FreeSans 400 0 0 0 gpio_dm0[35]
port 562 nsew
flabel metal3 s -400 231028 60 231098 0 FreeSans 400 0 0 0 gpio_dm2[35]
port 650 nsew
flabel metal3 s -400 230384 60 230454 0 FreeSans 400 0 0 0 gpio_holdover[35]
port 386 nsew
flabel metal3 s -400 227348 60 227418 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[35]
port 254 nsew
flabel metal3 s -400 234156 60 234226 0 FreeSans 400 0 0 0 gpio_inp_dis[35]
port 210 nsew
flabel metal3 s -400 226704 60 226774 0 FreeSans 400 0 0 0 gpio_oeb[35]
port 166 nsew
flabel metal3 s -400 229832 60 229902 0 FreeSans 400 0 0 0 gpio_out[35]
port 122 nsew
flabel metal3 s -400 227992 60 228062 0 FreeSans 400 0 0 0 gpio_vtrip_sel[35]
port 298 nsew
flabel metal3 s -400 226152 60 226222 0 FreeSans 400 0 0 0 gpio_in_h[35]
port 738 nsew
flabel metal3 s -400 237192 60 237262 0 FreeSans 400 0 0 0 gpio_dm1[35]
port 606 nsew
flabel metal3 s -400 239032 60 239102 0 FreeSans 400 0 0 0 gpio_slow_sel[35]
port 342 nsew
flabel metal3 s -400 240872 60 240942 0 FreeSans 400 0 0 0 gpio_in[35]
port 694 nsew
flabel metal3 s -400 279196 60 279266 0 FreeSans 400 0 0 0 gpio_analog_en[34]
port 431 nsew
flabel metal3 s -400 277908 60 277978 0 FreeSans 400 0 0 0 gpio_analog_pol[34]
port 519 nsew
flabel metal3 s -400 274872 60 274942 0 FreeSans 400 0 0 0 gpio_analog_sel[34]
port 475 nsew
flabel metal3 s -400 278552 60 278622 0 FreeSans 400 0 0 0 gpio_dm0[34]
port 563 nsew
flabel metal3 s -400 274228 60 274298 0 FreeSans 400 0 0 0 gpio_dm2[34]
port 651 nsew
flabel metal3 s -400 273584 60 273654 0 FreeSans 400 0 0 0 gpio_holdover[34]
port 387 nsew
flabel metal3 s -400 270548 60 270618 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[34]
port 255 nsew
flabel metal3 s -400 277356 60 277426 0 FreeSans 400 0 0 0 gpio_inp_dis[34]
port 211 nsew
flabel metal3 s -400 269904 60 269974 0 FreeSans 400 0 0 0 gpio_oeb[34]
port 167 nsew
flabel metal3 s -400 273032 60 273102 0 FreeSans 400 0 0 0 gpio_out[34]
port 123 nsew
flabel metal3 s -400 271192 60 271262 0 FreeSans 400 0 0 0 gpio_vtrip_sel[34]
port 299 nsew
flabel metal3 s -400 269352 60 269422 0 FreeSans 400 0 0 0 gpio_in_h[34]
port 739 nsew
flabel metal3 s -400 280392 60 280462 0 FreeSans 400 0 0 0 gpio_dm1[34]
port 607 nsew
flabel metal3 s -400 282232 60 282302 0 FreeSans 400 0 0 0 gpio_slow_sel[34]
port 343 nsew
flabel metal3 s -400 284072 60 284142 0 FreeSans 400 0 0 0 gpio_in[34]
port 695 nsew
flabel metal3 s -400 322396 60 322466 0 FreeSans 400 0 0 0 gpio_analog_en[33]
port 432 nsew
flabel metal3 s -400 318072 60 318142 0 FreeSans 400 0 0 0 gpio_analog_sel[33]
port 476 nsew
flabel metal3 s -400 317428 60 317498 0 FreeSans 400 0 0 0 gpio_dm2[33]
port 652 nsew
flabel metal3 s -400 321752 60 321822 0 FreeSans 400 0 0 0 gpio_dm0[33]
port 564 nsew
flabel metal3 s -400 316784 60 316854 0 FreeSans 400 0 0 0 gpio_holdover[33]
port 388 nsew
flabel metal3 s -400 313748 60 313818 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[33]
port 256 nsew
flabel metal3 s -400 320556 60 320626 0 FreeSans 400 0 0 0 gpio_inp_dis[33]
port 212 nsew
flabel metal3 s -400 313104 60 313174 0 FreeSans 400 0 0 0 gpio_oeb[33]
port 168 nsew
flabel metal3 s -400 316232 60 316302 0 FreeSans 400 0 0 0 gpio_out[33]
port 124 nsew
flabel metal3 s -400 314392 60 314462 0 FreeSans 400 0 0 0 gpio_vtrip_sel[33]
port 300 nsew
flabel metal3 s -400 312552 60 312622 0 FreeSans 400 0 0 0 gpio_in_h[33]
port 740 nsew
flabel metal3 s -400 321108 60 321178 0 FreeSans 400 0 0 0 gpio_analog_pol[33]
port 520 nsew
flabel metal3 s -400 323592 60 323662 0 FreeSans 400 0 0 0 gpio_dm1[33]
port 608 nsew
flabel metal3 s -400 325432 60 325502 0 FreeSans 400 0 0 0 gpio_slow_sel[33]
port 344 nsew
flabel metal3 s -400 327272 60 327342 0 FreeSans 400 0 0 0 gpio_in[33]
port 696 nsew
flabel metal3 s -400 365596 60 365666 0 FreeSans 400 0 0 0 gpio_analog_en[32]
port 433 nsew
flabel metal3 s -400 364308 60 364378 0 FreeSans 400 0 0 0 gpio_analog_pol[32]
port 521 nsew
flabel metal3 s -400 361272 60 361342 0 FreeSans 400 0 0 0 gpio_analog_sel[32]
port 477 nsew
flabel metal3 s -400 364952 60 365022 0 FreeSans 400 0 0 0 gpio_dm0[32]
port 565 nsew
flabel metal3 s -400 360628 60 360698 0 FreeSans 400 0 0 0 gpio_dm2[32]
port 653 nsew
flabel metal3 s -400 359984 60 360054 0 FreeSans 400 0 0 0 gpio_holdover[32]
port 389 nsew
flabel metal3 s -400 356948 60 357018 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[32]
port 257 nsew
flabel metal3 s -400 363756 60 363826 0 FreeSans 400 0 0 0 gpio_inp_dis[32]
port 213 nsew
flabel metal3 s -400 356304 60 356374 0 FreeSans 400 0 0 0 gpio_oeb[32]
port 169 nsew
flabel metal3 s -400 359432 60 359502 0 FreeSans 400 0 0 0 gpio_out[32]
port 125 nsew
flabel metal3 s -400 357592 60 357662 0 FreeSans 400 0 0 0 gpio_vtrip_sel[32]
port 301 nsew
flabel metal3 s -400 355752 60 355822 0 FreeSans 400 0 0 0 gpio_in_h[32]
port 741 nsew
flabel metal3 s -400 366792 60 366862 0 FreeSans 400 0 0 0 gpio_dm1[32]
port 609 nsew
flabel metal3 s -400 368632 60 368702 0 FreeSans 400 0 0 0 gpio_slow_sel[32]
port 345 nsew
flabel metal3 s -400 370472 60 370542 0 FreeSans 400 0 0 0 gpio_in[32]
port 697 nsew
flabel metal3 s -400 493196 60 493266 0 FreeSans 400 0 0 0 gpio_analog_en[31]
port 434 nsew
flabel metal3 s -400 491908 60 491978 0 FreeSans 400 0 0 0 gpio_analog_pol[31]
port 522 nsew
flabel metal3 s -400 488872 60 488942 0 FreeSans 400 0 0 0 gpio_analog_sel[31]
port 478 nsew
flabel metal3 s -400 492552 60 492622 0 FreeSans 400 0 0 0 gpio_dm0[31]
port 566 nsew
flabel metal3 s -400 488228 60 488298 0 FreeSans 400 0 0 0 gpio_dm2[31]
port 654 nsew
flabel metal3 s -400 487584 60 487654 0 FreeSans 400 0 0 0 gpio_holdover[31]
port 390 nsew
flabel metal3 s -400 484548 60 484618 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[31]
port 258 nsew
flabel metal3 s -400 491356 60 491426 0 FreeSans 400 0 0 0 gpio_inp_dis[31]
port 214 nsew
flabel metal3 s -400 483904 60 483974 0 FreeSans 400 0 0 0 gpio_oeb[31]
port 170 nsew
flabel metal3 s -400 487032 60 487102 0 FreeSans 400 0 0 0 gpio_out[31]
port 126 nsew
flabel metal3 s -400 485192 60 485262 0 FreeSans 400 0 0 0 gpio_vtrip_sel[31]
port 302 nsew
flabel metal3 s -400 483352 60 483422 0 FreeSans 400 0 0 0 gpio_in_h[31]
port 742 nsew
flabel metal3 s -400 494392 60 494462 0 FreeSans 400 0 0 0 gpio_dm1[31]
port 610 nsew
flabel metal3 s -400 496232 60 496302 0 FreeSans 400 0 0 0 gpio_slow_sel[31]
port 346 nsew
flabel metal3 s -400 498072 60 498142 0 FreeSans 400 0 0 0 gpio_in[31]
port 698 nsew
flabel metal3 s -400 535752 60 535822 0 FreeSans 400 0 0 0 gpio_dm0[30]
port 567 nsew
flabel metal3 s -400 531428 60 531498 0 FreeSans 400 0 0 0 gpio_dm2[30]
port 655 nsew
flabel metal3 s -400 530784 60 530854 0 FreeSans 400 0 0 0 gpio_holdover[30]
port 391 nsew
flabel metal3 s -400 527748 60 527818 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[30]
port 259 nsew
flabel metal3 s -400 534556 60 534626 0 FreeSans 400 0 0 0 gpio_inp_dis[30]
port 215 nsew
flabel metal3 s -400 527104 60 527174 0 FreeSans 400 0 0 0 gpio_oeb[30]
port 171 nsew
flabel metal3 s -400 530232 60 530302 0 FreeSans 400 0 0 0 gpio_out[30]
port 127 nsew
flabel metal3 s -400 528392 60 528462 0 FreeSans 400 0 0 0 gpio_vtrip_sel[30]
port 303 nsew
flabel metal3 s -400 536396 60 536466 0 FreeSans 400 0 0 0 gpio_analog_en[30]
port 435 nsew
flabel metal3 s -400 535108 60 535178 0 FreeSans 400 0 0 0 gpio_analog_pol[30]
port 523 nsew
flabel metal3 s -400 532072 60 532142 0 FreeSans 400 0 0 0 gpio_analog_sel[30]
port 479 nsew
flabel metal3 s -400 526552 60 526622 0 FreeSans 400 0 0 0 gpio_in_h[30]
port 743 nsew
flabel metal3 s -400 537592 60 537662 0 FreeSans 400 0 0 0 gpio_dm1[30]
port 611 nsew
flabel metal3 s -400 539432 60 539502 0 FreeSans 400 0 0 0 gpio_slow_sel[30]
port 347 nsew
flabel metal3 s -400 541272 60 541342 0 FreeSans 400 0 0 0 gpio_in[30]
port 699 nsew
flabel metal3 s -400 575272 60 575342 0 FreeSans 400 0 0 0 gpio_analog_sel[29]
port 480 nsew
flabel metal3 s -400 574628 60 574698 0 FreeSans 400 0 0 0 gpio_dm2[29]
port 656 nsew
flabel metal3 s -400 573984 60 574054 0 FreeSans 400 0 0 0 gpio_holdover[29]
port 392 nsew
flabel metal3 s -400 570948 60 571018 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[29]
port 260 nsew
flabel metal3 s -400 570304 60 570374 0 FreeSans 400 0 0 0 gpio_oeb[29]
port 172 nsew
flabel metal3 s -400 573432 60 573502 0 FreeSans 400 0 0 0 gpio_out[29]
port 128 nsew
flabel metal3 s -400 571592 60 571662 0 FreeSans 400 0 0 0 gpio_vtrip_sel[29]
port 304 nsew
flabel metal3 s -400 569752 60 569822 0 FreeSans 400 0 0 0 gpio_in_h[29]
port 744 nsew
flabel metal3 s -400 579596 60 579666 0 FreeSans 400 0 0 0 gpio_analog_en[29]
port 436 nsew
flabel metal3 s -400 578308 60 578378 0 FreeSans 400 0 0 0 gpio_analog_pol[29]
port 524 nsew
flabel metal3 s -400 578952 60 579022 0 FreeSans 400 0 0 0 gpio_dm0[29]
port 568 nsew
flabel metal3 s -400 577756 60 577826 0 FreeSans 400 0 0 0 gpio_inp_dis[29]
port 216 nsew
flabel metal3 s -400 580792 60 580862 0 FreeSans 400 0 0 0 gpio_dm1[29]
port 612 nsew
flabel metal3 s -400 582632 60 582702 0 FreeSans 400 0 0 0 gpio_slow_sel[29]
port 348 nsew
flabel metal3 s -400 584472 60 584542 0 FreeSans 400 0 0 0 gpio_in[29]
port 700 nsew
flabel metal3 s -400 622796 60 622866 0 FreeSans 400 0 0 0 gpio_analog_en[28]
port 437 nsew
flabel metal3 s -400 621508 60 621578 0 FreeSans 400 0 0 0 gpio_analog_pol[28]
port 525 nsew
flabel metal3 s -400 618472 60 618542 0 FreeSans 400 0 0 0 gpio_analog_sel[28]
port 481 nsew
flabel metal3 s -400 622152 60 622222 0 FreeSans 400 0 0 0 gpio_dm0[28]
port 569 nsew
flabel metal3 s -400 617828 60 617898 0 FreeSans 400 0 0 0 gpio_dm2[28]
port 657 nsew
flabel metal3 s -400 617184 60 617254 0 FreeSans 400 0 0 0 gpio_holdover[28]
port 393 nsew
flabel metal3 s -400 614148 60 614218 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[28]
port 261 nsew
flabel metal3 s -400 620956 60 621026 0 FreeSans 400 0 0 0 gpio_inp_dis[28]
port 217 nsew
flabel metal3 s -400 613504 60 613574 0 FreeSans 400 0 0 0 gpio_oeb[28]
port 173 nsew
flabel metal3 s -400 616632 60 616702 0 FreeSans 400 0 0 0 gpio_out[28]
port 129 nsew
flabel metal3 s -400 614792 60 614862 0 FreeSans 400 0 0 0 gpio_vtrip_sel[28]
port 305 nsew
flabel metal3 s -400 612952 60 613022 0 FreeSans 400 0 0 0 gpio_in_h[28]
port 745 nsew
flabel metal3 s -400 623992 60 624062 0 FreeSans 400 0 0 0 gpio_dm1[28]
port 613 nsew
flabel metal3 s -400 625832 60 625902 0 FreeSans 400 0 0 0 gpio_slow_sel[28]
port 349 nsew
flabel metal3 s -400 627672 60 627742 0 FreeSans 400 0 0 0 gpio_in[28]
port 701 nsew
flabel metal3 s -400 665996 60 666066 0 FreeSans 400 0 0 0 gpio_analog_en[27]
port 438 nsew
flabel metal3 s -400 664708 60 664778 0 FreeSans 400 0 0 0 gpio_analog_pol[27]
port 526 nsew
flabel metal3 s -400 661672 60 661742 0 FreeSans 400 0 0 0 gpio_analog_sel[27]
port 482 nsew
flabel metal3 s -400 665352 60 665422 0 FreeSans 400 0 0 0 gpio_dm0[27]
port 570 nsew
flabel metal3 s -400 661028 60 661098 0 FreeSans 400 0 0 0 gpio_dm2[27]
port 658 nsew
flabel metal3 s -400 660384 60 660454 0 FreeSans 400 0 0 0 gpio_holdover[27]
port 394 nsew
flabel metal3 s -400 657348 60 657418 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[27]
port 262 nsew
flabel metal3 s -400 664156 60 664226 0 FreeSans 400 0 0 0 gpio_inp_dis[27]
port 218 nsew
flabel metal3 s -400 656704 60 656774 0 FreeSans 400 0 0 0 gpio_oeb[27]
port 174 nsew
flabel metal3 s -400 659832 60 659902 0 FreeSans 400 0 0 0 gpio_out[27]
port 130 nsew
flabel metal3 s -400 657992 60 658062 0 FreeSans 400 0 0 0 gpio_vtrip_sel[27]
port 306 nsew
flabel metal3 s -400 656152 60 656222 0 FreeSans 400 0 0 0 gpio_in_h[27]
port 746 nsew
flabel metal3 s -400 667192 60 667262 0 FreeSans 400 0 0 0 gpio_dm1[27]
port 614 nsew
flabel metal3 s -400 669032 60 669102 0 FreeSans 400 0 0 0 gpio_slow_sel[27]
port 350 nsew
flabel metal3 s -400 670872 60 670942 0 FreeSans 400 0 0 0 gpio_in[27]
port 702 nsew
flabel metal3 -400 450940 60 455720 0 FreeSans 3200 90 0 0 vdda2
port 25 nsew
flabel metal3 -400 408814 60 413604 0 FreeSans 3200 90 0 0 vssd2
port 31 nsew
flabel metal3 -400 403862 60 408514 0 FreeSans 3200 90 0 0 vccd2
port 29 nsew
flabel metal3 -400 398762 60 403562 0 FreeSans 3200 90 0 0 vssd2
port 31 nsew
flabel metal3 -400 78140 60 82920 0 FreeSans 3200 90 0 0 vddio
port 18 nsew
flabel metal3 -400 36014 60 40804 0 FreeSans 3200 90 0 0 vccd
port 20 nsew
flabel metal3 -400 25962 60 30762 0 FreeSans 3200 90 0 0 vccd
port 20 nsew
flabel metal3 36806 -400 41586 60 0 FreeSans 3200 0 0 0 vssa
port 23 nsew
flabel metal3 199284 -400 203914 60 0 FreeSans 3200 0 0 0 vssd
port 21 nsew
flabel metal3 209164 -400 213964 60 0 FreeSans 3200 0 0 0 vssd
port 21 nsew
flabel metal3 527006 -400 531786 60 0 FreeSans 3200 0 0 0 vssio
port 19 nsew
flabel metal3 580806 -400 585586 60 0 FreeSans 3200 0 0 0 vdda
port 22 nsew
flabel metal3 633266 929006 633726 929068 0 FreeSans 400 0 0 0 gpio_loopback_zero[14]
port 803 nsew
flabel metal3 633266 839006 633726 839068 0 FreeSans 400 0 0 0 gpio_loopback_zero[13]
port 804 nsew
flabel metal3 633266 750006 633726 750068 0 FreeSans 400 0 0 0 gpio_loopback_zero[12]
port 805 nsew
flabel metal3 633266 705006 633726 705068 0 FreeSans 400 0 0 0 gpio_loopback_zero[11]
port 806 nsew
flabel metal3 633266 660006 633726 660068 0 FreeSans 400 0 0 0 gpio_loopback_zero[10]
port 807 nsew
flabel metal3 633266 615006 633726 615068 0 FreeSans 400 0 0 0 gpio_loopback_zero[9]
port 808 nsew
flabel metal3 633266 570006 633726 570068 0 FreeSans 400 0 0 0 gpio_loopback_zero[8]
port 809 nsew
flabel metal3 633266 525006 633726 525068 0 FreeSans 400 0 0 0 gpio_loopback_zero[7]
port 810 nsew
flabel metal3 633266 348006 633726 348068 0 FreeSans 400 0 0 0 gpio_loopback_zero[6]
port 811 nsew
flabel metal3 633266 303006 633726 303068 0 FreeSans 400 0 0 0 gpio_loopback_zero[5]
port 812 nsew
flabel metal3 633266 258006 633726 258068 0 FreeSans 400 0 0 0 gpio_loopback_zero[4]
port 813 nsew
flabel metal3 633266 213006 633726 213068 0 FreeSans 400 0 0 0 gpio_loopback_zero[3]
port 814 nsew
flabel metal3 633266 168006 633726 168068 0 FreeSans 400 0 0 0 gpio_loopback_zero[2]
port 815 nsew
flabel metal3 633266 123006 633726 123068 0 FreeSans 400 0 0 0 gpio_loopback_zero[1]
port 816 nsew
flabel metal3 633266 78006 633726 78068 0 FreeSans 400 0 0 0 gpio_loopback_zero[0]
port 817 nsew
flabel metal3 s 633266 60624 633726 60694 0 FreeSans 400 0 0 0 gpio_slow_sel[0]
port 377 nsew
flabel metal3 s 633266 58784 633726 58854 0 FreeSans 400 0 0 0 gpio_in[0]
port 729 nsew
flabel metal3 s 633266 62464 633726 62534 0 FreeSans 400 0 0 0 gpio_dm1[0]
port 641 nsew
flabel metal3 s 633266 63660 633726 63730 0 FreeSans 400 0 0 0 gpio_analog_en[0]
port 465 nsew
flabel metal3 s 633266 64948 633726 65018 0 FreeSans 400 0 0 0 gpio_analog_pol[0]
port 553 nsew
flabel metal3 s 633266 67984 633726 68054 0 FreeSans 400 0 0 0 gpio_analog_sel[0]
port 509 nsew
flabel metal3 s 633266 64304 633726 64374 0 FreeSans 400 0 0 0 gpio_dm0[0]
port 597 nsew
flabel metal3 s 633266 68628 633726 68698 0 FreeSans 400 0 0 0 gpio_dm2[0]
port 685 nsew
flabel metal3 s 633266 69272 633726 69342 0 FreeSans 400 0 0 0 gpio_holdover[0]
port 421 nsew
flabel metal3 s 633266 72308 633726 72378 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[0]
port 289 nsew
flabel metal3 s 633266 65500 633726 65570 0 FreeSans 400 0 0 0 gpio_inp_dis[0]
port 245 nsew
flabel metal3 s 633266 72952 633726 73022 0 FreeSans 400 0 0 0 gpio_oeb[0]
port 201 nsew
flabel metal3 s 633266 69824 633726 69894 0 FreeSans 400 0 0 0 gpio_out[0]
port 157 nsew
flabel metal3 s 633266 71664 633726 71734 0 FreeSans 400 0 0 0 gpio_vtrip_sel[0]
port 333 nsew
flabel metal3 633266 73504 633726 73574 0 FreeSans 400 0 0 0 gpio_in_h[0]
port 773 nsew
flabel metal3 s 633266 105824 633726 105894 0 FreeSans 400 0 0 0 gpio_slow_sel[1]
port 376 nsew
flabel metal3 s 633266 103984 633726 104054 0 FreeSans 400 0 0 0 gpio_in[1]
port 728 nsew
flabel metal3 s 633266 107664 633726 107734 0 FreeSans 400 0 0 0 gpio_dm1[1]
port 640 nsew
flabel metal3 s 633266 108860 633726 108930 0 FreeSans 400 0 0 0 gpio_analog_en[1]
port 464 nsew
flabel metal3 s 633266 110148 633726 110218 0 FreeSans 400 0 0 0 gpio_analog_pol[1]
port 552 nsew
flabel metal3 s 633266 113184 633726 113254 0 FreeSans 400 0 0 0 gpio_analog_sel[1]
port 508 nsew
flabel metal3 s 633266 109504 633726 109574 0 FreeSans 400 0 0 0 gpio_dm0[1]
port 596 nsew
flabel metal3 s 633266 113828 633726 113898 0 FreeSans 400 0 0 0 gpio_dm2[1]
port 684 nsew
flabel metal3 s 633266 114472 633726 114542 0 FreeSans 400 0 0 0 gpio_holdover[1]
port 420 nsew
flabel metal3 s 633266 117508 633726 117578 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[1]
port 288 nsew
flabel metal3 s 633266 110700 633726 110770 0 FreeSans 400 0 0 0 gpio_inp_dis[1]
port 244 nsew
flabel metal3 s 633266 118152 633726 118222 0 FreeSans 400 0 0 0 gpio_oeb[1]
port 200 nsew
flabel metal3 s 633266 115024 633726 115094 0 FreeSans 400 0 0 0 gpio_out[1]
port 156 nsew
flabel metal3 s 633266 116864 633726 116934 0 FreeSans 400 0 0 0 gpio_vtrip_sel[1]
port 332 nsew
flabel metal3 633266 118704 633726 118774 0 FreeSans 400 0 0 0 gpio_in_h[1]
port 772 nsew
flabel metal3 s 633266 150824 633726 150894 0 FreeSans 400 0 0 0 gpio_slow_sel[2]
port 375 nsew
flabel metal3 s 633266 148984 633726 149054 0 FreeSans 400 0 0 0 gpio_in[2]
port 727 nsew
flabel metal3 s 633266 152664 633726 152734 0 FreeSans 400 0 0 0 gpio_dm1[2]
port 639 nsew
flabel metal3 s 633266 153860 633726 153930 0 FreeSans 400 0 0 0 gpio_analog_en[2]
port 463 nsew
flabel metal3 s 633266 155148 633726 155218 0 FreeSans 400 0 0 0 gpio_analog_pol[2]
port 551 nsew
flabel metal3 s 633266 158184 633726 158254 0 FreeSans 400 0 0 0 gpio_analog_sel[2]
port 507 nsew
flabel metal3 s 633266 154504 633726 154574 0 FreeSans 400 0 0 0 gpio_dm0[2]
port 595 nsew
flabel metal3 s 633266 158828 633726 158898 0 FreeSans 400 0 0 0 gpio_dm2[2]
port 683 nsew
flabel metal3 s 633266 159472 633726 159542 0 FreeSans 400 0 0 0 gpio_holdover[2]
port 419 nsew
flabel metal3 s 633266 162508 633726 162578 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[2]
port 287 nsew
flabel metal3 s 633266 155700 633726 155770 0 FreeSans 400 0 0 0 gpio_inp_dis[2]
port 243 nsew
flabel metal3 s 633266 163152 633726 163222 0 FreeSans 400 0 0 0 gpio_oeb[2]
port 199 nsew
flabel metal3 s 633266 160024 633726 160094 0 FreeSans 400 0 0 0 gpio_out[2]
port 155 nsew
flabel metal3 s 633266 161864 633726 161934 0 FreeSans 400 0 0 0 gpio_vtrip_sel[2]
port 331 nsew
flabel metal3 633266 163704 633726 163774 0 FreeSans 400 0 0 0 gpio_in_h[2]
port 771 nsew
flabel metal3 s 633266 196024 633726 196094 0 FreeSans 400 0 0 0 gpio_slow_sel[3]
port 374 nsew
flabel metal3 s 633266 194184 633726 194254 0 FreeSans 400 0 0 0 gpio_in[3]
port 726 nsew
flabel metal3 s 633266 197864 633726 197934 0 FreeSans 400 0 0 0 gpio_dm1[3]
port 638 nsew
flabel metal3 s 633266 199060 633726 199130 0 FreeSans 400 0 0 0 gpio_analog_en[3]
port 462 nsew
flabel metal3 s 633266 200348 633726 200418 0 FreeSans 400 0 0 0 gpio_analog_pol[3]
port 550 nsew
flabel metal3 s 633266 203384 633726 203454 0 FreeSans 400 0 0 0 gpio_analog_sel[3]
port 506 nsew
flabel metal3 s 633266 204028 633726 204098 0 FreeSans 400 0 0 0 gpio_dm2[3]
port 682 nsew
flabel metal3 s 633266 199704 633726 199774 0 FreeSans 400 0 0 0 gpio_dm0[3]
port 594 nsew
flabel metal3 s 633266 204672 633726 204742 0 FreeSans 400 0 0 0 gpio_holdover[3]
port 418 nsew
flabel metal3 s 633266 207708 633726 207778 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[3]
port 286 nsew
flabel metal3 s 633266 200900 633726 200970 0 FreeSans 400 0 0 0 gpio_inp_dis[3]
port 242 nsew
flabel metal3 s 633266 208352 633726 208422 0 FreeSans 400 0 0 0 gpio_oeb[3]
port 198 nsew
flabel metal3 s 633266 205224 633726 205294 0 FreeSans 400 0 0 0 gpio_out[3]
port 154 nsew
flabel metal3 s 633266 207064 633726 207134 0 FreeSans 400 0 0 0 gpio_vtrip_sel[3]
port 330 nsew
flabel metal3 633266 208904 633726 208974 0 FreeSans 400 0 0 0 gpio_in_h[3]
port 770 nsew
flabel metal3 s 633266 241024 633726 241094 0 FreeSans 400 0 0 0 gpio_slow_sel[4]
port 373 nsew
flabel metal3 s 633266 239184 633726 239254 0 FreeSans 400 0 0 0 gpio_in[4]
port 725 nsew
flabel metal3 s 633266 242864 633726 242934 0 FreeSans 400 0 0 0 gpio_dm1[4]
port 637 nsew
flabel metal3 s 633266 244060 633726 244130 0 FreeSans 400 0 0 0 gpio_analog_en[4]
port 461 nsew
flabel metal3 s 633266 245348 633726 245418 0 FreeSans 400 0 0 0 gpio_analog_pol[4]
port 549 nsew
flabel metal3 s 633266 248384 633726 248454 0 FreeSans 400 0 0 0 gpio_analog_sel[4]
port 505 nsew
flabel metal3 s 633266 244704 633726 244774 0 FreeSans 400 0 0 0 gpio_dm0[4]
port 593 nsew
flabel metal3 s 633266 249028 633726 249098 0 FreeSans 400 0 0 0 gpio_dm2[4]
port 681 nsew
flabel metal3 s 633266 249672 633726 249742 0 FreeSans 400 0 0 0 gpio_holdover[4]
port 417 nsew
flabel metal3 s 633266 252708 633726 252778 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[4]
port 285 nsew
flabel metal3 s 633266 245900 633726 245970 0 FreeSans 400 0 0 0 gpio_inp_dis[4]
port 241 nsew
flabel metal3 s 633266 253352 633726 253422 0 FreeSans 400 0 0 0 gpio_oeb[4]
port 197 nsew
flabel metal3 s 633266 250224 633726 250294 0 FreeSans 400 0 0 0 gpio_out[4]
port 153 nsew
flabel metal3 s 633266 252064 633726 252134 0 FreeSans 400 0 0 0 gpio_vtrip_sel[4]
port 329 nsew
flabel metal3 633266 253904 633726 253974 0 FreeSans 400 0 0 0 gpio_in_h[4]
port 769 nsew
flabel metal3 s 633266 286024 633726 286094 0 FreeSans 400 0 0 0 gpio_slow_sel[5]
port 372 nsew
flabel metal3 s 633266 284184 633726 284254 0 FreeSans 400 0 0 0 gpio_in[5]
port 724 nsew
flabel metal3 s 633266 287864 633726 287934 0 FreeSans 400 0 0 0 gpio_dm1[5]
port 636 nsew
flabel metal3 s 633266 289060 633726 289130 0 FreeSans 400 0 0 0 gpio_analog_en[5]
port 460 nsew
flabel metal3 s 633266 290348 633726 290418 0 FreeSans 400 0 0 0 gpio_analog_pol[5]
port 548 nsew
flabel metal3 s 633266 293384 633726 293454 0 FreeSans 400 0 0 0 gpio_analog_sel[5]
port 504 nsew
flabel metal3 s 633266 289704 633726 289774 0 FreeSans 400 0 0 0 gpio_dm0[5]
port 592 nsew
flabel metal3 s 633266 294028 633726 294098 0 FreeSans 400 0 0 0 gpio_dm2[5]
port 680 nsew
flabel metal3 s 633266 294672 633726 294742 0 FreeSans 400 0 0 0 gpio_holdover[5]
port 416 nsew
flabel metal3 s 633266 297708 633726 297778 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[5]
port 284 nsew
flabel metal3 s 633266 290900 633726 290970 0 FreeSans 400 0 0 0 gpio_inp_dis[5]
port 240 nsew
flabel metal3 s 633266 298352 633726 298422 0 FreeSans 400 0 0 0 gpio_oeb[5]
port 196 nsew
flabel metal3 s 633266 295224 633726 295294 0 FreeSans 400 0 0 0 gpio_out[5]
port 152 nsew
flabel metal3 s 633266 297064 633726 297134 0 FreeSans 400 0 0 0 gpio_vtrip_sel[5]
port 328 nsew
flabel metal3 633266 298904 633726 298974 0 FreeSans 400 0 0 0 gpio_in_h[5]
port 768 nsew
flabel metal3 s 633266 331224 633726 331294 0 FreeSans 400 0 0 0 gpio_slow_sel[6]
port 371 nsew
flabel metal3 s 633266 329384 633726 329454 0 FreeSans 400 0 0 0 gpio_in[6]
port 723 nsew
flabel metal3 s 633266 333064 633726 333134 0 FreeSans 400 0 0 0 gpio_dm1[6]
port 635 nsew
flabel metal3 s 633266 334260 633726 334330 0 FreeSans 400 0 0 0 gpio_analog_en[6]
port 459 nsew
flabel metal3 s 633266 335548 633726 335618 0 FreeSans 400 0 0 0 gpio_analog_pol[6]
port 547 nsew
flabel metal3 s 633266 338584 633726 338654 0 FreeSans 400 0 0 0 gpio_analog_sel[6]
port 503 nsew
flabel metal3 s 633266 334904 633726 334974 0 FreeSans 400 0 0 0 gpio_dm0[6]
port 591 nsew
flabel metal3 s 633266 339228 633726 339298 0 FreeSans 400 0 0 0 gpio_dm2[6]
port 679 nsew
flabel metal3 s 633266 339872 633726 339942 0 FreeSans 400 0 0 0 gpio_holdover[6]
port 415 nsew
flabel metal3 s 633266 342908 633726 342978 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[6]
port 283 nsew
flabel metal3 s 633266 336100 633726 336170 0 FreeSans 400 0 0 0 gpio_inp_dis[6]
port 239 nsew
flabel metal3 s 633266 343552 633726 343622 0 FreeSans 400 0 0 0 gpio_oeb[6]
port 195 nsew
flabel metal3 s 633266 340424 633726 340494 0 FreeSans 400 0 0 0 gpio_out[6]
port 151 nsew
flabel metal3 s 633266 342264 633726 342334 0 FreeSans 400 0 0 0 gpio_vtrip_sel[6]
port 327 nsew
flabel metal3 633266 344104 633726 344174 0 FreeSans 400 0 0 0 gpio_in_h[6]
port 767 nsew
flabel metal3 s 633266 508424 633726 508494 0 FreeSans 400 0 0 0 gpio_slow_sel[7]
port 370 nsew
flabel metal3 s 633266 506584 633726 506654 0 FreeSans 400 0 0 0 gpio_in[7]
port 722 nsew
flabel metal3 s 633266 510264 633726 510334 0 FreeSans 400 0 0 0 gpio_dm1[7]
port 634 nsew
flabel metal3 s 633266 511460 633726 511530 0 FreeSans 400 0 0 0 gpio_analog_en[7]
port 458 nsew
flabel metal3 s 633266 512748 633726 512818 0 FreeSans 400 0 0 0 gpio_analog_pol[7]
port 546 nsew
flabel metal3 s 633266 515784 633726 515854 0 FreeSans 400 0 0 0 gpio_analog_sel[7]
port 502 nsew
flabel metal3 s 633266 512104 633726 512174 0 FreeSans 400 0 0 0 gpio_dm0[7]
port 590 nsew
flabel metal3 s 633266 516428 633726 516498 0 FreeSans 400 0 0 0 gpio_dm2[7]
port 678 nsew
flabel metal3 s 633266 517072 633726 517142 0 FreeSans 400 0 0 0 gpio_holdover[7]
port 414 nsew
flabel metal3 s 633266 520108 633726 520178 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[7]
port 282 nsew
flabel metal3 s 633266 513300 633726 513370 0 FreeSans 400 0 0 0 gpio_inp_dis[7]
port 238 nsew
flabel metal3 s 633266 520752 633726 520822 0 FreeSans 400 0 0 0 gpio_oeb[7]
port 194 nsew
flabel metal3 s 633266 517624 633726 517694 0 FreeSans 400 0 0 0 gpio_out[7]
port 150 nsew
flabel metal3 s 633266 519464 633726 519534 0 FreeSans 400 0 0 0 gpio_vtrip_sel[7]
port 326 nsew
flabel metal3 s 633266 521304 633726 521374 0 FreeSans 400 0 0 0 gpio_in_h[7]
port 766 nsew
flabel metal3 s 633266 553624 633726 553694 0 FreeSans 400 0 0 0 gpio_slow_sel[8]
port 369 nsew
flabel metal3 s 633266 551784 633726 551854 0 FreeSans 400 0 0 0 gpio_in[8]
port 721 nsew
flabel metal3 s 633266 555464 633726 555534 0 FreeSans 400 0 0 0 gpio_dm1[8]
port 633 nsew
flabel metal3 s 633266 556660 633726 556730 0 FreeSans 400 0 0 0 gpio_analog_en[8]
port 457 nsew
flabel metal3 s 633266 557948 633726 558018 0 FreeSans 400 0 0 0 gpio_analog_pol[8]
port 545 nsew
flabel metal3 s 633266 560984 633726 561054 0 FreeSans 400 0 0 0 gpio_analog_sel[8]
port 501 nsew
flabel metal3 s 633266 557304 633726 557374 0 FreeSans 400 0 0 0 gpio_dm0[8]
port 589 nsew
flabel metal3 s 633266 561628 633726 561698 0 FreeSans 400 0 0 0 gpio_dm2[8]
port 677 nsew
flabel metal3 s 633266 562272 633726 562342 0 FreeSans 400 0 0 0 gpio_holdover[8]
port 413 nsew
flabel metal3 s 633266 565308 633726 565378 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[8]
port 281 nsew
flabel metal3 s 633266 558500 633726 558570 0 FreeSans 400 0 0 0 gpio_inp_dis[8]
port 237 nsew
flabel metal3 s 633266 565952 633726 566022 0 FreeSans 400 0 0 0 gpio_oeb[8]
port 193 nsew
flabel metal3 s 633266 562824 633726 562894 0 FreeSans 400 0 0 0 gpio_out[8]
port 149 nsew
flabel metal3 s 633266 564664 633726 564734 0 FreeSans 400 0 0 0 gpio_vtrip_sel[8]
port 325 nsew
flabel metal3 s 633266 566504 633726 566574 0 FreeSans 400 0 0 0 gpio_in_h[8]
port 765 nsew
flabel metal3 s 633266 598624 633726 598694 0 FreeSans 400 0 0 0 gpio_slow_sel[9]
port 368 nsew
flabel metal3 s 633266 596784 633726 596854 0 FreeSans 400 0 0 0 gpio_in[9]
port 720 nsew
flabel metal3 s 633266 600464 633726 600534 0 FreeSans 400 0 0 0 gpio_dm1[9]
port 632 nsew
flabel metal3 s 633266 601660 633726 601730 0 FreeSans 400 0 0 0 gpio_analog_en[9]
port 456 nsew
flabel metal3 s 633266 602948 633726 603018 0 FreeSans 400 0 0 0 gpio_analog_pol[9]
port 544 nsew
flabel metal3 s 633266 605984 633726 606054 0 FreeSans 400 0 0 0 gpio_analog_sel[9]
port 500 nsew
flabel metal3 s 633266 602304 633726 602374 0 FreeSans 400 0 0 0 gpio_dm0[9]
port 588 nsew
flabel metal3 s 633266 606628 633726 606698 0 FreeSans 400 0 0 0 gpio_dm2[9]
port 676 nsew
flabel metal3 s 633266 607272 633726 607342 0 FreeSans 400 0 0 0 gpio_holdover[9]
port 412 nsew
flabel metal3 s 633266 610308 633726 610378 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[9]
port 280 nsew
flabel metal3 s 633266 603500 633726 603570 0 FreeSans 400 0 0 0 gpio_inp_dis[9]
port 236 nsew
flabel metal3 s 633266 610952 633726 611022 0 FreeSans 400 0 0 0 gpio_oeb[9]
port 192 nsew
flabel metal3 s 633266 607824 633726 607894 0 FreeSans 400 0 0 0 gpio_out[9]
port 148 nsew
flabel metal3 s 633266 609664 633726 609734 0 FreeSans 400 0 0 0 gpio_vtrip_sel[9]
port 324 nsew
flabel metal3 s 633266 611504 633726 611574 0 FreeSans 400 0 0 0 gpio_in_h[9]
port 764 nsew
flabel metal3 s 633266 643824 633726 643894 0 FreeSans 400 0 0 0 gpio_slow_sel[10]
port 367 nsew
flabel metal3 s 633266 641984 633726 642054 0 FreeSans 400 0 0 0 gpio_in[10]
port 719 nsew
flabel metal3 s 633266 645664 633726 645734 0 FreeSans 400 0 0 0 gpio_dm1[10]
port 631 nsew
flabel metal3 s 633266 646860 633726 646930 0 FreeSans 400 0 0 0 gpio_analog_en[10]
port 455 nsew
flabel metal3 s 633266 648148 633726 648218 0 FreeSans 400 0 0 0 gpio_analog_pol[10]
port 543 nsew
flabel metal3 s 633266 651184 633726 651254 0 FreeSans 400 0 0 0 gpio_analog_sel[10]
port 499 nsew
flabel metal3 s 633266 647504 633726 647574 0 FreeSans 400 0 0 0 gpio_dm0[10]
port 587 nsew
flabel metal3 s 633266 651828 633726 651898 0 FreeSans 400 0 0 0 gpio_dm2[10]
port 675 nsew
flabel metal3 s 633266 652472 633726 652542 0 FreeSans 400 0 0 0 gpio_holdover[10]
port 411 nsew
flabel metal3 s 633266 655508 633726 655578 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[10]
port 279 nsew
flabel metal3 s 633266 648700 633726 648770 0 FreeSans 400 0 0 0 gpio_inp_dis[10]
port 235 nsew
flabel metal3 s 633266 656152 633726 656222 0 FreeSans 400 0 0 0 gpio_oeb[10]
port 191 nsew
flabel metal3 s 633266 653024 633726 653094 0 FreeSans 400 0 0 0 gpio_out[10]
port 147 nsew
flabel metal3 s 633266 654864 633726 654934 0 FreeSans 400 0 0 0 gpio_vtrip_sel[10]
port 323 nsew
flabel metal3 s 633266 656704 633726 656774 0 FreeSans 400 0 0 0 gpio_in_h[10]
port 763 nsew
flabel metal3 s 633266 688824 633726 688894 0 FreeSans 400 0 0 0 gpio_slow_sel[11]
port 366 nsew
flabel metal3 s 633266 686984 633726 687054 0 FreeSans 400 0 0 0 gpio_in[11]
port 718 nsew
flabel metal3 s 633266 690664 633726 690734 0 FreeSans 400 0 0 0 gpio_dm1[11]
port 630 nsew
flabel metal3 s 633266 697472 633726 697542 0 FreeSans 400 0 0 0 gpio_holdover[11]
port 410 nsew
flabel metal3 s 633266 700508 633726 700578 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[11]
port 278 nsew
flabel metal3 s 633266 693700 633726 693770 0 FreeSans 400 0 0 0 gpio_inp_dis[11]
port 234 nsew
flabel metal3 s 633266 701152 633726 701222 0 FreeSans 400 0 0 0 gpio_oeb[11]
port 190 nsew
flabel metal3 s 633266 698024 633726 698094 0 FreeSans 400 0 0 0 gpio_out[11]
port 146 nsew
flabel metal3 s 633266 699864 633726 699934 0 FreeSans 400 0 0 0 gpio_vtrip_sel[11]
port 322 nsew
flabel metal3 s 633266 691860 633726 691930 0 FreeSans 400 0 0 0 gpio_analog_en[11]
port 454 nsew
flabel metal3 s 633266 693148 633726 693218 0 FreeSans 400 0 0 0 gpio_analog_pol[11]
port 542 nsew
flabel metal3 s 633266 696184 633726 696254 0 FreeSans 400 0 0 0 gpio_analog_sel[11]
port 498 nsew
flabel metal3 s 633266 692504 633726 692574 0 FreeSans 400 0 0 0 gpio_dm0[11]
port 586 nsew
flabel metal3 s 633266 696828 633726 696898 0 FreeSans 400 0 0 0 gpio_dm2[11]
port 674 nsew
flabel metal3 s 633266 701704 633726 701774 0 FreeSans 400 0 0 0 gpio_in_h[11]
port 762 nsew
flabel metal3 s 633266 733824 633726 733894 0 FreeSans 400 0 0 0 gpio_slow_sel[12]
port 365 nsew
flabel metal3 s 633266 731984 633726 732054 0 FreeSans 400 0 0 0 gpio_in[12]
port 717 nsew
flabel metal3 s 633266 735664 633726 735734 0 FreeSans 400 0 0 0 gpio_dm1[12]
port 629 nsew
flabel metal3 s 633266 736860 633726 736930 0 FreeSans 400 0 0 0 gpio_analog_en[12]
port 453 nsew
flabel metal3 s 633266 738148 633726 738218 0 FreeSans 400 0 0 0 gpio_analog_pol[12]
port 541 nsew
flabel metal3 s 633266 741184 633726 741254 0 FreeSans 400 0 0 0 gpio_analog_sel[12]
port 497 nsew
flabel metal3 s 633266 737504 633726 737574 0 FreeSans 400 0 0 0 gpio_dm0[12]
port 585 nsew
flabel metal3 s 633266 741828 633726 741898 0 FreeSans 400 0 0 0 gpio_dm2[12]
port 673 nsew
flabel metal3 s 633266 742472 633726 742542 0 FreeSans 400 0 0 0 gpio_holdover[12]
port 409 nsew
flabel metal3 s 633266 745508 633726 745578 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[12]
port 277 nsew
flabel metal3 s 633266 738700 633726 738770 0 FreeSans 400 0 0 0 gpio_inp_dis[12]
port 233 nsew
flabel metal3 s 633266 746152 633726 746222 0 FreeSans 400 0 0 0 gpio_oeb[12]
port 189 nsew
flabel metal3 s 633266 743024 633726 743094 0 FreeSans 400 0 0 0 gpio_out[12]
port 145 nsew
flabel metal3 s 633266 744864 633726 744934 0 FreeSans 400 0 0 0 gpio_vtrip_sel[12]
port 321 nsew
flabel metal3 s 633266 746704 633726 746774 0 FreeSans 400 0 0 0 gpio_in_h[12]
port 761 nsew
flabel metal3 s 633266 823024 633726 823094 0 FreeSans 400 0 0 0 gpio_slow_sel[13]
port 364 nsew
flabel metal3 s 633266 821184 633726 821254 0 FreeSans 400 0 0 0 gpio_in[13]
port 716 nsew
flabel metal3 s 633266 824864 633726 824934 0 FreeSans 400 0 0 0 gpio_dm1[13]
port 628 nsew
flabel metal3 s 633266 826060 633726 826130 0 FreeSans 400 0 0 0 gpio_analog_en[13]
port 452 nsew
flabel metal3 s 633266 827348 633726 827418 0 FreeSans 400 0 0 0 gpio_analog_pol[13]
port 540 nsew
flabel metal3 s 633266 830384 633726 830454 0 FreeSans 400 0 0 0 gpio_analog_sel[13]
port 496 nsew
flabel metal3 s 633266 826704 633726 826774 0 FreeSans 400 0 0 0 gpio_dm0[13]
port 584 nsew
flabel metal3 s 633266 831028 633726 831098 0 FreeSans 400 0 0 0 gpio_dm2[13]
port 672 nsew
flabel metal3 s 633266 831672 633726 831742 0 FreeSans 400 0 0 0 gpio_holdover[13]
port 408 nsew
flabel metal3 s 633266 834708 633726 834778 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[13]
port 276 nsew
flabel metal3 s 633266 827900 633726 827970 0 FreeSans 400 0 0 0 gpio_inp_dis[13]
port 232 nsew
flabel metal3 s 633266 835352 633726 835422 0 FreeSans 400 0 0 0 gpio_oeb[13]
port 188 nsew
flabel metal3 s 633266 832224 633726 832294 0 FreeSans 400 0 0 0 gpio_out[13]
port 144 nsew
flabel metal3 s 633266 834064 633726 834134 0 FreeSans 400 0 0 0 gpio_vtrip_sel[13]
port 320 nsew
flabel metal3 s 633266 835904 633726 835974 0 FreeSans 400 0 0 0 gpio_in_h[13]
port 760 nsew
flabel metal3 s 633266 912224 633726 912294 0 FreeSans 400 0 0 0 gpio_slow_sel[14]
port 363 nsew
flabel metal3 s 633266 910384 633726 910454 0 FreeSans 400 0 0 0 gpio_in[14]
port 715 nsew
flabel metal3 s 633266 914064 633726 914134 0 FreeSans 400 0 0 0 gpio_dm1[14]
port 627 nsew
flabel metal3 s 633266 915260 633726 915330 0 FreeSans 400 0 0 0 gpio_analog_en[14]
port 451 nsew
flabel metal3 s 633266 916548 633726 916618 0 FreeSans 400 0 0 0 gpio_analog_pol[14]
port 539 nsew
flabel metal3 s 633266 919584 633726 919654 0 FreeSans 400 0 0 0 gpio_analog_sel[14]
port 495 nsew
flabel metal3 s 633266 915904 633726 915974 0 FreeSans 400 0 0 0 gpio_dm0[14]
port 583 nsew
flabel metal3 s 633266 920228 633726 920298 0 FreeSans 400 0 0 0 gpio_dm2[14]
port 671 nsew
flabel metal3 s 633266 920872 633726 920942 0 FreeSans 400 0 0 0 gpio_holdover[14]
port 407 nsew
flabel metal3 s 633266 923908 633726 923978 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[14]
port 275 nsew
flabel metal3 s 633266 917100 633726 917170 0 FreeSans 400 0 0 0 gpio_inp_dis[14]
port 231 nsew
flabel metal3 s 633266 924552 633726 924622 0 FreeSans 400 0 0 0 gpio_oeb[14]
port 187 nsew
flabel metal3 s 633266 921424 633726 921494 0 FreeSans 400 0 0 0 gpio_out[14]
port 143 nsew
flabel metal3 s 633266 923264 633726 923334 0 FreeSans 400 0 0 0 gpio_vtrip_sel[14]
port 319 nsew
flabel metal3 s 633266 925104 633726 925174 0 FreeSans 400 0 0 0 gpio_in_h[14]
port 759 nsew
flabel metal3 s -400 927072 60 927142 0 FreeSans 400 0 0 0 gpio_in[24]
port 705 nsew
flabel metal3 s -400 925232 60 925302 0 FreeSans 400 0 0 0 gpio_slow_sel[24]
port 353 nsew
flabel metal3 s -400 923392 60 923462 0 FreeSans 400 0 0 0 gpio_dm1[24]
port 617 nsew
flabel metal3 s -400 922196 60 922266 0 FreeSans 400 0 0 0 gpio_analog_en[24]
port 441 nsew
flabel metal3 s -400 921552 60 921622 0 FreeSans 400 0 0 0 gpio_dm0[24]
port 573 nsew
flabel metal3 s -400 920908 60 920978 0 FreeSans 400 0 0 0 gpio_analog_pol[24]
port 529 nsew
flabel metal3 s -400 920356 60 920426 0 FreeSans 400 0 0 0 gpio_inp_dis[24]
port 221 nsew
flabel metal3 s -400 917872 60 917942 0 FreeSans 400 0 0 0 gpio_analog_sel[24]
port 485 nsew
flabel metal3 s -400 917228 60 917298 0 FreeSans 400 0 0 0 gpio_dm2[24]
port 661 nsew
flabel metal3 s -400 916584 60 916654 0 FreeSans 400 0 0 0 gpio_holdover[24]
port 397 nsew
flabel metal3 s -400 916032 60 916102 0 FreeSans 400 0 0 0 gpio_out[24]
port 133 nsew
flabel metal3 s -400 914192 60 914262 0 FreeSans 400 0 0 0 gpio_vtrip_sel[24]
port 309 nsew
flabel metal3 s -400 913548 60 913618 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[24]
port 265 nsew
flabel metal3 s -400 912904 60 912974 0 FreeSans 400 0 0 0 gpio_oeb[24]
port 177 nsew
flabel metal3 s -400 912352 60 912422 0 FreeSans 400 0 0 0 gpio_in_h[24]
port 749 nsew
flabel metal3 s -400 924560 60 924688 0 FreeSans 400 0 0 0 analog_io[24]
port 881 nsew
flabel metal3 s -400 922677 60 922891 0 FreeSans 400 0 0 0 analog_noesd_io[24]
port 925 nsew
flabel metal2 27498 953270 27558 953726 0 FreeSans 400 90 0 0 gpio_loopback_zero[23]
port 794 nsew
flabel metal2 78698 953270 78758 953726 0 FreeSans 400 90 0 0 gpio_loopback_zero[22]
port 795 nsew
flabel metal2 129898 953270 129958 953726 0 FreeSans 400 90 0 0 gpio_loopback_zero[21]
port 796 nsew
flabel metal2 181098 953270 181158 953726 0 FreeSans 400 90 0 0 gpio_loopback_zero[20]
port 797 nsew
flabel metal2 232298 953270 232358 953726 0 FreeSans 400 90 0 0 gpio_loopback_zero[19]
port 798 nsew
flabel metal2 336698 953270 336758 953726 0 FreeSans 400 90 0 0 gpio_loopback_zero[18]
port 799 nsew
flabel metal2 425698 953270 425758 953726 0 FreeSans 400 90 0 0 gpio_loopback_zero[17]
port 800 nsew
flabel metal2 476898 953270 476958 953726 0 FreeSans 400 90 0 0 gpio_loopback_zero[16]
port 801 nsew
flabel metal2 576298 953270 576358 953726 0 FreeSans 400 90 0 0 gpio_loopback_zero[15]
port 802 nsew
<< properties >>
string FIXED_BBOX 0 0 633326 953326
<< end >>
