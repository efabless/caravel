VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO simple_por
  CLASS BLOCK ;
  FOREIGN simple_por ;
  ORIGIN 0.000 0.000 ;
  SIZE 56.720 BY 41.690 ;
  PIN vdd3v3
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.350 36.720 34.910 41.690 ;
        RECT 37.005 33.995 54.465 36.505 ;
        RECT 37.005 33.905 38.675 33.995 ;
        RECT 41.220 33.905 54.465 33.995 ;
      LAYER li1 ;
        RECT 0.205 41.300 0.915 41.440 ;
        RECT 34.455 41.300 35.670 41.430 ;
        RECT 0.205 41.130 35.670 41.300 ;
        RECT 0.205 37.280 0.915 41.130 ;
        RECT 3.170 37.280 3.340 41.130 ;
        RECT 3.840 38.185 4.010 40.225 ;
        RECT 6.020 38.185 6.190 40.225 ;
        RECT 8.200 38.185 8.370 40.225 ;
        RECT 10.380 38.185 10.550 40.225 ;
        RECT 12.560 38.185 12.730 40.225 ;
        RECT 13.230 37.280 13.400 41.130 ;
        RECT 13.900 38.185 14.070 40.225 ;
        RECT 15.660 37.280 15.830 41.130 ;
        RECT 18.090 37.280 18.260 41.130 ;
        RECT 20.520 37.280 20.690 41.130 ;
        RECT 21.190 38.185 21.360 40.225 ;
        RECT 23.370 38.185 23.540 40.225 ;
        RECT 25.550 38.185 25.720 40.225 ;
        RECT 27.730 38.185 27.900 40.225 ;
        RECT 29.490 37.280 29.660 41.130 ;
        RECT 30.160 38.185 30.330 40.225 ;
        RECT 31.920 37.280 32.090 41.130 ;
        RECT 34.350 37.280 35.670 41.130 ;
        RECT 0.205 36.610 35.670 37.280 ;
        RECT 0.205 36.525 54.145 36.610 ;
        RECT 15.215 36.005 54.145 36.525 ;
        RECT 15.215 35.025 35.670 36.005 ;
        RECT 40.465 35.425 41.905 35.755 ;
        RECT 40.570 34.340 41.905 35.425 ;
        RECT 43.230 35.645 52.120 35.815 ;
        RECT 43.230 34.465 44.480 35.645 ;
        RECT 45.380 34.405 46.050 35.645 ;
        RECT 46.720 34.405 47.610 35.645 ;
        RECT 48.280 34.405 49.170 35.645 ;
        RECT 49.840 34.405 50.730 35.645 ;
        RECT 51.520 35.495 52.120 35.645 ;
        RECT 51.750 34.405 52.120 35.495 ;
        RECT 51.010 27.990 51.700 30.150 ;
      LAYER mcon ;
        RECT 0.285 40.950 0.845 41.375 ;
        RECT 1.135 41.130 2.945 41.300 ;
        RECT 3.835 41.130 12.735 41.300 ;
        RECT 13.625 41.130 15.435 41.300 ;
        RECT 16.055 41.130 17.865 41.300 ;
        RECT 18.485 41.130 20.295 41.300 ;
        RECT 21.130 41.130 29.050 41.300 ;
        RECT 29.885 41.130 31.695 41.300 ;
        RECT 32.315 41.130 34.125 41.300 ;
        RECT 3.170 39.205 3.340 41.130 ;
        RECT 3.840 39.310 4.010 40.060 ;
        RECT 6.020 39.310 6.190 40.060 ;
        RECT 8.200 39.310 8.370 40.060 ;
        RECT 10.380 39.310 10.550 40.060 ;
        RECT 12.560 39.310 12.730 40.060 ;
        RECT 13.230 39.205 13.400 41.130 ;
        RECT 13.900 38.265 14.070 40.145 ;
        RECT 20.520 39.395 20.690 41.130 ;
        RECT 21.190 39.310 21.360 40.060 ;
        RECT 23.370 39.310 23.540 40.060 ;
        RECT 25.550 39.310 25.720 40.060 ;
        RECT 27.730 39.310 27.900 40.060 ;
        RECT 29.490 39.395 29.660 41.130 ;
        RECT 30.160 38.265 30.330 40.145 ;
        RECT 34.680 40.560 35.585 41.365 ;
        RECT 34.635 35.110 35.550 37.175 ;
        RECT 37.490 36.005 37.660 36.175 ;
        RECT 37.970 36.005 38.140 36.175 ;
        RECT 38.450 36.005 38.620 36.175 ;
        RECT 38.930 36.005 39.100 36.175 ;
        RECT 39.410 36.005 39.580 36.175 ;
        RECT 39.890 36.005 40.060 36.175 ;
        RECT 40.370 36.005 40.540 36.175 ;
        RECT 40.850 36.005 41.020 36.175 ;
        RECT 41.330 36.005 41.500 36.175 ;
        RECT 41.810 36.005 41.980 36.175 ;
        RECT 42.290 36.005 42.460 36.175 ;
        RECT 42.770 36.005 42.940 36.175 ;
        RECT 43.250 36.005 43.420 36.175 ;
        RECT 43.730 36.005 43.900 36.175 ;
        RECT 44.210 36.005 44.380 36.175 ;
        RECT 44.690 36.005 44.860 36.175 ;
        RECT 45.170 36.005 45.340 36.175 ;
        RECT 45.650 36.005 45.820 36.175 ;
        RECT 46.130 36.005 46.300 36.175 ;
        RECT 46.610 36.005 46.780 36.175 ;
        RECT 47.090 36.005 47.260 36.175 ;
        RECT 47.570 36.005 47.740 36.175 ;
        RECT 48.050 36.005 48.220 36.175 ;
        RECT 48.530 36.005 48.700 36.175 ;
        RECT 49.010 36.005 49.180 36.175 ;
        RECT 49.490 36.005 49.660 36.175 ;
        RECT 49.970 36.005 50.140 36.175 ;
        RECT 50.450 36.005 50.620 36.175 ;
        RECT 50.930 36.005 51.100 36.175 ;
        RECT 51.410 36.005 51.580 36.175 ;
        RECT 51.890 36.005 52.060 36.175 ;
        RECT 52.370 36.005 52.540 36.175 ;
        RECT 52.850 36.005 53.020 36.175 ;
        RECT 53.330 36.005 53.500 36.175 ;
        RECT 53.810 36.005 53.980 36.175 ;
        RECT 40.560 35.495 40.730 35.665 ;
        RECT 40.920 35.495 41.090 35.665 ;
        RECT 41.280 35.495 41.450 35.665 ;
        RECT 41.640 35.495 41.810 35.665 ;
        RECT 43.230 35.495 43.400 35.665 ;
        RECT 43.590 35.495 43.760 35.665 ;
        RECT 43.950 35.495 44.120 35.665 ;
        RECT 44.310 35.495 44.480 35.665 ;
        RECT 45.385 35.495 45.555 35.665 ;
        RECT 45.745 35.495 45.915 35.665 ;
        RECT 46.720 35.495 46.890 35.665 ;
        RECT 47.080 35.495 47.250 35.665 ;
        RECT 47.440 35.495 47.610 35.665 ;
        RECT 48.280 35.495 48.450 35.665 ;
        RECT 48.640 35.495 48.810 35.665 ;
        RECT 49.000 35.495 49.170 35.665 ;
        RECT 49.845 35.495 50.015 35.665 ;
        RECT 50.560 35.495 50.730 35.665 ;
        RECT 51.880 35.495 52.050 35.665 ;
      LAYER met1 ;
        RECT 0.200 41.045 35.665 41.430 ;
        RECT 0.200 40.895 35.670 41.045 ;
        RECT 3.140 40.140 3.370 40.895 ;
        RECT 13.200 40.140 13.430 40.895 ;
        RECT 13.870 40.140 14.100 40.205 ;
        RECT 20.490 40.165 20.720 40.895 ;
        RECT 29.460 40.165 29.690 40.895 ;
        RECT 30.130 40.165 30.360 40.205 ;
        RECT 3.135 39.460 14.105 40.140 ;
        RECT 3.140 39.145 3.370 39.460 ;
        RECT 3.810 39.250 4.040 39.460 ;
        RECT 5.990 39.250 6.220 39.460 ;
        RECT 8.170 39.250 8.400 39.460 ;
        RECT 10.350 39.250 10.580 39.460 ;
        RECT 12.530 39.250 12.760 39.460 ;
        RECT 13.200 39.145 13.430 39.460 ;
        RECT 13.870 38.205 14.100 39.460 ;
        RECT 20.490 39.360 30.360 40.165 ;
        RECT 20.490 39.335 20.720 39.360 ;
        RECT 21.160 39.250 21.390 39.360 ;
        RECT 23.340 39.250 23.570 39.360 ;
        RECT 25.520 39.250 25.750 39.360 ;
        RECT 27.700 39.250 27.930 39.360 ;
        RECT 29.460 39.335 29.690 39.360 ;
        RECT 30.130 38.205 30.360 39.360 ;
        RECT 34.550 36.620 35.670 40.895 ;
        RECT 34.550 35.470 54.160 36.620 ;
        RECT 34.550 34.970 35.670 35.470 ;
        RECT 37.335 35.465 54.160 35.470 ;
        RECT 51.105 30.880 53.580 31.350 ;
        RECT 51.105 30.225 51.575 30.880 ;
        RECT 50.935 27.910 51.765 30.225 ;
      LAYER via ;
        RECT 0.300 41.005 3.120 41.345 ;
        RECT 5.130 40.965 35.465 41.300 ;
        RECT 35.855 35.620 41.600 36.495 ;
        RECT 43.010 35.620 53.750 36.495 ;
        RECT 51.165 30.935 53.500 31.300 ;
      LAYER met2 ;
        RECT 4.925 41.430 35.660 41.435 ;
        RECT 0.190 40.935 35.660 41.430 ;
        RECT 0.190 40.305 3.270 40.935 ;
        RECT 4.330 40.300 35.660 40.935 ;
        RECT 35.705 35.470 41.775 36.620 ;
        RECT 42.835 35.470 53.990 36.620 ;
        RECT 51.105 31.350 52.155 35.470 ;
        RECT 51.105 30.880 53.580 31.350 ;
      LAYER via2 ;
        RECT 0.385 40.520 3.170 41.305 ;
        RECT 4.430 40.520 35.455 41.305 ;
      LAYER met3 ;
        RECT 0.190 39.825 35.630 41.415 ;
      LAYER via3 ;
        RECT 0.365 40.000 35.365 41.220 ;
      LAYER met4 ;
        RECT 0.190 39.825 35.630 41.415 ;
    END
  END vdd3v3
  PIN vdd1v8
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 37.055 39.075 54.515 41.675 ;
      LAYER li1 ;
        RECT 37.385 41.175 54.185 41.345 ;
        RECT 38.000 40.815 46.890 40.985 ;
        RECT 38.000 39.635 39.250 40.815 ;
        RECT 40.150 39.575 40.820 40.815 ;
        RECT 41.490 39.575 42.380 40.815 ;
        RECT 43.050 39.575 43.940 40.815 ;
        RECT 44.610 39.575 45.500 40.815 ;
        RECT 46.290 40.665 46.890 40.815 ;
        RECT 46.520 39.575 46.890 40.665 ;
        RECT 47.080 40.815 54.010 40.985 ;
        RECT 47.080 39.635 47.970 40.815 ;
        RECT 48.760 39.575 49.650 40.815 ;
        RECT 50.320 39.575 51.210 40.815 ;
        RECT 51.880 39.575 52.770 40.815 ;
        RECT 53.440 39.575 54.010 40.815 ;
      LAYER mcon ;
        RECT 37.540 41.175 37.710 41.345 ;
        RECT 38.020 41.175 38.190 41.345 ;
        RECT 38.500 41.175 38.670 41.345 ;
        RECT 38.980 41.175 39.150 41.345 ;
        RECT 39.460 41.175 39.630 41.345 ;
        RECT 39.940 41.175 40.110 41.345 ;
        RECT 40.420 41.175 40.590 41.345 ;
        RECT 40.900 41.175 41.070 41.345 ;
        RECT 41.380 41.175 41.550 41.345 ;
        RECT 41.860 41.175 42.030 41.345 ;
        RECT 42.340 41.175 42.510 41.345 ;
        RECT 42.820 41.175 42.990 41.345 ;
        RECT 43.300 41.175 43.470 41.345 ;
        RECT 43.780 41.175 43.950 41.345 ;
        RECT 44.260 41.175 44.430 41.345 ;
        RECT 44.740 41.175 44.910 41.345 ;
        RECT 45.220 41.175 45.390 41.345 ;
        RECT 45.700 41.175 45.870 41.345 ;
        RECT 46.180 41.175 46.350 41.345 ;
        RECT 46.660 41.175 46.830 41.345 ;
        RECT 47.140 41.175 47.310 41.345 ;
        RECT 47.620 41.175 47.790 41.345 ;
        RECT 48.100 41.175 48.270 41.345 ;
        RECT 48.580 41.175 48.750 41.345 ;
        RECT 49.060 41.175 49.230 41.345 ;
        RECT 49.540 41.175 49.710 41.345 ;
        RECT 50.020 41.175 50.190 41.345 ;
        RECT 50.500 41.175 50.670 41.345 ;
        RECT 50.980 41.175 51.150 41.345 ;
        RECT 51.460 41.175 51.630 41.345 ;
        RECT 51.940 41.175 52.110 41.345 ;
        RECT 52.420 41.175 52.590 41.345 ;
        RECT 52.900 41.175 53.070 41.345 ;
        RECT 53.380 41.175 53.550 41.345 ;
        RECT 53.860 41.175 54.030 41.345 ;
        RECT 38.000 40.665 38.170 40.835 ;
        RECT 38.360 40.665 38.530 40.835 ;
        RECT 38.720 40.665 38.890 40.835 ;
        RECT 39.080 40.665 39.250 40.835 ;
        RECT 40.155 40.665 40.325 40.835 ;
        RECT 40.515 40.665 40.685 40.835 ;
        RECT 41.490 40.665 41.660 40.835 ;
        RECT 41.850 40.665 42.020 40.835 ;
        RECT 42.210 40.665 42.380 40.835 ;
        RECT 43.050 40.665 43.220 40.835 ;
        RECT 43.410 40.665 43.580 40.835 ;
        RECT 43.770 40.665 43.940 40.835 ;
        RECT 44.615 40.665 44.785 40.835 ;
        RECT 45.330 40.665 45.500 40.835 ;
        RECT 46.650 40.665 46.820 40.835 ;
        RECT 47.080 40.665 47.250 40.835 ;
        RECT 47.440 40.665 47.610 40.835 ;
        RECT 47.800 40.665 47.970 40.835 ;
        RECT 48.760 40.665 48.930 40.835 ;
        RECT 49.120 40.665 49.290 40.835 ;
        RECT 49.480 40.665 49.650 40.835 ;
        RECT 50.320 40.665 50.490 40.835 ;
        RECT 50.680 40.665 50.850 40.835 ;
        RECT 51.040 40.665 51.210 40.835 ;
        RECT 51.880 40.665 52.050 40.835 ;
        RECT 52.240 40.665 52.410 40.835 ;
        RECT 52.600 40.665 52.770 40.835 ;
        RECT 53.440 40.665 53.610 40.835 ;
        RECT 53.840 40.665 54.010 40.835 ;
      LAYER met1 ;
        RECT 36.420 40.625 54.205 41.390 ;
      LAYER via ;
        RECT 36.590 40.765 54.010 41.260 ;
      LAYER met2 ;
        RECT 36.420 40.625 54.205 41.390 ;
      LAYER via2 ;
        RECT 36.590 40.765 54.010 41.260 ;
      LAYER met3 ;
        RECT 36.420 40.625 54.205 41.390 ;
      LAYER via3 ;
        RECT 36.590 40.765 54.010 41.260 ;
      LAYER met4 ;
        RECT 36.205 39.810 55.900 41.455 ;
    END
  END vdd1v8
  PIN vss3v3
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 37.500 37.405 46.890 38.775 ;
        RECT 47.250 37.405 54.150 38.775 ;
        RECT 37.255 36.975 54.315 37.405 ;
        RECT 11.760 36.135 14.840 36.140 ;
        RECT 0.315 31.560 14.840 36.135 ;
        RECT 38.855 33.605 40.910 33.695 ;
        RECT 37.525 33.595 40.910 33.605 ;
        RECT 37.525 33.435 41.275 33.595 ;
        RECT 37.525 32.235 42.595 33.435 ;
        RECT 42.730 32.235 52.120 33.605 ;
        RECT 37.205 31.805 54.265 32.235 ;
        RECT 0.315 31.555 12.385 31.560 ;
        RECT 0.000 0.000 54.460 30.980 ;
      LAYER li1 ;
        RECT 38.060 37.740 39.310 38.575 ;
        RECT 40.150 37.950 40.880 38.635 ;
        RECT 39.990 37.740 40.880 37.950 ;
        RECT 41.430 37.740 42.440 38.635 ;
        RECT 42.990 37.740 44.000 38.635 ;
        RECT 44.550 37.740 45.560 38.635 ;
        RECT 46.520 37.790 46.890 38.635 ;
        RECT 46.360 37.740 46.890 37.790 ;
        RECT 38.060 37.570 46.890 37.740 ;
        RECT 47.080 37.740 47.970 38.575 ;
        RECT 48.560 37.740 49.570 38.235 ;
        RECT 50.120 37.740 51.130 38.235 ;
        RECT 51.680 37.740 52.730 38.235 ;
        RECT 53.720 37.740 54.090 38.235 ;
        RECT 47.080 37.570 54.090 37.740 ;
        RECT 37.385 37.105 54.185 37.275 ;
        RECT 12.000 35.895 14.600 35.900 ;
        RECT 0.175 35.730 14.600 35.895 ;
        RECT 0.175 35.725 12.170 35.730 ;
        RECT 0.175 31.965 0.725 35.725 ;
        RECT 2.315 32.825 2.485 34.865 ;
        RECT 2.985 31.965 3.175 35.725 ;
        RECT 4.765 32.825 4.935 34.865 ;
        RECT 6.945 32.825 7.115 34.865 ;
        RECT 9.125 32.825 9.295 34.865 ;
        RECT 11.305 32.825 11.475 34.865 ;
        RECT 11.975 31.970 12.170 35.725 ;
        RECT 12.670 32.830 12.840 34.870 ;
        RECT 14.430 34.190 14.600 35.730 ;
        RECT 14.430 31.970 35.670 34.190 ;
        RECT 40.455 32.395 41.965 33.305 ;
        RECT 43.290 32.570 44.540 33.405 ;
        RECT 45.380 32.780 46.110 33.465 ;
        RECT 45.220 32.570 46.110 32.780 ;
        RECT 46.660 32.570 47.670 33.465 ;
        RECT 48.220 32.570 49.230 33.465 ;
        RECT 49.780 32.570 50.790 33.465 ;
        RECT 51.750 32.620 52.120 33.465 ;
        RECT 51.590 32.570 52.120 32.620 ;
        RECT 43.290 32.400 52.120 32.570 ;
        RECT 11.975 31.965 35.670 31.970 ;
        RECT 0.175 31.940 35.670 31.965 ;
        RECT 37.335 31.940 54.135 32.105 ;
        RECT 0.175 30.715 54.300 31.940 ;
        RECT 0.175 30.630 54.280 30.715 ;
        RECT 0.175 30.150 3.445 30.630 ;
        RECT 0.175 29.065 3.450 30.150 ;
        RECT 0.180 1.905 0.350 29.065 ;
        RECT 0.830 27.990 1.520 29.065 ;
        RECT 2.760 27.990 3.450 29.065 ;
        RECT 52.940 30.145 53.630 30.150 ;
        RECT 54.110 30.145 54.280 30.630 ;
        RECT 52.940 29.065 54.280 30.145 ;
        RECT 52.940 27.990 53.630 29.065 ;
        RECT 0.830 1.905 1.520 2.990 ;
        RECT 0.180 0.830 1.520 1.905 ;
        RECT 52.940 1.905 53.630 2.990 ;
        RECT 54.110 1.905 54.280 29.065 ;
        RECT 52.940 0.830 54.280 1.905 ;
        RECT 0.180 0.825 1.170 0.830 ;
        RECT 53.275 0.825 54.280 0.830 ;
        RECT 0.180 0.350 0.350 0.825 ;
        RECT 54.110 0.350 54.280 0.825 ;
        RECT 0.180 0.180 54.280 0.350 ;
      LAYER mcon ;
        RECT 38.420 37.570 38.590 37.740 ;
        RECT 38.780 37.570 38.950 37.740 ;
        RECT 39.140 37.570 39.310 37.740 ;
        RECT 39.990 37.570 40.160 37.740 ;
        RECT 40.350 37.570 40.520 37.740 ;
        RECT 40.710 37.570 40.880 37.740 ;
        RECT 41.455 37.570 41.625 37.740 ;
        RECT 41.815 37.570 41.985 37.740 ;
        RECT 42.175 37.570 42.345 37.740 ;
        RECT 43.055 37.570 43.225 37.740 ;
        RECT 43.415 37.570 43.585 37.740 ;
        RECT 43.775 37.570 43.945 37.740 ;
        RECT 44.620 37.570 44.790 37.740 ;
        RECT 44.980 37.570 45.150 37.740 ;
        RECT 45.340 37.570 45.510 37.740 ;
        RECT 46.360 37.570 46.530 37.740 ;
        RECT 46.720 37.570 46.890 37.740 ;
        RECT 47.440 37.570 47.610 37.740 ;
        RECT 47.800 37.570 47.970 37.740 ;
        RECT 48.160 37.570 48.330 37.740 ;
        RECT 48.520 37.570 48.690 37.740 ;
        RECT 48.880 37.570 49.050 37.740 ;
        RECT 49.240 37.570 49.410 37.740 ;
        RECT 49.600 37.570 49.770 37.740 ;
        RECT 49.960 37.570 50.130 37.740 ;
        RECT 50.320 37.570 50.490 37.740 ;
        RECT 50.680 37.570 50.850 37.740 ;
        RECT 51.040 37.570 51.210 37.740 ;
        RECT 51.400 37.570 51.570 37.740 ;
        RECT 51.760 37.570 51.930 37.740 ;
        RECT 52.120 37.570 52.290 37.740 ;
        RECT 52.480 37.570 52.650 37.740 ;
        RECT 52.840 37.570 53.010 37.740 ;
        RECT 53.200 37.570 53.370 37.740 ;
        RECT 53.560 37.570 53.730 37.740 ;
        RECT 53.920 37.570 54.090 37.740 ;
        RECT 37.540 37.105 37.710 37.275 ;
        RECT 38.020 37.105 38.190 37.275 ;
        RECT 38.500 37.105 38.670 37.275 ;
        RECT 38.980 37.105 39.150 37.275 ;
        RECT 39.460 37.105 39.630 37.275 ;
        RECT 39.940 37.105 40.110 37.275 ;
        RECT 40.420 37.105 40.590 37.275 ;
        RECT 40.900 37.105 41.070 37.275 ;
        RECT 41.380 37.105 41.550 37.275 ;
        RECT 41.860 37.105 42.030 37.275 ;
        RECT 42.340 37.105 42.510 37.275 ;
        RECT 42.820 37.105 42.990 37.275 ;
        RECT 43.300 37.105 43.470 37.275 ;
        RECT 43.780 37.105 43.950 37.275 ;
        RECT 44.260 37.105 44.430 37.275 ;
        RECT 44.740 37.105 44.910 37.275 ;
        RECT 45.220 37.105 45.390 37.275 ;
        RECT 45.700 37.105 45.870 37.275 ;
        RECT 46.180 37.105 46.350 37.275 ;
        RECT 46.660 37.105 46.830 37.275 ;
        RECT 47.140 37.105 47.310 37.275 ;
        RECT 47.620 37.105 47.790 37.275 ;
        RECT 48.100 37.105 48.270 37.275 ;
        RECT 48.580 37.105 48.750 37.275 ;
        RECT 49.060 37.105 49.230 37.275 ;
        RECT 49.540 37.105 49.710 37.275 ;
        RECT 50.020 37.105 50.190 37.275 ;
        RECT 50.500 37.105 50.670 37.275 ;
        RECT 50.980 37.105 51.150 37.275 ;
        RECT 51.460 37.105 51.630 37.275 ;
        RECT 51.940 37.105 52.110 37.275 ;
        RECT 52.420 37.105 52.590 37.275 ;
        RECT 52.900 37.105 53.070 37.275 ;
        RECT 53.380 37.105 53.550 37.275 ;
        RECT 53.860 37.105 54.030 37.275 ;
        RECT 2.315 32.905 2.485 34.785 ;
        RECT 3.005 32.530 3.175 35.160 ;
        RECT 4.765 32.990 4.935 33.740 ;
        RECT 6.945 32.990 7.115 33.740 ;
        RECT 9.125 32.990 9.295 33.740 ;
        RECT 11.305 32.990 11.475 33.740 ;
        RECT 12.000 31.970 12.170 33.660 ;
        RECT 12.670 32.910 12.840 34.790 ;
        RECT 0.240 30.960 1.430 31.590 ;
        RECT 2.525 30.955 14.755 31.600 ;
        RECT 16.100 31.265 30.580 33.465 ;
        RECT 40.545 32.445 40.715 32.615 ;
        RECT 40.905 32.445 41.075 32.615 ;
        RECT 41.315 32.445 41.485 32.615 ;
        RECT 41.745 32.445 41.915 32.615 ;
        RECT 43.650 32.400 43.820 32.570 ;
        RECT 44.010 32.400 44.180 32.570 ;
        RECT 44.370 32.400 44.540 32.570 ;
        RECT 45.220 32.400 45.390 32.570 ;
        RECT 45.580 32.400 45.750 32.570 ;
        RECT 45.940 32.400 46.110 32.570 ;
        RECT 46.685 32.400 46.855 32.570 ;
        RECT 47.045 32.400 47.215 32.570 ;
        RECT 47.405 32.400 47.575 32.570 ;
        RECT 48.285 32.400 48.455 32.570 ;
        RECT 48.645 32.400 48.815 32.570 ;
        RECT 49.005 32.400 49.175 32.570 ;
        RECT 49.850 32.400 50.020 32.570 ;
        RECT 50.210 32.400 50.380 32.570 ;
        RECT 50.570 32.400 50.740 32.570 ;
        RECT 51.590 32.400 51.760 32.570 ;
        RECT 51.950 32.400 52.120 32.570 ;
        RECT 37.490 31.935 37.660 32.105 ;
        RECT 37.970 31.935 38.140 32.105 ;
        RECT 38.450 31.935 38.620 32.105 ;
        RECT 38.930 31.935 39.100 32.105 ;
        RECT 39.410 31.935 39.580 32.105 ;
        RECT 39.890 31.935 40.060 32.105 ;
        RECT 40.370 31.935 40.540 32.105 ;
        RECT 40.850 31.935 41.020 32.105 ;
        RECT 41.330 31.935 41.500 32.105 ;
        RECT 41.810 31.935 41.980 32.105 ;
        RECT 42.290 31.935 42.460 32.105 ;
        RECT 42.770 31.935 42.940 32.105 ;
        RECT 43.250 31.935 43.420 32.105 ;
        RECT 43.730 31.935 43.900 32.105 ;
        RECT 44.210 31.935 44.380 32.105 ;
        RECT 44.690 31.935 44.860 32.105 ;
        RECT 45.170 31.935 45.340 32.105 ;
        RECT 45.650 31.935 45.820 32.105 ;
        RECT 46.130 31.935 46.300 32.105 ;
        RECT 46.610 31.935 46.780 32.105 ;
        RECT 47.090 31.935 47.260 32.105 ;
        RECT 47.570 31.935 47.740 32.105 ;
        RECT 48.050 31.935 48.220 32.105 ;
        RECT 48.530 31.935 48.700 32.105 ;
        RECT 49.010 31.935 49.180 32.105 ;
        RECT 49.490 31.935 49.660 32.105 ;
        RECT 49.970 31.935 50.140 32.105 ;
        RECT 50.450 31.935 50.620 32.105 ;
        RECT 50.930 31.935 51.100 32.105 ;
        RECT 51.410 31.935 51.580 32.105 ;
        RECT 51.890 31.935 52.060 32.105 ;
        RECT 52.370 31.935 52.540 32.105 ;
        RECT 52.850 31.935 53.020 32.105 ;
        RECT 53.330 31.935 53.500 32.105 ;
        RECT 53.810 31.935 53.980 32.105 ;
        RECT 0.180 1.865 0.350 29.115 ;
        RECT 54.110 1.865 54.280 29.115 ;
        RECT 3.040 0.180 51.420 0.350 ;
      LAYER met1 ;
        RECT 36.395 37.815 54.180 37.850 ;
        RECT 36.395 37.445 54.185 37.815 ;
        RECT 36.395 37.305 54.180 37.445 ;
        RECT 36.395 37.085 54.185 37.305 ;
        RECT 37.385 37.075 54.185 37.085 ;
        RECT 2.975 34.860 3.205 35.220 ;
        RECT 2.315 34.845 3.205 34.860 ;
        RECT 2.285 33.725 3.205 34.845 ;
        RECT 4.735 33.725 4.965 33.800 ;
        RECT 6.915 33.725 7.145 33.800 ;
        RECT 9.095 33.725 9.325 33.800 ;
        RECT 11.275 33.725 11.505 33.800 ;
        RECT 12.640 33.725 12.870 34.850 ;
        RECT 2.285 32.895 12.870 33.725 ;
        RECT 2.285 32.845 3.205 32.895 ;
        RECT 2.525 32.470 3.205 32.845 ;
        RECT 2.525 31.630 3.170 32.470 ;
        RECT 11.970 31.910 12.200 32.895 ;
        RECT 12.640 32.850 12.870 32.895 ;
        RECT 15.835 32.655 30.870 34.210 ;
        RECT 15.835 31.630 54.135 32.655 ;
        RECT 0.125 30.925 1.505 31.630 ;
        RECT 2.465 31.595 54.135 31.630 ;
        RECT 2.465 31.185 30.870 31.595 ;
        RECT 2.465 30.925 30.875 31.185 ;
        RECT 0.125 26.740 0.665 30.925 ;
        RECT 54.025 26.740 54.335 30.395 ;
        RECT 0.125 23.740 54.335 26.740 ;
        RECT 0.125 21.740 0.665 23.740 ;
        RECT 54.025 21.740 54.335 23.740 ;
        RECT 0.125 18.740 54.335 21.740 ;
        RECT 0.125 16.740 0.665 18.740 ;
        RECT 54.025 16.740 54.335 18.740 ;
        RECT 0.125 13.740 54.335 16.740 ;
        RECT 0.125 11.740 0.665 13.740 ;
        RECT 54.025 11.740 54.335 13.740 ;
        RECT 0.125 8.740 54.335 11.740 ;
        RECT 0.125 6.740 0.665 8.740 ;
        RECT 54.025 6.740 54.335 8.740 ;
        RECT 0.125 3.740 54.335 6.740 ;
        RECT 0.125 0.495 0.665 3.740 ;
        RECT 54.025 0.495 54.335 3.740 ;
        RECT 0.125 0.055 54.335 0.495 ;
      LAYER via ;
        RECT 36.530 37.245 41.715 37.715 ;
        RECT 43.090 37.245 53.245 37.715 ;
        RECT 21.655 31.350 26.390 34.095 ;
      LAYER met2 ;
        RECT 36.395 37.085 41.870 37.850 ;
        RECT 42.940 37.715 53.335 37.850 ;
        RECT 42.935 37.245 53.335 37.715 ;
        RECT 42.940 37.085 53.335 37.245 ;
        RECT 21.540 31.245 26.490 34.340 ;
      LAYER via2 ;
        RECT 36.530 37.245 41.715 37.715 ;
        RECT 43.090 37.245 53.245 37.715 ;
        RECT 21.655 32.610 26.390 34.245 ;
      LAYER met3 ;
        RECT 36.395 37.085 53.335 37.850 ;
        RECT 20.555 32.470 26.495 36.585 ;
        RECT 20.555 31.255 21.535 32.470 ;
        RECT 19.455 0.255 50.815 31.255 ;
      LAYER via3 ;
        RECT 36.530 37.245 53.245 37.715 ;
        RECT 21.750 32.790 26.340 36.385 ;
        RECT 19.555 0.395 19.875 31.115 ;
      LAYER met4 ;
        RECT 0.190 36.275 53.335 38.275 ;
        RECT 19.085 32.610 26.495 36.275 ;
        RECT 19.085 0.255 20.055 32.610 ;
      LAYER via4 ;
        RECT 21.750 32.790 26.340 36.235 ;
      LAYER met5 ;
        RECT 21.565 32.470 26.495 36.585 ;
        RECT 22.535 30.675 26.495 32.470 ;
        RECT 24.535 0.835 51.415 30.675 ;
    END
  END vss3v3
  PIN porb_h
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER li1 ;
        RECT 46.220 34.225 46.550 35.465 ;
        RECT 47.780 34.225 48.110 35.465 ;
        RECT 49.340 34.225 49.670 35.465 ;
        RECT 50.900 35.250 51.350 35.465 ;
        RECT 50.900 34.225 51.580 35.250 ;
        RECT 46.220 34.055 51.580 34.225 ;
        RECT 46.280 33.645 51.170 33.815 ;
        RECT 46.280 32.825 46.490 33.645 ;
        RECT 47.840 32.825 48.050 33.645 ;
        RECT 49.400 32.825 49.610 33.645 ;
        RECT 50.960 32.995 51.170 33.645 ;
        RECT 51.350 32.995 51.580 34.055 ;
        RECT 50.960 32.825 51.580 32.995 ;
      LAYER mcon ;
        RECT 51.350 33.675 51.580 34.480 ;
      LAYER met1 ;
        RECT 51.320 34.170 51.610 34.540 ;
        RECT 51.320 33.825 53.410 34.170 ;
        RECT 51.320 33.615 51.610 33.825 ;
      LAYER via ;
        RECT 52.535 33.825 53.360 34.170 ;
      LAYER met2 ;
        RECT 52.490 33.825 54.590 34.170 ;
      LAYER via2 ;
        RECT 53.785 33.825 54.545 34.170 ;
      LAYER met3 ;
        RECT 53.735 34.170 54.590 34.200 ;
        RECT 53.735 33.825 56.710 34.170 ;
        RECT 53.735 33.790 54.590 33.825 ;
    END
  END porb_h
  PIN por_l
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER li1 ;
        RECT 48.260 39.395 48.590 40.635 ;
        RECT 49.820 39.395 50.150 40.635 ;
        RECT 51.380 39.395 51.710 40.635 ;
        RECT 52.940 39.395 53.270 40.635 ;
        RECT 48.260 39.225 54.095 39.395 ;
        RECT 48.180 38.585 53.210 38.590 ;
        RECT 53.925 38.585 54.095 39.225 ;
        RECT 48.180 38.420 54.095 38.585 ;
        RECT 48.180 37.920 48.390 38.420 ;
        RECT 49.740 37.920 49.950 38.420 ;
        RECT 51.300 37.920 51.510 38.420 ;
        RECT 52.900 38.415 54.095 38.420 ;
        RECT 52.900 37.920 53.550 38.415 ;
      LAYER mcon ;
        RECT 53.925 38.415 54.095 39.395 ;
      LAYER met1 ;
        RECT 53.895 38.640 54.125 39.455 ;
        RECT 53.715 38.370 54.575 38.640 ;
        RECT 53.895 38.355 54.125 38.370 ;
      LAYER via ;
        RECT 53.765 38.370 54.525 38.640 ;
      LAYER met2 ;
        RECT 53.765 38.305 54.525 38.705 ;
      LAYER via2 ;
        RECT 53.765 38.355 54.525 38.655 ;
      LAYER met3 ;
        RECT 53.715 38.330 54.550 38.695 ;
        RECT 53.960 37.755 54.260 38.330 ;
        RECT 53.960 37.455 56.720 37.755 ;
    END
  END por_l
  PIN porb_l
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER li1 ;
        RECT 40.990 39.395 41.320 40.635 ;
        RECT 42.550 39.395 42.880 40.635 ;
        RECT 44.110 39.395 44.440 40.635 ;
        RECT 45.670 40.420 46.120 40.635 ;
        RECT 45.670 39.395 46.350 40.420 ;
        RECT 40.990 39.225 46.350 39.395 ;
        RECT 41.050 38.815 45.940 38.985 ;
        RECT 41.050 37.995 41.260 38.815 ;
        RECT 42.610 37.995 42.820 38.815 ;
        RECT 44.170 37.995 44.380 38.815 ;
        RECT 45.730 38.165 45.940 38.815 ;
        RECT 46.120 38.165 46.350 39.225 ;
        RECT 45.730 37.995 46.350 38.165 ;
      LAYER mcon ;
        RECT 46.120 39.270 46.350 40.300 ;
      LAYER met1 ;
        RECT 46.090 40.255 46.380 40.360 ;
        RECT 50.640 40.255 51.500 40.265 ;
        RECT 46.090 40.005 51.500 40.255 ;
        RECT 46.090 39.210 46.380 40.005 ;
        RECT 50.640 39.995 51.500 40.005 ;
      LAYER via ;
        RECT 50.690 39.995 51.450 40.265 ;
      LAYER met2 ;
        RECT 50.690 39.930 51.450 40.330 ;
      LAYER via2 ;
        RECT 50.690 39.980 51.450 40.280 ;
      LAYER met3 ;
        RECT 50.640 40.280 51.475 40.320 ;
        RECT 50.640 39.980 52.155 40.280 ;
        RECT 50.640 39.955 51.475 39.980 ;
        RECT 51.855 39.580 52.155 39.980 ;
        RECT 51.855 39.280 56.715 39.580 ;
    END
  END porb_l
  PIN vss1v8
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT -0.070 42.760 56.090 43.380 ;
      LAYER mcon ;
        RECT 0.130 42.760 55.890 43.380 ;
      LAYER met1 ;
        RECT -0.070 42.720 56.090 43.420 ;
    END
  END vss1v8
  OBS
      LAYER li1 ;
        RECT 1.640 40.440 2.440 40.610 ;
        RECT 4.070 40.440 4.870 40.610 ;
        RECT 5.160 40.440 5.960 40.610 ;
        RECT 6.250 40.440 7.050 40.610 ;
        RECT 7.340 40.440 8.140 40.610 ;
        RECT 8.430 40.440 9.230 40.610 ;
        RECT 9.520 40.440 10.320 40.610 ;
        RECT 10.610 40.440 11.410 40.610 ;
        RECT 11.700 40.440 12.500 40.610 ;
        RECT 14.130 40.440 14.930 40.610 ;
        RECT 16.560 40.440 17.360 40.610 ;
        RECT 18.990 40.440 19.790 40.610 ;
        RECT 21.420 40.440 22.220 40.610 ;
        RECT 22.510 40.440 23.310 40.610 ;
        RECT 23.600 40.440 24.400 40.610 ;
        RECT 24.690 40.440 25.490 40.610 ;
        RECT 25.780 40.440 26.580 40.610 ;
        RECT 26.870 40.440 27.670 40.610 ;
        RECT 27.960 40.440 28.760 40.610 ;
        RECT 30.390 40.440 31.190 40.610 ;
        RECT 32.820 40.440 33.620 40.610 ;
        RECT 1.410 38.185 1.580 40.225 ;
        RECT 2.500 38.185 2.670 40.225 ;
        RECT 4.930 38.185 5.100 40.225 ;
        RECT 7.110 38.185 7.280 40.225 ;
        RECT 9.290 38.185 9.460 40.225 ;
        RECT 11.470 38.185 11.640 40.225 ;
        RECT 14.990 38.185 15.160 40.225 ;
        RECT 16.330 38.185 16.500 40.225 ;
        RECT 17.420 38.185 17.590 40.225 ;
        RECT 18.760 38.185 18.930 40.225 ;
        RECT 19.850 38.185 20.020 40.225 ;
        RECT 22.280 38.185 22.450 40.225 ;
        RECT 24.460 38.185 24.630 40.225 ;
        RECT 26.640 38.185 26.810 40.225 ;
        RECT 28.820 38.185 28.990 40.225 ;
        RECT 31.250 38.185 31.420 40.225 ;
        RECT 32.590 38.185 32.760 40.225 ;
        RECT 33.680 38.185 33.850 40.225 ;
        RECT 37.630 39.455 37.820 40.735 ;
        RECT 39.430 39.455 39.980 40.635 ;
        RECT 37.630 39.285 39.980 39.455 ;
        RECT 37.630 38.665 37.820 39.285 ;
        RECT 39.810 39.145 39.980 39.285 ;
        RECT 38.020 38.770 39.630 39.005 ;
        RECT 39.810 38.815 40.765 39.145 ;
        RECT 37.630 37.995 37.840 38.665 ;
        RECT 39.810 38.590 39.980 38.815 ;
        RECT 47.295 38.770 53.745 39.005 ;
        RECT 39.490 38.420 39.980 38.590 ;
        RECT 1.640 37.800 2.440 37.970 ;
        RECT 4.070 37.800 4.870 37.970 ;
        RECT 5.160 37.800 5.960 37.970 ;
        RECT 6.250 37.800 7.050 37.970 ;
        RECT 7.340 37.800 8.140 37.970 ;
        RECT 8.430 37.800 9.230 37.970 ;
        RECT 9.520 37.800 10.320 37.970 ;
        RECT 10.610 37.800 11.410 37.970 ;
        RECT 11.700 37.800 12.500 37.970 ;
        RECT 14.130 37.800 14.930 37.970 ;
        RECT 16.560 37.800 17.360 37.970 ;
        RECT 18.990 37.800 19.790 37.970 ;
        RECT 21.420 37.800 22.220 37.970 ;
        RECT 22.510 37.800 23.310 37.970 ;
        RECT 23.600 37.800 24.400 37.970 ;
        RECT 24.690 37.800 25.490 37.970 ;
        RECT 25.780 37.800 26.580 37.970 ;
        RECT 26.870 37.800 27.670 37.970 ;
        RECT 27.960 37.800 28.760 37.970 ;
        RECT 30.390 37.800 31.190 37.970 ;
        RECT 32.820 37.800 33.620 37.970 ;
        RECT 39.490 37.920 39.700 38.420 ;
        RECT 38.075 35.675 38.365 35.755 ;
        RECT 37.420 35.505 38.365 35.675 ;
        RECT 1.455 35.035 2.255 35.205 ;
        RECT 3.905 35.035 4.705 35.205 ;
        RECT 4.995 35.035 5.795 35.205 ;
        RECT 6.085 35.035 6.885 35.205 ;
        RECT 7.175 35.035 7.975 35.205 ;
        RECT 8.265 35.035 9.065 35.205 ;
        RECT 9.355 35.035 10.155 35.205 ;
        RECT 10.445 35.035 11.245 35.205 ;
        RECT 12.900 35.040 13.700 35.210 ;
        RECT 1.225 32.825 1.395 34.865 ;
        RECT 3.675 32.825 3.845 34.865 ;
        RECT 5.855 32.825 6.025 34.865 ;
        RECT 8.035 32.825 8.205 34.865 ;
        RECT 10.215 32.825 10.385 34.865 ;
        RECT 13.760 32.830 13.930 34.870 ;
        RECT 37.420 33.995 37.590 35.505 ;
        RECT 38.075 35.425 38.365 35.505 ;
        RECT 38.535 35.255 40.125 35.425 ;
        RECT 37.765 34.355 38.015 35.105 ;
        RECT 37.765 34.185 38.210 34.355 ;
        RECT 38.535 34.315 38.795 35.255 ;
        RECT 38.990 34.350 39.345 35.085 ;
        RECT 37.420 33.825 37.865 33.995 ;
        RECT 37.615 33.110 37.865 33.825 ;
        RECT 38.040 32.815 38.210 34.185 ;
        RECT 38.990 34.005 39.170 34.350 ;
        RECT 39.795 34.340 40.125 35.255 ;
        RECT 38.380 33.705 39.170 34.005 ;
        RECT 39.350 33.875 40.640 34.170 ;
        RECT 41.190 33.705 42.025 34.075 ;
        RECT 38.380 33.675 42.025 33.705 ;
        RECT 38.935 33.665 42.025 33.675 ;
        RECT 38.935 33.525 41.545 33.665 ;
        RECT 38.395 33.165 38.725 33.430 ;
        RECT 38.935 33.335 39.275 33.525 ;
        RECT 39.725 33.165 40.055 33.355 ;
        RECT 38.395 32.995 40.055 33.165 ;
        RECT 1.455 32.485 2.255 32.655 ;
        RECT 3.905 32.485 4.705 32.655 ;
        RECT 4.995 32.485 5.795 32.655 ;
        RECT 6.085 32.485 6.885 32.655 ;
        RECT 7.175 32.485 7.975 32.655 ;
        RECT 8.265 32.485 9.065 32.655 ;
        RECT 9.355 32.485 10.155 32.655 ;
        RECT 10.445 32.485 11.245 32.655 ;
        RECT 12.900 32.490 13.700 32.660 ;
        RECT 38.040 32.590 39.345 32.815 ;
        RECT 42.195 32.535 42.530 35.735 ;
        RECT 42.860 34.285 43.050 35.565 ;
        RECT 44.660 34.285 45.210 35.465 ;
        RECT 42.860 34.115 45.210 34.285 ;
        RECT 42.860 33.495 43.050 34.115 ;
        RECT 45.040 33.975 45.210 34.115 ;
        RECT 43.250 33.600 44.860 33.835 ;
        RECT 45.040 33.645 45.995 33.975 ;
        RECT 42.860 32.825 43.070 33.495 ;
        RECT 45.040 33.420 45.210 33.645 ;
        RECT 44.720 33.250 45.210 33.420 ;
        RECT 44.720 32.750 44.930 33.250 ;
        RECT 4.690 30.145 5.380 30.150 ;
        RECT 6.620 30.145 7.310 30.150 ;
        RECT 4.690 29.065 7.310 30.145 ;
        RECT 4.690 27.990 5.380 29.065 ;
        RECT 6.620 27.990 7.310 29.065 ;
        RECT 8.550 30.145 9.240 30.150 ;
        RECT 10.480 30.145 11.170 30.150 ;
        RECT 8.550 29.065 11.170 30.145 ;
        RECT 8.550 27.990 9.240 29.065 ;
        RECT 10.480 27.990 11.170 29.065 ;
        RECT 12.410 30.145 13.100 30.150 ;
        RECT 14.340 30.145 15.030 30.150 ;
        RECT 12.410 29.065 15.030 30.145 ;
        RECT 12.410 27.990 13.100 29.065 ;
        RECT 14.340 27.990 15.030 29.065 ;
        RECT 16.270 30.145 16.960 30.150 ;
        RECT 18.200 30.145 18.890 30.150 ;
        RECT 16.270 29.065 18.890 30.145 ;
        RECT 16.270 27.990 16.960 29.065 ;
        RECT 18.200 27.990 18.890 29.065 ;
        RECT 20.130 30.145 20.820 30.150 ;
        RECT 22.060 30.145 22.750 30.150 ;
        RECT 20.130 29.065 22.750 30.145 ;
        RECT 20.130 27.990 20.820 29.065 ;
        RECT 22.060 27.990 22.750 29.065 ;
        RECT 23.990 30.145 24.680 30.150 ;
        RECT 25.920 30.145 26.610 30.150 ;
        RECT 23.990 29.065 26.610 30.145 ;
        RECT 23.990 27.990 24.680 29.065 ;
        RECT 25.920 27.990 26.610 29.065 ;
        RECT 27.850 30.145 28.540 30.150 ;
        RECT 29.780 30.145 30.470 30.150 ;
        RECT 27.850 29.065 30.470 30.145 ;
        RECT 27.850 27.990 28.540 29.065 ;
        RECT 29.780 27.990 30.470 29.065 ;
        RECT 31.710 30.145 32.400 30.150 ;
        RECT 33.640 30.145 34.330 30.150 ;
        RECT 31.710 29.065 34.330 30.145 ;
        RECT 31.710 27.990 32.400 29.065 ;
        RECT 33.640 27.990 34.330 29.065 ;
        RECT 35.570 30.145 36.260 30.150 ;
        RECT 37.500 30.145 38.190 30.150 ;
        RECT 35.570 29.065 38.190 30.145 ;
        RECT 35.570 27.990 36.260 29.065 ;
        RECT 37.500 27.990 38.190 29.065 ;
        RECT 39.430 30.145 40.120 30.150 ;
        RECT 41.360 30.145 42.050 30.150 ;
        RECT 39.430 29.065 42.050 30.145 ;
        RECT 39.430 27.990 40.120 29.065 ;
        RECT 41.360 27.990 42.050 29.065 ;
        RECT 43.290 30.145 43.980 30.150 ;
        RECT 45.220 30.145 45.910 30.150 ;
        RECT 43.290 29.065 45.910 30.145 ;
        RECT 43.290 27.990 43.980 29.065 ;
        RECT 45.220 27.990 45.910 29.065 ;
        RECT 47.150 30.145 47.840 30.150 ;
        RECT 49.080 30.145 49.770 30.150 ;
        RECT 47.150 29.065 49.770 30.145 ;
        RECT 47.150 27.990 47.840 29.065 ;
        RECT 49.080 27.990 49.770 29.065 ;
        RECT 2.760 1.905 3.450 2.990 ;
        RECT 4.690 1.905 5.380 2.990 ;
        RECT 2.760 0.830 5.380 1.905 ;
        RECT 6.620 1.905 7.310 2.990 ;
        RECT 8.550 1.905 9.240 2.990 ;
        RECT 6.620 0.830 9.240 1.905 ;
        RECT 10.480 1.905 11.170 2.990 ;
        RECT 12.410 1.905 13.100 2.990 ;
        RECT 10.480 0.830 13.100 1.905 ;
        RECT 14.340 1.905 15.030 2.990 ;
        RECT 16.270 1.905 16.960 2.990 ;
        RECT 14.340 0.830 16.960 1.905 ;
        RECT 18.200 1.905 18.890 2.990 ;
        RECT 20.130 1.905 20.820 2.990 ;
        RECT 18.200 0.830 20.820 1.905 ;
        RECT 22.060 1.905 22.750 2.990 ;
        RECT 23.990 1.905 24.680 2.990 ;
        RECT 22.060 0.830 24.680 1.905 ;
        RECT 25.920 1.905 26.610 2.990 ;
        RECT 27.850 1.905 28.540 2.990 ;
        RECT 25.920 0.830 28.540 1.905 ;
        RECT 29.780 1.905 30.470 2.990 ;
        RECT 31.710 1.905 32.400 2.990 ;
        RECT 29.780 0.830 32.400 1.905 ;
        RECT 33.640 1.905 34.330 2.990 ;
        RECT 35.570 1.905 36.260 2.990 ;
        RECT 33.640 0.830 36.260 1.905 ;
        RECT 37.500 1.905 38.190 2.990 ;
        RECT 39.430 1.905 40.120 2.990 ;
        RECT 37.500 0.830 40.120 1.905 ;
        RECT 41.360 1.905 42.050 2.990 ;
        RECT 43.290 1.905 43.980 2.990 ;
        RECT 41.360 0.830 43.980 1.905 ;
        RECT 45.220 1.905 45.910 2.990 ;
        RECT 47.150 1.905 47.840 2.990 ;
        RECT 45.220 0.830 47.840 1.905 ;
        RECT 49.080 1.905 49.770 2.990 ;
        RECT 51.010 1.905 51.700 2.990 ;
        RECT 49.080 0.830 51.700 1.905 ;
        RECT 3.095 0.825 5.030 0.830 ;
        RECT 6.955 0.825 8.890 0.830 ;
        RECT 10.815 0.825 12.750 0.830 ;
        RECT 14.675 0.825 16.610 0.830 ;
        RECT 18.535 0.825 20.470 0.830 ;
        RECT 22.395 0.825 24.330 0.830 ;
        RECT 26.255 0.825 28.190 0.830 ;
        RECT 30.115 0.825 32.050 0.830 ;
        RECT 33.975 0.825 35.910 0.830 ;
        RECT 37.835 0.825 39.770 0.830 ;
        RECT 41.695 0.825 43.630 0.830 ;
        RECT 45.555 0.825 47.490 0.830 ;
        RECT 49.415 0.825 51.350 0.830 ;
      LAYER mcon ;
        RECT 1.720 40.440 2.360 40.610 ;
        RECT 4.150 40.440 4.790 40.610 ;
        RECT 5.240 40.440 5.880 40.610 ;
        RECT 6.330 40.440 6.970 40.610 ;
        RECT 7.420 40.440 8.060 40.610 ;
        RECT 8.510 40.440 9.150 40.610 ;
        RECT 9.600 40.440 10.240 40.610 ;
        RECT 10.690 40.440 11.330 40.610 ;
        RECT 11.780 40.440 12.420 40.610 ;
        RECT 14.210 40.440 14.850 40.610 ;
        RECT 16.640 40.440 17.280 40.610 ;
        RECT 19.070 40.440 19.710 40.610 ;
        RECT 21.500 40.440 22.140 40.610 ;
        RECT 22.590 40.440 23.230 40.610 ;
        RECT 23.680 40.440 24.320 40.610 ;
        RECT 24.770 40.440 25.410 40.610 ;
        RECT 25.860 40.440 26.500 40.610 ;
        RECT 26.950 40.440 27.590 40.610 ;
        RECT 28.040 40.440 28.680 40.610 ;
        RECT 30.470 40.440 31.110 40.610 ;
        RECT 32.900 40.440 33.540 40.610 ;
        RECT 1.410 38.265 1.580 40.145 ;
        RECT 2.500 38.265 2.670 40.145 ;
        RECT 4.930 38.350 5.100 39.100 ;
        RECT 7.110 38.350 7.280 39.100 ;
        RECT 9.290 38.350 9.460 39.100 ;
        RECT 11.470 38.350 11.640 39.100 ;
        RECT 14.990 38.265 15.160 40.145 ;
        RECT 16.330 38.265 16.500 40.145 ;
        RECT 17.420 38.265 17.590 40.145 ;
        RECT 18.760 38.265 18.930 40.145 ;
        RECT 19.850 38.265 20.020 40.145 ;
        RECT 22.280 38.350 22.450 39.100 ;
        RECT 24.460 38.350 24.630 39.100 ;
        RECT 26.640 38.350 26.810 39.100 ;
        RECT 28.820 38.350 28.990 39.100 ;
        RECT 31.250 38.265 31.420 40.145 ;
        RECT 32.590 38.265 32.760 40.145 ;
        RECT 33.680 38.265 33.850 40.145 ;
        RECT 1.720 37.800 2.360 37.970 ;
        RECT 4.150 37.800 4.790 37.970 ;
        RECT 5.240 37.800 5.880 37.970 ;
        RECT 6.330 37.800 6.970 37.970 ;
        RECT 7.420 37.800 8.060 37.970 ;
        RECT 8.510 37.800 9.150 37.970 ;
        RECT 9.600 37.800 10.240 37.970 ;
        RECT 10.690 37.800 11.330 37.970 ;
        RECT 11.780 37.800 12.420 37.970 ;
        RECT 14.210 37.800 14.850 37.970 ;
        RECT 16.640 37.800 17.280 37.970 ;
        RECT 19.070 37.800 19.710 37.970 ;
        RECT 21.500 37.800 22.140 37.970 ;
        RECT 22.590 37.800 23.230 37.970 ;
        RECT 23.680 37.800 24.320 37.970 ;
        RECT 24.770 37.800 25.410 37.970 ;
        RECT 25.860 37.800 26.500 37.970 ;
        RECT 26.950 37.800 27.590 37.970 ;
        RECT 28.040 37.800 28.680 37.970 ;
        RECT 30.470 37.800 31.110 37.970 ;
        RECT 32.900 37.800 33.540 37.970 ;
        RECT 1.535 35.035 2.175 35.205 ;
        RECT 3.985 35.035 4.625 35.205 ;
        RECT 5.075 35.035 5.715 35.205 ;
        RECT 6.165 35.035 6.805 35.205 ;
        RECT 7.255 35.035 7.895 35.205 ;
        RECT 8.345 35.035 8.985 35.205 ;
        RECT 9.435 35.035 10.075 35.205 ;
        RECT 10.525 35.035 11.165 35.205 ;
        RECT 12.980 35.040 13.620 35.210 ;
        RECT 1.225 32.905 1.395 34.785 ;
        RECT 3.675 33.950 3.845 34.700 ;
        RECT 5.855 33.950 6.025 34.700 ;
        RECT 8.035 33.950 8.205 34.700 ;
        RECT 10.215 33.950 10.385 34.700 ;
        RECT 13.760 32.910 13.930 34.790 ;
        RECT 39.350 33.875 40.640 34.170 ;
        RECT 42.195 33.420 42.530 34.390 ;
        RECT 1.535 32.485 2.175 32.655 ;
        RECT 3.985 32.485 4.625 32.655 ;
        RECT 5.075 32.485 5.715 32.655 ;
        RECT 6.165 32.485 6.805 32.655 ;
        RECT 7.255 32.485 7.895 32.655 ;
        RECT 8.345 32.485 8.985 32.655 ;
        RECT 9.435 32.485 10.075 32.655 ;
        RECT 10.525 32.485 11.165 32.655 ;
        RECT 12.980 32.490 13.620 32.660 ;
        RECT 13.240 29.145 14.200 30.075 ;
      LAYER met1 ;
        RECT 3.545 40.645 4.090 40.720 ;
        RECT 1.660 40.635 2.420 40.640 ;
        RECT 1.090 40.410 2.420 40.635 ;
        RECT 3.545 40.425 12.490 40.645 ;
        RECT 14.145 40.425 14.950 40.645 ;
        RECT 3.545 40.410 4.850 40.425 ;
        RECT 5.180 40.410 5.940 40.425 ;
        RECT 6.270 40.410 7.030 40.425 ;
        RECT 7.360 40.410 8.120 40.425 ;
        RECT 8.450 40.410 9.210 40.425 ;
        RECT 9.540 40.410 10.300 40.425 ;
        RECT 10.630 40.410 11.390 40.425 ;
        RECT 11.720 40.410 12.480 40.425 ;
        RECT 14.150 40.410 14.910 40.425 ;
        RECT 16.580 40.410 17.340 40.640 ;
        RECT 18.495 40.410 19.795 40.640 ;
        RECT 21.440 40.625 22.200 40.640 ;
        RECT 22.530 40.625 23.290 40.640 ;
        RECT 23.620 40.625 24.380 40.640 ;
        RECT 24.710 40.625 25.470 40.640 ;
        RECT 25.800 40.625 26.560 40.640 ;
        RECT 26.890 40.625 27.650 40.640 ;
        RECT 27.980 40.625 28.740 40.640 ;
        RECT 21.415 40.410 28.740 40.625 ;
        RECT 30.410 40.625 31.170 40.640 ;
        RECT 30.410 40.410 31.185 40.625 ;
        RECT 32.840 40.410 33.600 40.640 ;
        RECT 1.090 40.190 2.180 40.410 ;
        RECT 1.090 38.205 1.610 40.190 ;
        RECT 1.875 38.205 2.180 40.190 ;
        RECT 2.470 40.200 2.700 40.205 ;
        RECT 2.470 38.940 2.835 40.200 ;
        RECT 4.900 38.940 5.130 39.160 ;
        RECT 7.080 38.940 7.310 39.160 ;
        RECT 9.260 38.940 9.490 39.160 ;
        RECT 11.440 38.940 11.670 39.160 ;
        RECT 2.470 38.265 12.685 38.940 ;
        RECT 2.470 38.205 2.835 38.265 ;
        RECT 1.090 38.000 2.180 38.205 ;
        RECT 1.090 37.770 2.420 38.000 ;
        RECT 2.605 37.985 2.835 38.205 ;
        RECT 3.545 38.000 4.090 38.030 ;
        RECT 14.330 38.000 14.720 40.410 ;
        RECT 14.960 39.020 15.190 40.205 ;
        RECT 16.300 39.020 16.530 40.205 ;
        RECT 14.960 38.290 16.530 39.020 ;
        RECT 14.960 38.205 15.190 38.290 ;
        RECT 16.300 38.205 16.530 38.290 ;
        RECT 16.800 38.000 17.165 40.410 ;
        RECT 18.495 40.205 18.905 40.410 ;
        RECT 21.415 40.405 28.735 40.410 ;
        RECT 30.415 40.405 31.185 40.410 ;
        RECT 17.390 40.175 17.620 40.205 ;
        RECT 17.390 38.205 17.780 40.175 ;
        RECT 17.430 38.180 17.780 38.205 ;
        RECT 3.545 37.985 4.850 38.000 ;
        RECT 5.180 37.985 5.940 38.000 ;
        RECT 6.270 37.985 7.030 38.000 ;
        RECT 7.360 37.985 8.120 38.000 ;
        RECT 8.450 37.985 9.210 38.000 ;
        RECT 9.540 37.985 10.300 38.000 ;
        RECT 10.630 37.985 11.390 38.000 ;
        RECT 11.720 37.985 12.480 38.000 ;
        RECT 14.150 37.985 14.910 38.000 ;
        RECT 2.605 37.780 14.950 37.985 ;
        RECT 2.605 37.770 14.910 37.780 ;
        RECT 16.580 37.770 17.340 38.000 ;
        RECT 1.090 37.505 1.410 37.770 ;
        RECT 2.605 37.765 14.610 37.770 ;
        RECT 3.545 37.720 4.090 37.765 ;
        RECT 16.800 37.505 17.165 37.770 ;
        RECT 1.090 37.265 17.165 37.505 ;
        RECT 1.090 36.240 1.410 37.265 ;
        RECT 17.485 36.720 17.780 38.180 ;
        RECT 0.925 35.605 1.410 36.240 ;
        RECT 11.910 36.370 17.780 36.720 ;
        RECT 18.495 38.205 18.960 40.205 ;
        RECT 19.820 39.025 20.125 40.205 ;
        RECT 22.250 39.025 22.480 39.160 ;
        RECT 24.430 39.025 24.660 39.160 ;
        RECT 26.610 39.025 26.840 39.160 ;
        RECT 28.790 39.025 29.020 39.160 ;
        RECT 19.820 38.290 29.020 39.025 ;
        RECT 19.820 38.225 29.010 38.290 ;
        RECT 19.820 38.205 20.125 38.225 ;
        RECT 18.495 38.000 18.865 38.205 ;
        RECT 18.495 37.770 19.790 38.000 ;
        RECT 19.940 37.985 20.125 38.205 ;
        RECT 30.630 38.000 30.940 40.405 ;
        RECT 31.220 40.145 31.450 40.205 ;
        RECT 32.560 40.145 32.790 40.205 ;
        RECT 31.220 39.420 32.790 40.145 ;
        RECT 31.220 38.205 31.450 39.420 ;
        RECT 32.560 38.205 32.790 39.420 ;
        RECT 33.060 38.000 33.370 40.410 ;
        RECT 33.760 40.205 34.115 40.220 ;
        RECT 33.650 38.205 34.115 40.205 ;
        RECT 37.960 38.740 49.040 39.035 ;
        RECT 21.440 37.985 22.200 38.000 ;
        RECT 22.530 37.985 23.290 38.000 ;
        RECT 23.620 37.985 24.380 38.000 ;
        RECT 24.710 37.985 25.470 38.000 ;
        RECT 25.800 37.985 26.560 38.000 ;
        RECT 26.890 37.985 27.650 38.000 ;
        RECT 27.980 37.985 28.740 38.000 ;
        RECT 30.410 37.985 31.170 38.000 ;
        RECT 18.495 37.505 18.865 37.770 ;
        RECT 19.940 37.765 31.195 37.985 ;
        RECT 32.840 37.770 33.600 38.000 ;
        RECT 33.060 37.505 33.370 37.770 ;
        RECT 18.495 37.265 33.370 37.505 ;
        RECT 0.925 34.845 1.315 35.605 ;
        RECT 11.910 35.370 12.260 36.370 ;
        RECT 18.495 35.825 18.865 37.265 ;
        RECT 11.325 35.235 12.260 35.370 ;
        RECT 13.835 35.370 18.865 35.825 ;
        RECT 12.920 35.235 13.680 35.240 ;
        RECT 1.475 35.005 2.235 35.235 ;
        RECT 3.905 35.015 13.690 35.235 ;
        RECT 3.925 35.005 4.685 35.015 ;
        RECT 5.015 35.005 5.775 35.015 ;
        RECT 6.105 35.005 6.865 35.015 ;
        RECT 7.195 35.005 7.955 35.015 ;
        RECT 8.285 35.005 9.045 35.015 ;
        RECT 9.375 35.005 10.135 35.015 ;
        RECT 10.465 35.005 11.225 35.015 ;
        RECT 0.925 32.865 1.425 34.845 ;
        RECT 1.195 32.845 1.425 32.865 ;
        RECT 1.725 32.685 1.995 35.005 ;
        RECT 11.910 34.760 12.260 35.015 ;
        RECT 12.920 35.010 13.680 35.015 ;
        RECT 3.605 34.075 12.260 34.760 ;
        RECT 3.645 33.890 3.875 34.075 ;
        RECT 5.825 33.890 6.055 34.075 ;
        RECT 8.005 33.890 8.235 34.075 ;
        RECT 10.185 33.890 10.415 34.075 ;
        RECT 13.145 32.690 13.465 35.010 ;
        RECT 13.835 34.850 14.210 35.370 ;
        RECT 33.760 35.325 34.115 38.205 ;
        RECT 13.730 32.865 14.210 34.850 ;
        RECT 32.035 34.200 34.125 35.325 ;
        RECT 42.165 34.390 42.560 34.450 ;
        RECT 32.035 33.845 40.700 34.200 ;
        RECT 42.145 33.865 42.580 34.390 ;
        RECT 32.035 33.000 34.125 33.845 ;
        RECT 42.145 33.570 44.325 33.865 ;
        RECT 42.145 33.420 42.580 33.570 ;
        RECT 42.165 33.360 42.560 33.420 ;
        RECT 13.730 32.850 13.960 32.865 ;
        RECT 1.475 32.455 2.235 32.685 ;
        RECT 3.925 32.665 4.685 32.685 ;
        RECT 5.015 32.665 5.775 32.685 ;
        RECT 6.105 32.665 6.865 32.685 ;
        RECT 7.195 32.665 7.955 32.685 ;
        RECT 8.285 32.665 9.045 32.685 ;
        RECT 9.375 32.665 10.135 32.685 ;
        RECT 10.465 32.665 11.225 32.685 ;
        RECT 12.920 32.665 13.680 32.690 ;
        RECT 1.725 29.720 1.995 32.455 ;
        RECT 3.905 32.445 11.800 32.665 ;
        RECT 12.920 32.460 13.695 32.665 ;
        RECT 12.925 32.445 13.695 32.460 ;
        RECT 11.325 32.300 11.800 32.445 ;
        RECT 13.175 29.720 14.265 30.130 ;
        RECT 1.725 29.450 14.265 29.720 ;
        RECT 13.175 29.080 14.265 29.450 ;
      LAYER via ;
        RECT 3.595 40.410 4.005 40.720 ;
        RECT 3.595 37.720 4.005 38.030 ;
        RECT 41.695 38.740 42.595 39.035 ;
        RECT 11.375 35.015 11.755 35.370 ;
        RECT 32.160 33.115 34.015 35.180 ;
        RECT 42.195 33.420 42.530 34.390 ;
        RECT 11.375 32.300 11.750 32.665 ;
      LAYER met2 ;
        RECT 3.595 40.360 4.005 40.770 ;
        RECT 3.645 38.080 3.925 40.360 ;
        RECT 41.695 38.690 42.595 39.085 ;
        RECT 3.595 37.670 4.005 38.080 ;
        RECT 11.375 34.965 11.755 35.420 ;
        RECT 11.440 32.715 11.700 34.965 ;
        RECT 32.035 33.000 34.125 35.325 ;
        RECT 42.215 34.440 42.500 38.690 ;
        RECT 42.195 33.370 42.530 34.440 ;
        RECT 11.375 32.250 11.750 32.715 ;
      LAYER via2 ;
        RECT 32.160 33.115 34.015 35.180 ;
      LAYER met3 ;
        RECT 32.040 33.000 34.125 35.325 ;
      LAYER via3 ;
        RECT 32.160 33.115 34.015 35.180 ;
      LAYER met4 ;
        RECT 54.215 35.370 55.890 38.870 ;
        RECT 31.930 32.955 55.890 35.370 ;
        RECT 20.505 0.255 55.745 31.255 ;
      LAYER via4 ;
        RECT 54.395 33.075 55.730 38.775 ;
        RECT 54.465 0.460 55.645 31.050 ;
      LAYER met5 ;
        RECT 54.255 0.250 55.855 38.895 ;
  END
END simple_por
END LIBRARY

