magic
tech sky130A
timestamp 1724421276
use sky130_ef_sc_hd__fill_4  sky130_ef_sc_hd__fill_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1716601000
transform 1 0 0 0 1 0
box -19 -24 203 296
use sky130_ef_sc_hd__fill_8  sky130_ef_sc_hd__fill_8_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1716601000
transform 1 0 184 0 1 0
box -19 -24 387 296
<< end >>
