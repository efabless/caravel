* NGSPICE file created from housekeeping.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_2 abstract view
.subckt sky130_fd_sc_hd__ebufn_2 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_2 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtn_1 abstract view
.subckt sky130_fd_sc_hd__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4bb_1 abstract view
.subckt sky130_fd_sc_hd__nand4bb_1 A_N B_N C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

.subckt housekeeping VGND VPWR debug_in debug_mode debug_oeb debug_out irq[0] irq[1]
+ irq[2] mask_rev_in[0] mask_rev_in[10] mask_rev_in[11] mask_rev_in[12] mask_rev_in[13]
+ mask_rev_in[14] mask_rev_in[15] mask_rev_in[16] mask_rev_in[17] mask_rev_in[18]
+ mask_rev_in[19] mask_rev_in[1] mask_rev_in[20] mask_rev_in[21] mask_rev_in[22] mask_rev_in[23]
+ mask_rev_in[24] mask_rev_in[25] mask_rev_in[26] mask_rev_in[27] mask_rev_in[28]
+ mask_rev_in[29] mask_rev_in[2] mask_rev_in[30] mask_rev_in[31] mask_rev_in[3] mask_rev_in[4]
+ mask_rev_in[5] mask_rev_in[6] mask_rev_in[7] mask_rev_in[8] mask_rev_in[9] mgmt_gpio_in[0]
+ mgmt_gpio_in[10] mgmt_gpio_in[11] mgmt_gpio_in[12] mgmt_gpio_in[13] mgmt_gpio_in[14]
+ mgmt_gpio_in[15] mgmt_gpio_in[16] mgmt_gpio_in[17] mgmt_gpio_in[18] mgmt_gpio_in[19]
+ mgmt_gpio_in[1] mgmt_gpio_in[20] mgmt_gpio_in[21] mgmt_gpio_in[22] mgmt_gpio_in[23]
+ mgmt_gpio_in[24] mgmt_gpio_in[25] mgmt_gpio_in[26] mgmt_gpio_in[27] mgmt_gpio_in[28]
+ mgmt_gpio_in[29] mgmt_gpio_in[2] mgmt_gpio_in[30] mgmt_gpio_in[31] mgmt_gpio_in[32]
+ mgmt_gpio_in[33] mgmt_gpio_in[34] mgmt_gpio_in[35] mgmt_gpio_in[36] mgmt_gpio_in[37]
+ mgmt_gpio_in[3] mgmt_gpio_in[4] mgmt_gpio_in[5] mgmt_gpio_in[6] mgmt_gpio_in[7]
+ mgmt_gpio_in[8] mgmt_gpio_in[9] mgmt_gpio_oeb[0] mgmt_gpio_oeb[10] mgmt_gpio_oeb[11]
+ mgmt_gpio_oeb[12] mgmt_gpio_oeb[13] mgmt_gpio_oeb[14] mgmt_gpio_oeb[15] mgmt_gpio_oeb[16]
+ mgmt_gpio_oeb[17] mgmt_gpio_oeb[18] mgmt_gpio_oeb[19] mgmt_gpio_oeb[1] mgmt_gpio_oeb[20]
+ mgmt_gpio_oeb[21] mgmt_gpio_oeb[22] mgmt_gpio_oeb[23] mgmt_gpio_oeb[24] mgmt_gpio_oeb[25]
+ mgmt_gpio_oeb[26] mgmt_gpio_oeb[27] mgmt_gpio_oeb[28] mgmt_gpio_oeb[29] mgmt_gpio_oeb[2]
+ mgmt_gpio_oeb[30] mgmt_gpio_oeb[31] mgmt_gpio_oeb[32] mgmt_gpio_oeb[33] mgmt_gpio_oeb[34]
+ mgmt_gpio_oeb[35] mgmt_gpio_oeb[36] mgmt_gpio_oeb[37] mgmt_gpio_oeb[3] mgmt_gpio_oeb[4]
+ mgmt_gpio_oeb[5] mgmt_gpio_oeb[6] mgmt_gpio_oeb[7] mgmt_gpio_oeb[8] mgmt_gpio_oeb[9]
+ mgmt_gpio_out[0] mgmt_gpio_out[10] mgmt_gpio_out[11] mgmt_gpio_out[12] mgmt_gpio_out[13]
+ mgmt_gpio_out[14] mgmt_gpio_out[15] mgmt_gpio_out[16] mgmt_gpio_out[17] mgmt_gpio_out[18]
+ mgmt_gpio_out[19] mgmt_gpio_out[1] mgmt_gpio_out[20] mgmt_gpio_out[21] mgmt_gpio_out[22]
+ mgmt_gpio_out[23] mgmt_gpio_out[24] mgmt_gpio_out[25] mgmt_gpio_out[26] mgmt_gpio_out[27]
+ mgmt_gpio_out[28] mgmt_gpio_out[29] mgmt_gpio_out[2] mgmt_gpio_out[30] mgmt_gpio_out[31]
+ mgmt_gpio_out[32] mgmt_gpio_out[33] mgmt_gpio_out[34] mgmt_gpio_out[35] mgmt_gpio_out[36]
+ mgmt_gpio_out[37] mgmt_gpio_out[3] mgmt_gpio_out[4] mgmt_gpio_out[5] mgmt_gpio_out[6]
+ mgmt_gpio_out[7] mgmt_gpio_out[8] mgmt_gpio_out[9] pad_flash_clk pad_flash_clk_oeb
+ pad_flash_csb pad_flash_csb_oeb pad_flash_io0_di pad_flash_io0_do pad_flash_io0_ieb
+ pad_flash_io0_oeb pad_flash_io1_di pad_flash_io1_do pad_flash_io1_ieb pad_flash_io1_oeb
+ pll90_sel[0] pll90_sel[1] pll90_sel[2] pll_bypass pll_dco_ena pll_div[0] pll_div[1]
+ pll_div[2] pll_div[3] pll_div[4] pll_ena pll_sel[0] pll_sel[1] pll_sel[2] pll_trim[0]
+ pll_trim[10] pll_trim[11] pll_trim[12] pll_trim[13] pll_trim[14] pll_trim[15] pll_trim[16]
+ pll_trim[17] pll_trim[18] pll_trim[19] pll_trim[1] pll_trim[20] pll_trim[21] pll_trim[22]
+ pll_trim[23] pll_trim[24] pll_trim[25] pll_trim[2] pll_trim[3] pll_trim[4] pll_trim[5]
+ pll_trim[6] pll_trim[7] pll_trim[8] pll_trim[9] porb pwr_ctrl_out[0] pwr_ctrl_out[1]
+ pwr_ctrl_out[2] pwr_ctrl_out[3] qspi_enabled reset ser_rx ser_tx serial_clock serial_data_1
+ serial_data_2 serial_load serial_resetn spi_csb spi_enabled spi_sck spi_sdi spi_sdo
+ spi_sdoenb spimemio_flash_clk spimemio_flash_csb spimemio_flash_io0_di spimemio_flash_io0_do
+ spimemio_flash_io0_oeb spimemio_flash_io1_di spimemio_flash_io1_do spimemio_flash_io1_oeb
+ spimemio_flash_io2_di spimemio_flash_io2_do spimemio_flash_io2_oeb spimemio_flash_io3_di
+ spimemio_flash_io3_do spimemio_flash_io3_oeb sram_ro_addr[0] sram_ro_addr[1] sram_ro_addr[2]
+ sram_ro_addr[3] sram_ro_addr[4] sram_ro_addr[5] sram_ro_addr[6] sram_ro_addr[7]
+ sram_ro_clk sram_ro_csb sram_ro_data[0] sram_ro_data[10] sram_ro_data[11] sram_ro_data[12]
+ sram_ro_data[13] sram_ro_data[14] sram_ro_data[15] sram_ro_data[16] sram_ro_data[17]
+ sram_ro_data[18] sram_ro_data[19] sram_ro_data[1] sram_ro_data[20] sram_ro_data[21]
+ sram_ro_data[22] sram_ro_data[23] sram_ro_data[24] sram_ro_data[25] sram_ro_data[26]
+ sram_ro_data[27] sram_ro_data[28] sram_ro_data[29] sram_ro_data[2] sram_ro_data[30]
+ sram_ro_data[31] sram_ro_data[3] sram_ro_data[4] sram_ro_data[5] sram_ro_data[6]
+ sram_ro_data[7] sram_ro_data[8] sram_ro_data[9] trap uart_enabled user_clock usr1_vcc_pwrgood
+ usr1_vdd_pwrgood usr2_vcc_pwrgood usr2_vdd_pwrgood wb_ack_o wb_adr_i[0] wb_adr_i[10]
+ wb_adr_i[11] wb_adr_i[12] wb_adr_i[13] wb_adr_i[14] wb_adr_i[15] wb_adr_i[16] wb_adr_i[17]
+ wb_adr_i[18] wb_adr_i[19] wb_adr_i[1] wb_adr_i[20] wb_adr_i[21] wb_adr_i[22] wb_adr_i[23]
+ wb_adr_i[24] wb_adr_i[25] wb_adr_i[26] wb_adr_i[27] wb_adr_i[28] wb_adr_i[29] wb_adr_i[2]
+ wb_adr_i[30] wb_adr_i[31] wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6] wb_adr_i[7]
+ wb_adr_i[8] wb_adr_i[9] wb_clk_i wb_cyc_i wb_dat_i[0] wb_dat_i[10] wb_dat_i[11]
+ wb_dat_i[12] wb_dat_i[13] wb_dat_i[14] wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18]
+ wb_dat_i[19] wb_dat_i[1] wb_dat_i[20] wb_dat_i[21] wb_dat_i[22] wb_dat_i[23] wb_dat_i[24]
+ wb_dat_i[25] wb_dat_i[26] wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[2] wb_dat_i[30]
+ wb_dat_i[31] wb_dat_i[3] wb_dat_i[4] wb_dat_i[5] wb_dat_i[6] wb_dat_i[7] wb_dat_i[8]
+ wb_dat_i[9] wb_dat_o[0] wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13] wb_dat_o[14]
+ wb_dat_o[15] wb_dat_o[16] wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[1] wb_dat_o[20]
+ wb_dat_o[21] wb_dat_o[22] wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26] wb_dat_o[27]
+ wb_dat_o[28] wb_dat_o[29] wb_dat_o[2] wb_dat_o[30] wb_dat_o[31] wb_dat_o[3] wb_dat_o[4]
+ wb_dat_o[5] wb_dat_o[6] wb_dat_o[7] wb_dat_o[8] wb_dat_o[9] wb_rstn_i wb_sel_i[0]
+ wb_sel_i[1] wb_sel_i[2] wb_sel_i[3] wb_stb_i wb_we_i
XFILLER_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7963_ _7979_/A _7994_/B VGND VGND VPWR VPWR _8096_/B sky130_fd_sc_hd__or2_4
XFILLER_82_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9702_ _4446_/A1 _9702_/D _4981_/X VGND VGND VPWR VPWR _9702_/Q sky130_fd_sc_hd__dfrtp_1
X_6914_ _9287_/Q VGND VGND VPWR VPWR _6914_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_82_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7894_ _8583_/A _7894_/B _7903_/C _8193_/A VGND VGND VPWR VPWR _7895_/A sky130_fd_sc_hd__or4_1
XFILLER_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9633_ _9639_/CLK _9633_/D _9633_/SET_B VGND VGND VPWR VPWR _9633_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_22_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6845_ _9537_/Q VGND VGND VPWR VPWR _6845_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9564_ _9617_/CLK _9564_/D _9295_/SET_B VGND VGND VPWR VPWR _9564_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6776_ _6774_/Y _5121_/B _6775_/Y _5949_/B VGND VGND VPWR VPWR _6776_/X sky130_fd_sc_hd__o22a_1
X_8515_ _8515_/A _8515_/B VGND VGND VPWR VPWR _8703_/B sky130_fd_sc_hd__nor2_1
X_9495_ _9534_/CLK _9495_/D _9647_/SET_B VGND VGND VPWR VPWR _9495_/Q sky130_fd_sc_hd__dfstp_1
X_5727_ _7041_/A _7127_/C VGND VGND VPWR VPWR _5728_/A sky130_fd_sc_hd__or2_1
X_8446_ _7864_/X _8341_/B _8009_/X _8445_/X _8013_/X VGND VGND VPWR VPWR _8448_/C
+ sky130_fd_sc_hd__o2111ai_2
XFILLER_108_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5658_ _5658_/A VGND VGND VPWR VPWR _5658_/Y sky130_fd_sc_hd__inv_2
X_8377_ _8583_/C _8377_/B _8377_/C VGND VGND VPWR VPWR _8565_/A sky130_fd_sc_hd__or3_1
XFILLER_151_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5589_ _9316_/Q _5585_/A _8925_/A1 _5585_/Y VGND VGND VPWR VPWR _9316_/D sky130_fd_sc_hd__a22o_1
X_4609_ _9727_/Q _4604_/A _5966_/B1 _4604_/Y VGND VGND VPWR VPWR _9727_/D sky130_fd_sc_hd__a22o_1
XFILLER_104_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7328_ _6812_/Y _7126_/X _6868_/Y _7128_/X VGND VGND VPWR VPWR _7328_/X sky130_fd_sc_hd__o22a_1
XFILLER_117_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7259_ _6218_/Y _7059_/D _6152_/Y _7116_/X _7258_/X VGND VGND VPWR VPWR _7264_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_131_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4960_ _6022_/A _6022_/B _6022_/C _9708_/Q VGND VGND VPWR VPWR _4960_/X sky130_fd_sc_hd__o31a_1
X_4891_ _4891_/A _4911_/A VGND VGND VPWR VPWR _5450_/B sky130_fd_sc_hd__or2_4
X_6630_ _6149_/A _6629_/Y _9039_/Q _6149_/Y VGND VGND VPWR VPWR _9039_/D sky130_fd_sc_hd__o22a_1
XFILLER_20_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6561_ _6561_/A VGND VGND VPWR VPWR _6561_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_164_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5512_ _9369_/Q _5509_/A _8844_/X _5509_/Y VGND VGND VPWR VPWR _9369_/D sky130_fd_sc_hd__a22o_1
X_8300_ _8496_/A _8300_/B VGND VGND VPWR VPWR _8301_/A sky130_fd_sc_hd__or2_1
XFILLER_118_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6492_ _9207_/Q VGND VGND VPWR VPWR _8751_/A sky130_fd_sc_hd__inv_6
XFILLER_145_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9280_ _9280_/CLK _9280_/D _9757_/SET_B VGND VGND VPWR VPWR _9280_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_172_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5443_ _5443_/A VGND VGND VPWR VPWR _5444_/A sky130_fd_sc_hd__clkbuf_2
X_8231_ _8231_/A _8676_/B _8658_/B _8573_/B VGND VGND VPWR VPWR _8237_/A sky130_fd_sc_hd__or4_1
X_5374_ _5671_/A _5374_/B VGND VGND VPWR VPWR _5375_/A sky130_fd_sc_hd__or2_1
XFILLER_99_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8162_ _8162_/A _8370_/A VGND VGND VPWR VPWR _8163_/B sky130_fd_sc_hd__or2_1
X_7113_ _4742_/Y _7112_/X _4668_/Y _7077_/B VGND VGND VPWR VPWR _7113_/X sky130_fd_sc_hd__o22a_1
X_8093_ _8093_/A _8093_/B VGND VGND VPWR VPWR _8431_/A sky130_fd_sc_hd__nor2_1
XFILLER_141_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7044_ _7075_/A _7115_/B VGND VGND VPWR VPWR _7045_/A sky130_fd_sc_hd__or2_1
XFILLER_82_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8995_ _9563_/Q _8767_/A VGND VGND VPWR VPWR mgmt_gpio_out[18] sky130_fd_sc_hd__ebufn_8
XFILLER_103_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7946_ _8379_/C _8195_/A VGND VGND VPWR VPWR _8079_/C sky130_fd_sc_hd__or2_1
XFILLER_82_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7877_ _8515_/B _8232_/B VGND VGND VPWR VPWR _7877_/X sky130_fd_sc_hd__or2_2
X_9616_ _9788_/CLK _9616_/D _9646_/SET_B VGND VGND VPWR VPWR _9616_/Q sky130_fd_sc_hd__dfrtp_1
X_6828_ _6823_/Y _6027_/B _6824_/Y _5336_/B _6827_/X VGND VGND VPWR VPWR _6829_/D
+ sky130_fd_sc_hd__o221a_2
XFILLER_50_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6759_ _6759_/A _6759_/B _6759_/C VGND VGND VPWR VPWR _6784_/C sky130_fd_sc_hd__and3_1
X_9547_ _9639_/CLK _9547_/D _9757_/SET_B VGND VGND VPWR VPWR _9547_/Q sky130_fd_sc_hd__dfstp_1
X_9478_ _9483_/CLK _9478_/D _9685_/SET_B VGND VGND VPWR VPWR _9478_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_148_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8429_ _8703_/A _8585_/B VGND VGND VPWR VPWR _8560_/B sky130_fd_sc_hd__or2_1
XFILLER_163_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5090_ _5090_/A VGND VGND VPWR VPWR _5091_/A sky130_fd_sc_hd__buf_2
XFILLER_96_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8780_ _8780_/A VGND VGND VPWR VPWR _8780_/X sky130_fd_sc_hd__clkbuf_1
X_7800_ _8379_/C _7839_/A _8379_/D VGND VGND VPWR VPWR _8093_/A sky130_fd_sc_hd__or3_4
X_5992_ _9698_/Q _5992_/B VGND VGND VPWR VPWR _7008_/B sky130_fd_sc_hd__nand2_1
X_7731_ _7731_/A _8975_/S VGND VGND VPWR VPWR _7732_/A sky130_fd_sc_hd__and2_1
X_4943_ _6022_/A _6022_/D _6022_/C VGND VGND VPWR VPWR _4944_/A sky130_fd_sc_hd__or3_1
XFILLER_24_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7662_ _7662_/A _7662_/B _7662_/C _7662_/D VGND VGND VPWR VPWR _7662_/Y sky130_fd_sc_hd__nand4_4
X_6613_ _8771_/A _5420_/B _6612_/Y _5442_/B VGND VGND VPWR VPWR _6613_/X sky130_fd_sc_hd__o22a_1
X_9401_ _9758_/CLK _9401_/D _7011_/B VGND VGND VPWR VPWR _9401_/Q sky130_fd_sc_hd__dfrtp_2
X_4874_ _9726_/Q VGND VGND VPWR VPWR _4874_/Y sky130_fd_sc_hd__inv_2
X_7593_ _6129_/Y _7419_/X _6116_/Y _7421_/X VGND VGND VPWR VPWR _7593_/X sky130_fd_sc_hd__o22a_1
XFILLER_20_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6544_ _9635_/Q VGND VGND VPWR VPWR _6544_/Y sky130_fd_sc_hd__clkinv_2
X_9332_ _9545_/CLK _9332_/D _4628_/A VGND VGND VPWR VPWR _9332_/Q sky130_fd_sc_hd__dfstp_1
X_9263_ _9601_/CLK _9263_/D _9295_/SET_B VGND VGND VPWR VPWR _9263_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_165_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6475_ _6475_/A _6475_/B _6475_/C _6475_/D VGND VGND VPWR VPWR _6475_/Y sky130_fd_sc_hd__nand4_2
X_8214_ _8311_/B VGND VGND VPWR VPWR _8214_/Y sky130_fd_sc_hd__inv_2
XFILLER_161_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5426_ _9428_/Q _5422_/A _8925_/A1 _5422_/Y VGND VGND VPWR VPWR _9428_/D sky130_fd_sc_hd__a22o_1
Xoutput231 _8792_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[30] sky130_fd_sc_hd__buf_2
Xoutput220 _8772_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[20] sky130_fd_sc_hd__buf_2
XFILLER_160_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9194_ _9378_/CLK _9194_/D _9646_/SET_B VGND VGND VPWR VPWR _9194_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput242 _7702_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[6] sky130_fd_sc_hd__buf_2
Xoutput253 _8836_/X VGND VGND VPWR VPWR pad_flash_csb sky130_fd_sc_hd__buf_2
X_5357_ _5357_/A VGND VGND VPWR VPWR _5357_/Y sky130_fd_sc_hd__clkinv_2
X_8145_ _7987_/Y _8390_/B _8144_/X VGND VGND VPWR VPWR _8145_/X sky130_fd_sc_hd__a21o_1
Xoutput286 _9733_/Q VGND VGND VPWR VPWR pll_trim[1] sky130_fd_sc_hd__buf_2
Xoutput275 _9732_/Q VGND VGND VPWR VPWR pll_trim[0] sky130_fd_sc_hd__buf_2
Xoutput264 _9758_/Q VGND VGND VPWR VPWR pll_bypass sky130_fd_sc_hd__buf_2
X_5288_ _9520_/Q _5280_/A _8916_/A1 _5280_/Y VGND VGND VPWR VPWR _9520_/D sky130_fd_sc_hd__a22o_1
X_8076_ _8515_/B _8437_/B _8075_/Y VGND VGND VPWR VPWR _8078_/A sky130_fd_sc_hd__o21ai_1
Xoutput297 _9738_/Q VGND VGND VPWR VPWR pll_trim[6] sky130_fd_sc_hd__buf_2
XFILLER_87_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7027_ _7027_/A VGND VGND VPWR VPWR _7073_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8978_ _7482_/X _4875_/Y _8978_/S VGND VGND VPWR VPWR _8978_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7929_ _7929_/A _7929_/B VGND VGND VPWR VPWR _7929_/Y sky130_fd_sc_hd__nand2_1
XFILLER_43_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xnet299_3 _8837_/A1 VGND VGND VPWR VPWR _6359_/A1 sky130_fd_sc_hd__inv_4
XFILLER_187_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4590_ _5960_/A _4590_/B VGND VGND VPWR VPWR _4591_/A sky130_fd_sc_hd__or2_1
XFILLER_155_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6260_ _6258_/Y _4590_/B _6259_/Y _6086_/X VGND VGND VPWR VPWR _6260_/X sky130_fd_sc_hd__o22a_1
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6191_ input41/X _8930_/S _6190_/Y _5431_/B VGND VGND VPWR VPWR _6191_/X sky130_fd_sc_hd__o2bb2a_1
X_5211_ _9570_/Q _5203_/Y _8916_/X _5203_/A VGND VGND VPWR VPWR _9570_/D sky130_fd_sc_hd__o22a_1
XFILLER_130_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5142_ _9620_/Q _5136_/A _8955_/A1 _5136_/Y VGND VGND VPWR VPWR _9620_/D sky130_fd_sc_hd__a22o_1
XFILLER_96_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5073_ _5073_/A VGND VGND VPWR VPWR _9662_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8901_ _7728_/X _9698_/Q _9048_/Q VGND VGND VPWR VPWR _8901_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8832_ _6544_/Y _9058_/Q _8977_/S VGND VGND VPWR VPWR _8832_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8763_ _8763_/A VGND VGND VPWR VPWR _8764_/A sky130_fd_sc_hd__clkbuf_1
X_5975_ _9096_/Q _5970_/A _8929_/A1 _5970_/Y VGND VGND VPWR VPWR _9096_/D sky130_fd_sc_hd__a22o_1
XFILLER_12_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4926_ _9502_/Q VGND VGND VPWR VPWR _4926_/Y sky130_fd_sc_hd__clkinv_4
X_8694_ _8496_/A _8216_/X _8312_/D _7905_/X VGND VGND VPWR VPWR _8695_/B sky130_fd_sc_hd__o211ai_1
X_7714_ _9084_/Q _7713_/B _9085_/Q VGND VGND VPWR VPWR _7715_/B sky130_fd_sc_hd__a21oi_1
X_7645_ _6729_/Y _7408_/X _6685_/Y _7410_/X VGND VGND VPWR VPWR _7645_/X sky130_fd_sc_hd__o22a_1
X_4857_ _9778_/Q VGND VGND VPWR VPWR _4857_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7576_ _6182_/Y _7415_/X _6215_/Y _7417_/X _7575_/X VGND VGND VPWR VPWR _7590_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6527_ _9367_/Q VGND VGND VPWR VPWR _8799_/A sky130_fd_sc_hd__inv_6
XFILLER_146_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9315_ _9535_/CLK _9315_/D _9647_/SET_B VGND VGND VPWR VPWR _9315_/Q sky130_fd_sc_hd__dfrtp_1
X_4788_ _4784_/Y _5941_/B _4786_/Y _5488_/B VGND VGND VPWR VPWR _4788_/X sky130_fd_sc_hd__o22a_2
XFILLER_134_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6458_ _9105_/Q VGND VGND VPWR VPWR _6458_/Y sky130_fd_sc_hd__clkinv_4
X_9246_ _9279_/CLK _9246_/D _9779_/SET_B VGND VGND VPWR VPWR _9246_/Q sky130_fd_sc_hd__dfstp_2
X_9177_ _9613_/CLK _9177_/D _9646_/SET_B VGND VGND VPWR VPWR _9177_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_121_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5409_ _9439_/Q _5406_/A _5965_/B1 _5406_/Y VGND VGND VPWR VPWR _9439_/D sky130_fd_sc_hd__a22o_1
X_6389_ _6384_/Y _4564_/B _6385_/Y _4907_/X _6388_/X VGND VGND VPWR VPWR _6408_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_161_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8128_ _8130_/B _8640_/B VGND VGND VPWR VPWR _8676_/A sky130_fd_sc_hd__nor2_1
XFILLER_125_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8059_ _8085_/A VGND VGND VPWR VPWR _8064_/B sky130_fd_sc_hd__inv_2
XFILLER_87_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5760_ _9238_/Q _5759_/A _8846_/X _5759_/Y VGND VGND VPWR VPWR _9238_/D sky130_fd_sc_hd__a22o_1
XFILLER_187_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4711_ _4931_/A _4780_/B VGND VGND VPWR VPWR _5632_/B sky130_fd_sc_hd__or2_4
XFILLER_91_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5691_ _5691_/A _9055_/Q VGND VGND VPWR VPWR _5692_/A sky130_fd_sc_hd__or2_2
XFILLER_175_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4642_ _4642_/A VGND VGND VPWR VPWR _4642_/X sky130_fd_sc_hd__clkbuf_1
X_7430_ _7430_/A VGND VGND VPWR VPWR _7430_/X sky130_fd_sc_hd__buf_6
XFILLER_175_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7361_ _6577_/Y _7079_/B _6510_/Y _7059_/A VGND VGND VPWR VPWR _7361_/X sky130_fd_sc_hd__o22a_1
X_4573_ _9749_/Q _4566_/A _5966_/B1 _4566_/Y VGND VGND VPWR VPWR _9749_/D sky130_fd_sc_hd__a22o_1
X_9100_ _9652_/CLK _9100_/D _9647_/SET_B VGND VGND VPWR VPWR _9100_/Q sky130_fd_sc_hd__dfrtp_1
X_6312_ _6310_/Y _6081_/B _6311_/Y _5583_/B VGND VGND VPWR VPWR _6312_/X sky130_fd_sc_hd__o22a_1
X_7292_ _4761_/Y _7048_/B _4784_/Y _7077_/A _7291_/X VGND VGND VPWR VPWR _7299_/A
+ sky130_fd_sc_hd__o221a_1
X_9031_ _9039_/CLK _9031_/D VGND VGND VPWR VPWR _9031_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6243_ _9745_/Q VGND VGND VPWR VPWR _6243_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6174_ _6174_/A _6174_/B _6174_/C _6174_/D VGND VGND VPWR VPWR _6237_/A sky130_fd_sc_hd__and4_1
X_5125_ _9630_/Q _5123_/A _5964_/B1 _5123_/Y VGND VGND VPWR VPWR _9630_/D sky130_fd_sc_hd__a22o_1
X_5056_ _7733_/A _7734_/A _8810_/A VGND VGND VPWR VPWR _5062_/A sky130_fd_sc_hd__a21oi_1
XFILLER_84_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_1_wb_clk_i clkbuf_1_0_1_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_2_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_52_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5958_ _9107_/Q _5951_/A _8930_/A1 _5951_/Y VGND VGND VPWR VPWR _9107_/D sky130_fd_sc_hd__a22o_1
X_8746_ _8746_/A VGND VGND VPWR VPWR _8746_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4909_ _9758_/Q VGND VGND VPWR VPWR _4909_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8677_ _8677_/A _8677_/B _8677_/C _8677_/D VGND VGND VPWR VPWR _8731_/D sky130_fd_sc_hd__or4_4
X_5889_ _5849_/A _8885_/X _8924_/X _9144_/Q VGND VGND VPWR VPWR _9144_/D sky130_fd_sc_hd__o22a_1
XFILLER_21_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7628_ _6801_/Y _7400_/X _6927_/Y _7405_/X _7627_/X VGND VGND VPWR VPWR _7644_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_193_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7559_ _6246_/Y _7427_/X _6320_/Y _5699_/X VGND VGND VPWR VPWR _7559_/X sky130_fd_sc_hd__o22a_1
XFILLER_20_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_2_0_csclk clkbuf_2_3_0_csclk/A VGND VGND VPWR VPWR clkbuf_2_2_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_134_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9229_ _9440_/CLK _9229_/D _9685_/SET_B VGND VGND VPWR VPWR _9229_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_5 _7243_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6930_ _6928_/Y _5671_/B _6929_/Y _5960_/B VGND VGND VPWR VPWR _6930_/X sky130_fd_sc_hd__o22a_1
XFILLER_66_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_6_csclk clkbuf_leaf_6_csclk/A VGND VGND VPWR VPWR _9440_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_81_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6861_ _9741_/Q VGND VGND VPWR VPWR _6861_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8600_ _8600_/A _8600_/B VGND VGND VPWR VPWR _8662_/C sky130_fd_sc_hd__or2_1
X_5812_ _5812_/A VGND VGND VPWR VPWR _5812_/Y sky130_fd_sc_hd__inv_2
X_6792_ _6787_/Y _5355_/B _6788_/Y _5267_/B _6791_/X VGND VGND VPWR VPWR _6830_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_62_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9580_ _9620_/CLK _9580_/D _9633_/SET_B VGND VGND VPWR VPWR _9580_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5743_ _5743_/A VGND VGND VPWR VPWR _5744_/A sky130_fd_sc_hd__clkbuf_2
X_8531_ _8607_/A _8531_/B _8734_/D _8614_/D VGND VGND VPWR VPWR _8535_/A sky130_fd_sc_hd__or4_1
Xclkbuf_1_0_0_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR clkbuf_1_0_1_mgmt_gpio_in[4]/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_22_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5674_ _9268_/Q _5673_/A _8843_/X _5673_/Y VGND VGND VPWR VPWR _9268_/D sky130_fd_sc_hd__a22o_1
X_8462_ _7836_/B _8299_/B _7862_/Y _8544_/A _7987_/Y VGND VGND VPWR VPWR _8668_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_148_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8393_ _8393_/A VGND VGND VPWR VPWR _8393_/Y sky130_fd_sc_hd__inv_2
X_4625_ _4625_/A VGND VGND VPWR VPWR _9720_/D sky130_fd_sc_hd__clkbuf_1
X_7413_ _7413_/A _9253_/Q VGND VGND VPWR VPWR _7474_/C sky130_fd_sc_hd__or2_4
X_7344_ _6632_/Y _7112_/X _6750_/Y _7077_/B VGND VGND VPWR VPWR _7344_/X sky130_fd_sc_hd__o22a_1
X_4556_ _4556_/A VGND VGND VPWR VPWR _9758_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7275_ _6126_/Y _7068_/A _6083_/Y _7105_/X VGND VGND VPWR VPWR _7275_/X sky130_fd_sc_hd__o22a_1
X_4487_ _4661_/C _8938_/X _4801_/C VGND VGND VPWR VPWR _4488_/A sky130_fd_sc_hd__or3_1
X_9014_ _9027_/CLK _9014_/D VGND VGND VPWR VPWR _9014_/Q sky130_fd_sc_hd__dfxtp_1
X_6226_ _9768_/Q VGND VGND VPWR VPWR _6226_/Y sky130_fd_sc_hd__clkinv_2
X_6157_ _9652_/Q VGND VGND VPWR VPWR _6157_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5108_ _9061_/Q _9062_/Q _9063_/Q _9065_/D VGND VGND VPWR VPWR _5108_/X sky130_fd_sc_hd__or4_2
XFILLER_106_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater361 _8843_/X VGND VGND VPWR VPWR _8925_/A1 sky130_fd_sc_hd__buf_12
Xrepeater372 _9647_/SET_B VGND VGND VPWR VPWR _9295_/SET_B sky130_fd_sc_hd__buf_12
X_6088_ _6085_/Y _6086_/X _6087_/Y _4870_/X VGND VGND VPWR VPWR _6088_/X sky130_fd_sc_hd__o22a_1
XFILLER_38_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5039_ _8974_/X _4551_/B _9680_/Q _5062_/D VGND VGND VPWR VPWR _9680_/D sky130_fd_sc_hd__a22o_1
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9778_ _9785_/CLK _9778_/D _9779_/SET_B VGND VGND VPWR VPWR _9778_/Q sky130_fd_sc_hd__dfstp_1
X_8729_ _8729_/A VGND VGND VPWR VPWR _8729_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput120 sram_ro_data[5] VGND VGND VPWR VPWR _6270_/A sky130_fd_sc_hd__clkbuf_1
Xinput131 usr2_vdd_pwrgood VGND VGND VPWR VPWR _4867_/A sky130_fd_sc_hd__clkbuf_1
Xinput153 wb_adr_i[29] VGND VGND VPWR VPWR input153/X sky130_fd_sc_hd__clkbuf_1
Xinput142 wb_adr_i[19] VGND VGND VPWR VPWR _7768_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_163_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput164 wb_cyc_i VGND VGND VPWR VPWR input164/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput186 wb_dat_i[29] VGND VGND VPWR VPWR _7747_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput175 wb_dat_i[19] VGND VGND VPWR VPWR _7742_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_76_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput197 wb_rstn_i VGND VGND VPWR VPWR _6146_/A sky130_fd_sc_hd__buf_12
XFILLER_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5390_ _9452_/Q _5384_/A _8841_/X _5384_/Y VGND VGND VPWR VPWR _9452_/D sky130_fd_sc_hd__a22o_1
XFILLER_172_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7060_ _7104_/A _7127_/B _7073_/C VGND VGND VPWR VPWR _7061_/A sky130_fd_sc_hd__or3_1
XFILLER_140_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6011_ _9084_/Q _5995_/A _8899_/X _5995_/Y VGND VGND VPWR VPWR _9084_/D sky130_fd_sc_hd__a22o_1
XFILLER_140_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7962_ _8528_/A _7960_/Y _8193_/A _8193_/B VGND VGND VPWR VPWR _7994_/B sky130_fd_sc_hd__o22a_1
X_9701_ _4446_/A1 _9701_/D _4984_/X VGND VGND VPWR VPWR _9701_/Q sky130_fd_sc_hd__dfrtp_1
X_6913_ _9094_/Q VGND VGND VPWR VPWR _6913_/Y sky130_fd_sc_hd__clkinv_2
X_7893_ _8077_/A _8232_/B _8441_/A _7892_/X VGND VGND VPWR VPWR _7893_/X sky130_fd_sc_hd__o211a_1
X_9632_ _9639_/CLK _9632_/D _9633_/SET_B VGND VGND VPWR VPWR _9632_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_22_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6844_ _9779_/Q VGND VGND VPWR VPWR _6844_/Y sky130_fd_sc_hd__inv_2
X_9563_ _9617_/CLK _9563_/D _9295_/SET_B VGND VGND VPWR VPWR _9563_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6775_ _9108_/Q VGND VGND VPWR VPWR _6775_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8514_ _8514_/A _8514_/B _8514_/C VGND VGND VPWR VPWR _8605_/B sky130_fd_sc_hd__or3_1
X_9494_ _9534_/CLK _9494_/D _9647_/SET_B VGND VGND VPWR VPWR _9494_/Q sky130_fd_sc_hd__dfstp_1
X_5726_ _5726_/A VGND VGND VPWR VPWR _7127_/C sky130_fd_sc_hd__buf_4
X_8445_ _8272_/A _8521_/B _8164_/A _8525_/C _8085_/A VGND VGND VPWR VPWR _8445_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_184_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5657_ _9054_/Q _9056_/Q _5724_/B _5647_/X _5656_/Y VGND VGND VPWR VPWR _9278_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_184_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8376_ _8376_/A _8539_/A VGND VGND VPWR VPWR _8380_/B sky130_fd_sc_hd__or2_1
X_5588_ _9317_/Q _5585_/A _8844_/X _5585_/Y VGND VGND VPWR VPWR _9317_/D sky130_fd_sc_hd__a22o_1
XFILLER_2_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4608_ _9728_/Q _4604_/A _5965_/B1 _4604_/Y VGND VGND VPWR VPWR _9728_/D sky130_fd_sc_hd__a22o_1
XFILLER_190_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7327_ _6856_/Y _5728_/X _6902_/Y _7040_/A _7326_/X VGND VGND VPWR VPWR _7330_/C
+ sky130_fd_sc_hd__o221a_2
XFILLER_104_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4539_ _4539_/A VGND VGND VPWR VPWR _9761_/D sky130_fd_sc_hd__clkbuf_1
X_7258_ _6171_/Y _7118_/X _6205_/Y _7048_/C VGND VGND VPWR VPWR _7258_/X sky130_fd_sc_hd__o22a_1
XFILLER_131_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6209_ _6207_/Y _4822_/X _6208_/Y _4907_/X VGND VGND VPWR VPWR _6209_/X sky130_fd_sc_hd__o22a_1
X_7189_ _7189_/A _7189_/B _7189_/C _7189_/D VGND VGND VPWR VPWR _7199_/B sky130_fd_sc_hd__and4_1
XFILLER_58_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4890_ _9406_/Q VGND VGND VPWR VPWR _4890_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6560_ _6555_/Y _5518_/B _6556_/Y _5404_/B _6559_/X VGND VGND VPWR VPWR _6567_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_192_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5511_ _9370_/Q _5509_/A _8845_/X _5509_/Y VGND VGND VPWR VPWR _9370_/D sky130_fd_sc_hd__a22o_1
X_6491_ _9341_/Q VGND VGND VPWR VPWR _6491_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5442_ _5671_/A _5442_/B VGND VGND VPWR VPWR _5443_/A sky130_fd_sc_hd__or2_1
X_8230_ _8230_/A _8260_/B VGND VGND VPWR VPWR _8573_/B sky130_fd_sc_hd__nor2_1
XFILLER_8_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8161_ _8554_/A _8378_/B VGND VGND VPWR VPWR _8370_/A sky130_fd_sc_hd__nor2_1
X_5373_ _9463_/Q _5368_/A _5967_/B1 _5368_/Y VGND VGND VPWR VPWR _9463_/D sky130_fd_sc_hd__a22o_1
XFILLER_172_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_24_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR _9788_/CLK sky130_fd_sc_hd__clkbuf_16
X_8092_ _8093_/B VGND VGND VPWR VPWR _8092_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7112_ _7112_/A VGND VGND VPWR VPWR _7112_/X sky130_fd_sc_hd__buf_8
XFILLER_141_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7043_ _7043_/A VGND VGND VPWR VPWR _7048_/B sky130_fd_sc_hd__buf_8
XFILLER_67_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_39_csclk clkbuf_2_1_0_csclk/X VGND VGND VPWR VPWR _9655_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_67_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8994_ _9562_/Q _8765_/A VGND VGND VPWR VPWR mgmt_gpio_out[17] sky130_fd_sc_hd__ebufn_8
XFILLER_82_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7945_ _8077_/A _8188_/B _9068_/Q VGND VGND VPWR VPWR _8514_/B sky130_fd_sc_hd__o21ai_1
XFILLER_103_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7876_ _8226_/C _8230_/A VGND VGND VPWR VPWR _8232_/B sky130_fd_sc_hd__or2_2
XFILLER_23_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9615_ _9788_/CLK _9615_/D _9646_/SET_B VGND VGND VPWR VPWR _9615_/Q sky130_fd_sc_hd__dfrtp_1
X_6827_ _6825_/Y _5317_/B _6826_/Y _5412_/B VGND VGND VPWR VPWR _6827_/X sky130_fd_sc_hd__o22a_1
X_9546_ _9757_/CLK _9546_/D _9757_/SET_B VGND VGND VPWR VPWR _9546_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_50_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6758_ _6753_/Y _6081_/B _6754_/Y _5905_/B _6757_/X VGND VGND VPWR VPWR _6759_/C
+ sky130_fd_sc_hd__o221a_1
X_9477_ _9527_/CLK _9477_/D _9685_/SET_B VGND VGND VPWR VPWR _9477_/Q sky130_fd_sc_hd__dfstp_1
X_6689_ _6685_/Y _5024_/B _6686_/Y _5507_/B _6688_/X VGND VGND VPWR VPWR _6690_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_12_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5709_ _7476_/A _7401_/B VGND VGND VPWR VPWR _7472_/A sky130_fd_sc_hd__or2_4
XFILLER_148_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8428_ _8687_/B _8428_/B VGND VGND VPWR VPWR _8430_/A sky130_fd_sc_hd__or2_1
XFILLER_109_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8359_ _8359_/A _8359_/B VGND VGND VPWR VPWR _8574_/C sky130_fd_sc_hd__or2_1
XFILLER_151_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5991_ _5991_/A VGND VGND VPWR VPWR _5991_/X sky130_fd_sc_hd__clkbuf_1
X_4942_ _9090_/Q VGND VGND VPWR VPWR _6022_/C sky130_fd_sc_hd__clkinv_2
XFILLER_17_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7730_ _7727_/Y _7726_/Y _9700_/Q _7729_/Y VGND VGND VPWR VPWR _7730_/Y sky130_fd_sc_hd__a31oi_1
X_7661_ _7661_/A _7661_/B _7661_/C _7661_/D VGND VGND VPWR VPWR _7662_/D sky130_fd_sc_hd__and4_2
XFILLER_177_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6612_ _9414_/Q VGND VGND VPWR VPWR _6612_/Y sky130_fd_sc_hd__clkinv_2
X_9400_ _9758_/CLK _9400_/D _9633_/SET_B VGND VGND VPWR VPWR _9400_/Q sky130_fd_sc_hd__dfrtp_1
X_4873_ _4865_/Y _5336_/B _4867_/Y _4868_/X _4872_/X VGND VGND VPWR VPWR _4896_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_60_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7592_ _6091_/Y _7400_/X _6139_/Y _7405_/X _7591_/X VGND VGND VPWR VPWR _7608_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_32_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6543_ _9461_/Q VGND VGND VPWR VPWR _6543_/Y sky130_fd_sc_hd__clkinv_4
X_9331_ _9771_/CLK _9331_/D _4628_/A VGND VGND VPWR VPWR _9331_/Q sky130_fd_sc_hd__dfstp_1
X_9262_ _9601_/CLK _9262_/D _9295_/SET_B VGND VGND VPWR VPWR _9262_/Q sky130_fd_sc_hd__dfrtp_1
X_6474_ _6474_/A _6474_/B _6474_/C _6474_/D VGND VGND VPWR VPWR _6475_/D sky130_fd_sc_hd__and4_1
XFILLER_9_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8213_ _8213_/A _8213_/B VGND VGND VPWR VPWR _8311_/B sky130_fd_sc_hd__or2_1
X_5425_ _9429_/Q _5422_/A _8844_/X _5422_/Y VGND VGND VPWR VPWR _9429_/D sky130_fd_sc_hd__a22o_1
XFILLER_145_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput210 _8754_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[11] sky130_fd_sc_hd__buf_2
XFILLER_118_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput232 _8794_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[31] sky130_fd_sc_hd__buf_2
Xoutput221 _8774_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[21] sky130_fd_sc_hd__buf_2
XFILLER_133_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9193_ _9378_/CLK _9193_/D _9646_/SET_B VGND VGND VPWR VPWR _9193_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput243 _7700_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[7] sky130_fd_sc_hd__buf_2
X_5356_ _5356_/A VGND VGND VPWR VPWR _5357_/A sky130_fd_sc_hd__clkbuf_4
X_8144_ _8144_/A _8362_/A _8575_/A _8627_/B VGND VGND VPWR VPWR _8144_/X sky130_fd_sc_hd__or4_1
Xoutput265 _9720_/Q VGND VGND VPWR VPWR pll_dco_ena sky130_fd_sc_hd__buf_2
Xoutput254 _7010_/Y VGND VGND VPWR VPWR pad_flash_csb_oeb sky130_fd_sc_hd__buf_2
Xoutput276 _9742_/Q VGND VGND VPWR VPWR pll_trim[10] sky130_fd_sc_hd__buf_2
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5287_ _9521_/Q _5280_/A _8840_/X _5280_/Y VGND VGND VPWR VPWR _9521_/D sky130_fd_sc_hd__a22o_1
X_8075_ _8585_/B _8075_/B VGND VGND VPWR VPWR _8075_/Y sky130_fd_sc_hd__nor2_1
Xoutput298 _9739_/Q VGND VGND VPWR VPWR pll_trim[7] sky130_fd_sc_hd__buf_2
Xoutput287 _9752_/Q VGND VGND VPWR VPWR pll_trim[20] sky130_fd_sc_hd__buf_2
X_7026_ _9250_/Q _9249_/Q VGND VGND VPWR VPWR _7027_/A sky130_fd_sc_hd__or2_1
XFILLER_101_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8977_ _8930_/S _6322_/Y _8977_/S VGND VGND VPWR VPWR _8977_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7928_ _8325_/A _7928_/B VGND VGND VPWR VPWR _7929_/B sky130_fd_sc_hd__and2_1
XFILLER_82_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7859_ _8521_/B _8262_/B VGND VGND VPWR VPWR _8463_/A sky130_fd_sc_hd__nor2_1
XFILLER_11_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9529_ _9534_/CLK _9529_/D _9647_/SET_B VGND VGND VPWR VPWR _9529_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_109_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5210_ _9571_/Q _5203_/Y _8930_/X _5203_/A VGND VGND VPWR VPWR _9571_/D sky130_fd_sc_hd__o22a_1
XFILLER_115_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6190_ _9422_/Q VGND VGND VPWR VPWR _6190_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_130_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5141_ _9621_/Q _5136_/A _8929_/A1 _5136_/Y VGND VGND VPWR VPWR _9621_/D sky130_fd_sc_hd__a22o_1
X_5072_ _8964_/X _9662_/Q _5078_/S VGND VGND VPWR VPWR _5073_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8900_ _7710_/X _9082_/Q _9051_/Q VGND VGND VPWR VPWR _8900_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8831_ _6544_/Y input2/X input1/X VGND VGND VPWR VPWR _8831_/X sky130_fd_sc_hd__mux2_2
X_8762_ _8762_/A VGND VGND VPWR VPWR _8762_/X sky130_fd_sc_hd__clkbuf_1
X_5974_ _9097_/Q _5970_/A _8925_/A1 _5970_/Y VGND VGND VPWR VPWR _9097_/D sky130_fd_sc_hd__a22o_1
X_7713_ _9084_/Q _7713_/B _9085_/Q VGND VGND VPWR VPWR _7716_/B sky130_fd_sc_hd__and3_1
X_8693_ _8693_/A _8693_/B _8693_/C _7929_/A VGND VGND VPWR VPWR _8696_/B sky130_fd_sc_hd__or4b_1
XFILLER_100_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4925_ _4925_/A _4931_/B VGND VGND VPWR VPWR _5366_/B sky130_fd_sc_hd__or2_4
XFILLER_193_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7644_ _7644_/A _7644_/B _7644_/C _7644_/D VGND VGND VPWR VPWR _7644_/Y sky130_fd_sc_hd__nand4_4
XFILLER_20_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4856_ _4911_/A _4917_/A VGND VGND VPWR VPWR _5317_/B sky130_fd_sc_hd__or2_4
XFILLER_165_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7575_ _6232_/Y _7419_/X _6189_/Y _7421_/X VGND VGND VPWR VPWR _7575_/X sky130_fd_sc_hd__o22a_1
XFILLER_20_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9314_ _9534_/CLK _9314_/D _9647_/SET_B VGND VGND VPWR VPWR _9314_/Q sky130_fd_sc_hd__dfrtp_1
X_6526_ _6526_/A _6526_/B _6526_/C _6526_/D VGND VGND VPWR VPWR _6629_/B sky130_fd_sc_hd__and4_1
X_4787_ _4787_/A _4921_/A VGND VGND VPWR VPWR _5488_/B sky130_fd_sc_hd__or2_4
XFILLER_173_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6457_ _9181_/Q VGND VGND VPWR VPWR _6457_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9245_ _9279_/CLK _9245_/D _9633_/SET_B VGND VGND VPWR VPWR _9245_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_133_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5408_ _9440_/Q _5406_/A _5964_/B1 _5406_/Y VGND VGND VPWR VPWR _9440_/D sky130_fd_sc_hd__a22o_1
X_6388_ _6386_/Y _6086_/X _6387_/Y _5336_/B VGND VGND VPWR VPWR _6388_/X sky130_fd_sc_hd__o22a_1
X_9176_ _9279_/CLK _9176_/D _9757_/SET_B VGND VGND VPWR VPWR _9176_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_125_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8127_ _8354_/A _8127_/B _8571_/A _8683_/B VGND VGND VPWR VPWR _8131_/A sky130_fd_sc_hd__or4_1
XFILLER_87_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5339_ _9488_/Q _5338_/A _5963_/B1 _5338_/Y VGND VGND VPWR VPWR _9488_/D sky130_fd_sc_hd__a22o_1
XFILLER_125_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8058_ _8521_/B VGND VGND VPWR VPWR _8061_/A sky130_fd_sc_hd__inv_2
XFILLER_125_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7009_ _9051_/Q _5993_/B _9050_/Q _7008_/X VGND VGND VPWR VPWR _9050_/D sky130_fd_sc_hd__a22o_1
XFILLER_47_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4710_ _9281_/Q VGND VGND VPWR VPWR _7304_/A sky130_fd_sc_hd__inv_2
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5690_ _9053_/Q VGND VGND VPWR VPWR _5691_/A sky130_fd_sc_hd__inv_2
XFILLER_30_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4641_ _4994_/A VGND VGND VPWR VPWR _4642_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_175_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7360_ _6589_/Y _7095_/X _6477_/Y _7068_/D _7359_/X VGND VGND VPWR VPWR _7365_/B
+ sky130_fd_sc_hd__o221a_1
X_4572_ _9750_/Q _4566_/A _5965_/B1 _4566_/Y VGND VGND VPWR VPWR _9750_/D sky130_fd_sc_hd__a22o_1
XFILLER_155_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6311_ _9317_/Q VGND VGND VPWR VPWR _6311_/Y sky130_fd_sc_hd__inv_2
X_7291_ _4677_/Y _7040_/C _4775_/Y _7059_/C VGND VGND VPWR VPWR _7291_/X sky130_fd_sc_hd__o22a_1
X_9030_ _9039_/CLK _9030_/D VGND VGND VPWR VPWR _9030_/Q sky130_fd_sc_hd__dfxtp_1
X_6242_ _6240_/Y _5306_/B _6241_/Y _4491_/B VGND VGND VPWR VPWR _6242_/X sky130_fd_sc_hd__o22a_1
XFILLER_143_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6173_ _6168_/Y _5278_/B _6169_/Y _5306_/B _6172_/X VGND VGND VPWR VPWR _6174_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_130_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5124_ _9631_/Q _5123_/A _5963_/B1 _5123_/Y VGND VGND VPWR VPWR _9631_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5055_ _9667_/Q _5047_/A _8916_/A1 _5047_/Y VGND VGND VPWR VPWR _9667_/D sky130_fd_sc_hd__a22o_1
XFILLER_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8814_ _9791_/Q _6251_/Y _8916_/A1 _6251_/A _8939_/X VGND VGND VPWR VPWR _9791_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_80_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5957_ _9108_/Q _5951_/A _8955_/A1 _5951_/Y VGND VGND VPWR VPWR _9108_/D sky130_fd_sc_hd__a22o_1
XFILLER_71_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8745_ _8745_/A VGND VGND VPWR VPWR _8746_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_52_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8676_ _8676_/A _8676_/B VGND VGND VPWR VPWR _8677_/B sky130_fd_sc_hd__or2_1
X_4908_ _9740_/Q VGND VGND VPWR VPWR _4908_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7627_ _6866_/Y _7408_/X _6902_/Y _7410_/X VGND VGND VPWR VPWR _7627_/X sky130_fd_sc_hd__o22a_1
X_5888_ _5849_/X _8887_/X _8924_/X _9145_/Q VGND VGND VPWR VPWR _9145_/D sky130_fd_sc_hd__o22a_1
XFILLER_21_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4839_ _4831_/Y _4832_/X _4833_/Y _5431_/B _4838_/X VGND VGND VPWR VPWR _4864_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_181_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7558_ _6301_/Y _7415_/X _6297_/Y _7417_/X _7557_/X VGND VGND VPWR VPWR _7572_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_134_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6509_ _9323_/Q VGND VGND VPWR VPWR _8763_/A sky130_fd_sc_hd__clkinv_8
X_7489_ _6799_/Y _7430_/X _6860_/Y _7432_/X _7488_/X VGND VGND VPWR VPWR _7489_/X
+ sky130_fd_sc_hd__o221a_1
X_9228_ _9440_/CLK _9228_/D _9685_/SET_B VGND VGND VPWR VPWR _9228_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_20_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9159_ _9358_/CLK _9159_/D _9528_/SET_B VGND VGND VPWR VPWR _9159_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_121_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_6 _7265_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6860_ _9547_/Q VGND VGND VPWR VPWR _6860_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5811_ _5811_/A VGND VGND VPWR VPWR _5812_/A sky130_fd_sc_hd__clkbuf_2
X_6791_ _6789_/Y _4602_/B _6790_/Y _4524_/B VGND VGND VPWR VPWR _6791_/X sky130_fd_sc_hd__o22a_4
XFILLER_34_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5742_ _5960_/A _5742_/B VGND VGND VPWR VPWR _5743_/A sky130_fd_sc_hd__or2_1
X_8530_ _8472_/Y _8528_/Y _8518_/X _8459_/C VGND VGND VPWR VPWR _8614_/D sky130_fd_sc_hd__a31o_1
XFILLER_22_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5673_ _5673_/A VGND VGND VPWR VPWR _5673_/Y sky130_fd_sc_hd__inv_2
X_8461_ _8461_/A _8627_/A VGND VGND VPWR VPWR _8464_/B sky130_fd_sc_hd__or2_1
XFILLER_163_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8392_ _8392_/A VGND VGND VPWR VPWR _8708_/A sky130_fd_sc_hd__inv_2
X_7412_ _4877_/Y _7400_/X _4720_/Y _7405_/X _7411_/X VGND VGND VPWR VPWR _7481_/A
+ sky130_fd_sc_hd__o221a_1
X_4624_ _5966_/B1 _9720_/Q _4626_/S VGND VGND VPWR VPWR _4625_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7343_ _7343_/A _7343_/B _7343_/C _7343_/D VGND VGND VPWR VPWR _7353_/B sky130_fd_sc_hd__and4_1
X_4555_ _5967_/B1 _9758_/Q _4555_/S VGND VGND VPWR VPWR _4556_/A sky130_fd_sc_hd__mux2_1
X_4486_ _4486_/A VGND VGND VPWR VPWR _9786_/D sky130_fd_sc_hd__clkbuf_1
X_9013_ _9039_/CLK _9013_/D VGND VGND VPWR VPWR _9013_/Q sky130_fd_sc_hd__dfxtp_1
X_7274_ _6067_/Y _7059_/B _6081_/A _7068_/C _7273_/X VGND VGND VPWR VPWR _7277_/C
+ sky130_fd_sc_hd__o221a_1
X_6225_ _9430_/Q VGND VGND VPWR VPWR _6225_/Y sky130_fd_sc_hd__inv_2
X_6156_ _6151_/Y _5545_/B _6152_/Y _5496_/B _6155_/X VGND VGND VPWR VPWR _6174_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_97_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5107_ _9641_/Q _5102_/A _5967_/B1 _5102_/Y VGND VGND VPWR VPWR _9641_/D sky130_fd_sc_hd__a22o_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater362 _8842_/X VGND VGND VPWR VPWR _5964_/B1 sky130_fd_sc_hd__buf_12
X_6087_ _6087_/A VGND VGND VPWR VPWR _6087_/Y sky130_fd_sc_hd__inv_2
Xrepeater373 _9647_/SET_B VGND VGND VPWR VPWR _9528_/SET_B sky130_fd_sc_hd__buf_12
XFILLER_38_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5038_ _8975_/X _4551_/B _9681_/Q _5062_/D VGND VGND VPWR VPWR _9681_/D sky130_fd_sc_hd__a22o_1
XFILLER_167_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9777_ _9777_/CLK _9777_/D _7011_/B VGND VGND VPWR VPWR _9777_/Q sky130_fd_sc_hd__dfrtp_1
X_6989_ _8813_/A _8809_/A _6950_/B VGND VGND VPWR VPWR _9068_/D sky130_fd_sc_hd__o21ai_1
X_8728_ _8728_/A VGND VGND VPWR VPWR _8728_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8659_ _8659_/A _8659_/B _8659_/C _7893_/X VGND VGND VPWR VPWR _8727_/C sky130_fd_sc_hd__or4b_1
XFILLER_166_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput110 sram_ro_data[25] VGND VGND VPWR VPWR _6817_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput132 wb_adr_i[0] VGND VGND VPWR VPWR _7839_/A sky130_fd_sc_hd__clkbuf_4
Xinput154 wb_adr_i[2] VGND VGND VPWR VPWR _8379_/B sky130_fd_sc_hd__buf_4
Xinput143 wb_adr_i[1] VGND VGND VPWR VPWR _8394_/C sky130_fd_sc_hd__buf_4
XFILLER_76_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput121 sram_ro_data[6] VGND VGND VPWR VPWR _6233_/A sky130_fd_sc_hd__clkbuf_1
Xinput187 wb_dat_i[2] VGND VGND VPWR VPWR _8963_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput176 wb_dat_i[1] VGND VGND VPWR VPWR _8962_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput165 wb_dat_i[0] VGND VGND VPWR VPWR _8961_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_102_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput198 wb_sel_i[0] VGND VGND VPWR VPWR _5059_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_63_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6010_ _6010_/A VGND VGND VPWR VPWR _6010_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_79_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7961_ _7959_/A _8195_/B _7960_/Y VGND VGND VPWR VPWR _7979_/A sky130_fd_sc_hd__a21oi_1
XFILLER_94_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6912_ _6908_/Y _5089_/B _6909_/Y _5864_/B _6911_/X VGND VGND VPWR VPWR _6925_/B
+ sky130_fd_sc_hd__o221a_1
X_7892_ _8515_/B _8305_/A _8496_/A _8305_/B VGND VGND VPWR VPWR _7892_/X sky130_fd_sc_hd__a211o_1
X_9700_ _9709_/CLK _9700_/D _4987_/X VGND VGND VPWR VPWR _9700_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6843_ _9490_/Q VGND VGND VPWR VPWR _6843_/Y sky130_fd_sc_hd__clkinv_2
X_9631_ _9757_/CLK _9631_/D _9757_/SET_B VGND VGND VPWR VPWR _9631_/Q sky130_fd_sc_hd__dfstp_1
X_9562_ _9617_/CLK _9562_/D _9295_/SET_B VGND VGND VPWR VPWR _9562_/Q sky130_fd_sc_hd__dfrtp_1
X_6774_ _9629_/Q VGND VGND VPWR VPWR _6774_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8513_ _8513_/A VGND VGND VPWR VPWR _8513_/X sky130_fd_sc_hd__clkbuf_1
X_9493_ _9493_/CLK _9493_/D _4628_/A VGND VGND VPWR VPWR _9493_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5725_ _9250_/Q _5725_/B VGND VGND VPWR VPWR _5726_/A sky130_fd_sc_hd__or2_1
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8444_ _8444_/A _8444_/B VGND VGND VPWR VPWR _8448_/B sky130_fd_sc_hd__or2_1
X_5656_ _5647_/A _5658_/A _5751_/C VGND VGND VPWR VPWR _5656_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_163_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4607_ _9729_/Q _4604_/A _5964_/B1 _4604_/Y VGND VGND VPWR VPWR _9729_/D sky130_fd_sc_hd__a22o_1
X_8375_ _8375_/A _8582_/A _8678_/A _8646_/A VGND VGND VPWR VPWR _8380_/A sky130_fd_sc_hd__or4_1
X_5587_ _9318_/Q _5585_/A _8845_/X _5585_/Y VGND VGND VPWR VPWR _9318_/D sky130_fd_sc_hd__a22o_1
XFILLER_116_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7326_ _7326_/A _7392_/B VGND VGND VPWR VPWR _7326_/X sky130_fd_sc_hd__or2_1
XFILLER_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4538_ _5967_/B1 _9761_/Q _4540_/S VGND VGND VPWR VPWR _4539_/A sky130_fd_sc_hd__mux2_1
X_7257_ _6194_/Y _7040_/D _6154_/Y _7110_/X _7256_/X VGND VGND VPWR VPWR _7264_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_117_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4469_ _4456_/Y _8942_/X _8941_/X VGND VGND VPWR VPWR _4801_/C sky130_fd_sc_hd__a21bo_1
XFILLER_104_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6208_ _6208_/A VGND VGND VPWR VPWR _6208_/Y sky130_fd_sc_hd__inv_2
X_7188_ _8751_/A _7048_/D _6517_/Y _7040_/B _7187_/X VGND VGND VPWR VPWR _7189_/D
+ sky130_fd_sc_hd__o221a_1
X_6139_ _9263_/Q VGND VGND VPWR VPWR _6139_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_5_csclk clkbuf_2_2_0_csclk/X VGND VGND VPWR VPWR _9789_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_174_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5510_ _9371_/Q _5509_/A _8846_/X _5509_/Y VGND VGND VPWR VPWR _9371_/D sky130_fd_sc_hd__a22o_1
XFILLER_145_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6490_ _9096_/Q VGND VGND VPWR VPWR _7705_/A sky130_fd_sc_hd__inv_6
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5441_ _9416_/Q _5433_/A _8916_/A1 _5433_/Y VGND VGND VPWR VPWR _9416_/D sky130_fd_sc_hd__a22o_1
XFILLER_172_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8160_ _8160_/A _8645_/A VGND VGND VPWR VPWR _8162_/A sky130_fd_sc_hd__or2_1
X_5372_ _9464_/Q _5368_/A _5966_/B1 _5368_/Y VGND VGND VPWR VPWR _9464_/D sky130_fd_sc_hd__a22o_1
X_8091_ _8525_/A _8091_/B _8386_/A VGND VGND VPWR VPWR _8093_/B sky130_fd_sc_hd__or3_1
XFILLER_99_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7111_ _9246_/Q _9245_/Q _7111_/C _7127_/C VGND VGND VPWR VPWR _7112_/A sky130_fd_sc_hd__or4_2
XFILLER_141_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7042_ _7127_/A _7127_/B _7073_/C VGND VGND VPWR VPWR _7043_/A sky130_fd_sc_hd__or3_1
XFILLER_86_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8993_ _9561_/Q _8763_/A VGND VGND VPWR VPWR mgmt_gpio_out[16] sky130_fd_sc_hd__ebufn_8
XFILLER_67_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7944_ _7944_/A VGND VGND VPWR VPWR _7944_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_82_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7875_ _8525_/A _7894_/B _7903_/C _8193_/A VGND VGND VPWR VPWR _8230_/A sky130_fd_sc_hd__or4_4
X_9614_ _9788_/CLK _9614_/D _9295_/SET_B VGND VGND VPWR VPWR _9614_/Q sky130_fd_sc_hd__dfrtp_1
X_6826_ _9433_/Q VGND VGND VPWR VPWR _6826_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6757_ _6755_/Y _5872_/B _6756_/Y _5526_/B VGND VGND VPWR VPWR _6757_/X sky130_fd_sc_hd__o22a_1
XFILLER_11_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9545_ _9545_/CLK _9545_/D _4628_/A VGND VGND VPWR VPWR _9545_/Q sky130_fd_sc_hd__dfrtp_1
X_5708_ _9251_/Q VGND VGND VPWR VPWR _7401_/B sky130_fd_sc_hd__inv_2
X_9476_ _9527_/CLK _9476_/D _9685_/SET_B VGND VGND VPWR VPWR _9476_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_163_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6688_ input45/X _8926_/S _6687_/Y _5837_/B VGND VGND VPWR VPWR _6688_/X sky130_fd_sc_hd__o2bb2a_1
X_5639_ _9281_/Q _5634_/A _8839_/X _5634_/Y VGND VGND VPWR VPWR _9281_/D sky130_fd_sc_hd__a22o_1
X_8427_ _8427_/A _8601_/D VGND VGND VPWR VPWR _8428_/B sky130_fd_sc_hd__or2_1
XFILLER_12_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8358_ _8358_/A _8358_/B VGND VGND VPWR VPWR _8642_/C sky130_fd_sc_hd__or2_1
XFILLER_151_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7309_ _7309_/A _7309_/B _7309_/C VGND VGND VPWR VPWR _7309_/Y sky130_fd_sc_hd__nand3_4
XFILLER_2_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8289_ _8625_/A _8340_/B _8340_/C _8288_/X VGND VGND VPWR VPWR _8290_/B sky130_fd_sc_hd__a31o_1
XFILLER_144_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5990_ _6040_/A VGND VGND VPWR VPWR _5991_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_91_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4941_ _9091_/Q VGND VGND VPWR VPWR _6022_/D sky130_fd_sc_hd__inv_2
X_7660_ _6750_/Y _7471_/X _7348_/A _7473_/X _7659_/X VGND VGND VPWR VPWR _7661_/D
+ sky130_fd_sc_hd__o221a_1
X_4872_ _4869_/Y _4870_/X _4871_/Y _4558_/B VGND VGND VPWR VPWR _4872_/X sky130_fd_sc_hd__o22a_2
XFILLER_17_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6611_ _9427_/Q VGND VGND VPWR VPWR _8771_/A sky130_fd_sc_hd__inv_6
XFILLER_192_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7591_ _6078_/Y _7408_/X _6059_/Y _7410_/X VGND VGND VPWR VPWR _7591_/X sky130_fd_sc_hd__o22a_1
XFILLER_20_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9330_ _9776_/CLK _9330_/D _4628_/A VGND VGND VPWR VPWR _9330_/Q sky130_fd_sc_hd__dfrtp_1
X_6542_ _8799_/A _5507_/B _6530_/X _6536_/X _6541_/X VGND VGND VPWR VPWR _6629_/C
+ sky130_fd_sc_hd__o2111a_1
X_9261_ _9601_/CLK _9261_/D _9295_/SET_B VGND VGND VPWR VPWR _9261_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_145_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6473_ _6473_/A _6473_/B _6473_/C _6473_/D VGND VGND VPWR VPWR _6474_/D sky130_fd_sc_hd__and4_1
X_5424_ _9430_/Q _5422_/A _8845_/X _5422_/Y VGND VGND VPWR VPWR _9430_/D sky130_fd_sc_hd__a22o_1
X_8212_ _8341_/B _8260_/B _8312_/D VGND VGND VPWR VPWR _8224_/B sky130_fd_sc_hd__o21ai_1
X_9192_ _9378_/CLK _9192_/D _9646_/SET_B VGND VGND VPWR VPWR _9192_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput233 _8796_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[32] sky130_fd_sc_hd__buf_2
Xoutput222 _8776_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[22] sky130_fd_sc_hd__buf_2
XFILLER_133_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput211 _8756_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[12] sky130_fd_sc_hd__buf_2
Xoutput244 _8748_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[8] sky130_fd_sc_hd__buf_2
X_8143_ _8164_/A _8551_/A VGND VGND VPWR VPWR _8627_/B sky130_fd_sc_hd__nor2_1
X_5355_ _5545_/A _5355_/B VGND VGND VPWR VPWR _5356_/A sky130_fd_sc_hd__or2_1
Xoutput266 _9721_/Q VGND VGND VPWR VPWR pll_div[0] sky130_fd_sc_hd__buf_2
Xoutput255 _8838_/X VGND VGND VPWR VPWR pad_flash_io0_do sky130_fd_sc_hd__buf_2
Xoutput277 _9743_/Q VGND VGND VPWR VPWR pll_trim[11] sky130_fd_sc_hd__buf_2
X_5286_ _9522_/Q _5280_/A _8955_/A1 _5280_/Y VGND VGND VPWR VPWR _9522_/D sky130_fd_sc_hd__a22o_1
X_8074_ _8074_/A _8704_/A VGND VGND VPWR VPWR _8075_/B sky130_fd_sc_hd__or2_1
XFILLER_114_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput299 _9740_/Q VGND VGND VPWR VPWR pll_trim[8] sky130_fd_sc_hd__buf_2
Xoutput288 _9753_/Q VGND VGND VPWR VPWR pll_trim[21] sky130_fd_sc_hd__buf_2
XFILLER_141_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7025_ _7025_/A VGND VGND VPWR VPWR _7079_/B sky130_fd_sc_hd__buf_8
XFILLER_101_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8976_ _8926_/S _6322_/Y _8977_/S VGND VGND VPWR VPWR _8976_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7927_ _8615_/A _7927_/B VGND VGND VPWR VPWR _7928_/B sky130_fd_sc_hd__nor2_1
X_7858_ _7858_/A VGND VGND VPWR VPWR _8262_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6809_ _6807_/Y _4481_/B _6808_/Y _4893_/X VGND VGND VPWR VPWR _6809_/X sky130_fd_sc_hd__o22a_1
XFILLER_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7789_ _7903_/C _7823_/A _8528_/A _8193_/A _7787_/X VGND VGND VPWR VPWR _7900_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_156_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9528_ _9535_/CLK _9528_/D _9528_/SET_B VGND VGND VPWR VPWR _9528_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_139_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9459_ _9532_/CLK _9459_/D _9647_/SET_B VGND VGND VPWR VPWR _9459_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_151_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_23_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR _9617_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_38_csclk clkbuf_2_1_0_csclk/X VGND VGND VPWR VPWR _9757_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_6_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5140_ _9622_/Q _5136_/A _8925_/A1 _5136_/Y VGND VGND VPWR VPWR _9622_/D sky130_fd_sc_hd__a22o_1
X_5071_ _5071_/A VGND VGND VPWR VPWR _9663_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8830_ _9593_/Q input91/X _8835_/S VGND VGND VPWR VPWR _8830_/X sky130_fd_sc_hd__mux2_1
XFILLER_92_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8761_ _8761_/A VGND VGND VPWR VPWR _8762_/A sky130_fd_sc_hd__clkbuf_1
X_5973_ _9098_/Q _5970_/A _8844_/X _5970_/Y VGND VGND VPWR VPWR _9098_/D sky130_fd_sc_hd__a22o_1
XFILLER_25_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4924_ _9463_/Q VGND VGND VPWR VPWR _4924_/Y sky130_fd_sc_hd__clkinv_2
X_7712_ _9084_/Q _7713_/B _9084_/Q _7713_/B VGND VGND VPWR VPWR _7712_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_178_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8692_ _8671_/Y _8673_/X _8680_/Y _8682_/X _8691_/Y VGND VGND VPWR VPWR _8692_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_33_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4855_ _9494_/Q VGND VGND VPWR VPWR _4855_/Y sky130_fd_sc_hd__inv_2
X_7643_ _7643_/A _7643_/B _7643_/C _7643_/D VGND VGND VPWR VPWR _7644_/D sky130_fd_sc_hd__and4_1
XFILLER_20_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7574_ _6152_/Y _7400_/X _6178_/Y _7405_/X _7573_/X VGND VGND VPWR VPWR _7590_/A
+ sky130_fd_sc_hd__o221a_1
X_4786_ _9380_/Q VGND VGND VPWR VPWR _4786_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9313_ _9534_/CLK _9313_/D _9647_/SET_B VGND VGND VPWR VPWR _9313_/Q sky130_fd_sc_hd__dfstp_1
X_6525_ _8747_/A _5837_/B _6521_/Y _6135_/A _6524_/X VGND VGND VPWR VPWR _6526_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_134_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9244_ _9789_/CLK _9244_/D _9685_/SET_B VGND VGND VPWR VPWR _9244_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_109_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6456_ _9110_/Q VGND VGND VPWR VPWR _6456_/Y sky130_fd_sc_hd__clkinv_2
X_5407_ _9441_/Q _5406_/A _5963_/B1 _5406_/Y VGND VGND VPWR VPWR _9441_/D sky130_fd_sc_hd__a22o_1
X_6387_ _9488_/Q VGND VGND VPWR VPWR _6387_/Y sky130_fd_sc_hd__clkinv_4
X_9175_ _9280_/CLK _9175_/D _9757_/SET_B VGND VGND VPWR VPWR _9175_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_125_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8126_ _8164_/A _8130_/B VGND VGND VPWR VPWR _8683_/B sky130_fd_sc_hd__nor2_1
XFILLER_87_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5338_ _5338_/A VGND VGND VPWR VPWR _5338_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8057_ _8057_/A _8536_/A VGND VGND VPWR VPWR _8062_/A sky130_fd_sc_hd__nand2_1
XFILLER_102_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5269_ _5269_/A VGND VGND VPWR VPWR _5269_/Y sky130_fd_sc_hd__clkinv_2
X_7008_ _7008_/A _7008_/B VGND VGND VPWR VPWR _7008_/X sky130_fd_sc_hd__or2_1
XFILLER_47_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8959_ _7133_/X _4875_/Y _8959_/S VGND VGND VPWR VPWR _8959_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4640_ _9717_/Q _4636_/A _8948_/X _4636_/Y VGND VGND VPWR VPWR hold2/A sky130_fd_sc_hd__a22o_1
XFILLER_175_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6310_ _9395_/Q VGND VGND VPWR VPWR _6310_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_128_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4571_ _9751_/Q _4566_/A _5964_/B1 _4566_/Y VGND VGND VPWR VPWR _9751_/D sky130_fd_sc_hd__a22o_1
XFILLER_183_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7290_ _4888_/Y _7082_/X _4865_/Y _7084_/X _7289_/X VGND VGND VPWR VPWR _7309_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_89_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6241_ _9783_/Q VGND VGND VPWR VPWR _6241_/Y sky130_fd_sc_hd__inv_2
X_6172_ _6170_/Y _5621_/B _6171_/Y _5267_/B VGND VGND VPWR VPWR _6172_/X sky130_fd_sc_hd__o22a_1
XFILLER_131_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5123_ _5123_/A VGND VGND VPWR VPWR _5123_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5054_ _9668_/Q _5047_/A _8930_/A1 _5047_/Y VGND VGND VPWR VPWR _9668_/D sky130_fd_sc_hd__a22o_1
X_8813_ _8813_/A _8813_/B VGND VGND VPWR VPWR _9060_/D sky130_fd_sc_hd__nor2_1
XFILLER_65_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5956_ _9109_/Q _5951_/A _8929_/A1 _5951_/Y VGND VGND VPWR VPWR _9109_/D sky130_fd_sc_hd__a22o_1
XFILLER_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8744_ _8744_/A VGND VGND VPWR VPWR _8744_/X sky130_fd_sc_hd__clkbuf_1
X_8675_ _8675_/A _8675_/B _8675_/C _8675_/D VGND VGND VPWR VPWR _8716_/D sky130_fd_sc_hd__or4_4
X_5887_ _5849_/X _8889_/X _8924_/X _9146_/Q VGND VGND VPWR VPWR _9146_/D sky130_fd_sc_hd__o22a_1
XFILLER_33_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4907_ _6158_/A _6111_/B VGND VGND VPWR VPWR _4907_/X sky130_fd_sc_hd__or2_4
XFILLER_178_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7626_ _7626_/A _7626_/B _7626_/C _7626_/D VGND VGND VPWR VPWR _7626_/Y sky130_fd_sc_hd__nand4_4
X_4838_ _4835_/Y _4481_/B _4836_/Y _5232_/B VGND VGND VPWR VPWR _4838_/X sky130_fd_sc_hd__o22a_1
XFILLER_166_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4769_ _9646_/Q VGND VGND VPWR VPWR _4769_/Y sky130_fd_sc_hd__inv_2
X_7557_ _6282_/Y _7419_/X _6241_/Y _7421_/X VGND VGND VPWR VPWR _7557_/X sky130_fd_sc_hd__o22a_1
X_6508_ _9336_/Q VGND VGND VPWR VPWR _6508_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7488_ _6788_/Y _7434_/X _6854_/Y _7436_/X VGND VGND VPWR VPWR _7488_/X sky130_fd_sc_hd__o22a_1
XFILLER_134_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6439_ _9650_/Q VGND VGND VPWR VPWR _6439_/Y sky130_fd_sc_hd__clkinv_4
X_9227_ _9440_/CLK _9227_/D _9685_/SET_B VGND VGND VPWR VPWR _9227_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_161_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9158_ _9695_/CLK _9158_/D _9646_/SET_B VGND VGND VPWR VPWR _9158_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8109_ _8640_/A VGND VGND VPWR VPWR _8110_/C sky130_fd_sc_hd__inv_2
XFILLER_102_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9089_ _9089_/CLK _9089_/D _5991_/X VGND VGND VPWR VPWR _9089_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_7 _7265_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5810_ _5960_/A _5810_/B VGND VGND VPWR VPWR _5811_/A sky130_fd_sc_hd__or2_1
XFILLER_62_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6790_ _9763_/Q VGND VGND VPWR VPWR _6790_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5741_ _9245_/Q _5713_/A _5738_/B _5724_/B VGND VGND VPWR VPWR _9245_/D sky130_fd_sc_hd__o22a_1
X_8460_ _8460_/A VGND VGND VPWR VPWR _8627_/A sky130_fd_sc_hd__inv_2
X_5672_ _5672_/A VGND VGND VPWR VPWR _5673_/A sky130_fd_sc_hd__clkbuf_2
X_7411_ _4897_/Y _7408_/X _4842_/Y _7410_/X VGND VGND VPWR VPWR _7411_/X sky130_fd_sc_hd__o22a_1
XFILLER_30_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8391_ _8544_/C VGND VGND VPWR VPWR _8401_/B sky130_fd_sc_hd__clkinv_4
X_4623_ _5259_/A _4623_/B VGND VGND VPWR VPWR _4626_/S sky130_fd_sc_hd__or2_1
XFILLER_30_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7342_ _6646_/Y _7048_/D _6745_/Y _7040_/B _7341_/X VGND VGND VPWR VPWR _7343_/D
+ sky130_fd_sc_hd__o221a_1
X_4554_ _6158_/A _4925_/A _5259_/A VGND VGND VPWR VPWR _4555_/S sky130_fd_sc_hd__or3_1
XFILLER_143_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7273_ _6103_/Y _7079_/B _6066_/Y _7059_/A VGND VGND VPWR VPWR _7273_/X sky130_fd_sc_hd__o22a_1
XFILLER_116_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4485_ _8840_/X _9786_/Q _6018_/S VGND VGND VPWR VPWR _4486_/A sky130_fd_sc_hd__mux2_1
X_9012_ _9027_/CLK _9012_/D VGND VGND VPWR VPWR _9012_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6224_ _9131_/Q VGND VGND VPWR VPWR _6224_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_131_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6155_ _6153_/Y _4870_/X _6154_/Y _5534_/B VGND VGND VPWR VPWR _6155_/X sky130_fd_sc_hd__o22a_1
XFILLER_85_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5106_ _9642_/Q _5102_/A _5966_/B1 _5102_/Y VGND VGND VPWR VPWR _9642_/D sky130_fd_sc_hd__a22o_1
X_6086_ _6158_/A _6086_/B VGND VGND VPWR VPWR _6086_/X sky130_fd_sc_hd__or2_4
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5037_ _9049_/Q _5034_/Y _5985_/B _9682_/Q VGND VGND VPWR VPWR _9682_/D sky130_fd_sc_hd__a31o_1
Xrepeater363 _8842_/X VGND VGND VPWR VPWR _8929_/A1 sky130_fd_sc_hd__buf_12
Xrepeater374 _9685_/SET_B VGND VGND VPWR VPWR _9647_/SET_B sky130_fd_sc_hd__buf_12
XFILLER_122_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9776_ _9776_/CLK _9776_/D _7011_/B VGND VGND VPWR VPWR _9776_/Q sky130_fd_sc_hd__dfrtp_1
X_6988_ _8812_/A _8809_/A _6962_/B VGND VGND VPWR VPWR _9067_/D sky130_fd_sc_hd__o21ai_1
X_8727_ _8727_/A _8727_/B _8727_/C _8727_/D VGND VGND VPWR VPWR _8728_/A sky130_fd_sc_hd__or4_1
XFILLER_40_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5939_ _5939_/A _5939_/B VGND VGND VPWR VPWR _5939_/X sky130_fd_sc_hd__or2_1
X_8658_ _8676_/B _8658_/B VGND VGND VPWR VPWR _8659_/B sky130_fd_sc_hd__or2_1
XFILLER_21_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8589_ _8650_/B _8650_/C _8651_/B _8588_/X VGND VGND VPWR VPWR _8589_/X sky130_fd_sc_hd__or4b_2
XFILLER_154_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7609_ _4924_/Y _7408_/X _4692_/A _7410_/X VGND VGND VPWR VPWR _7609_/X sky130_fd_sc_hd__o22a_1
XFILLER_147_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput111 sram_ro_data[26] VGND VGND VPWR VPWR _6669_/A sky130_fd_sc_hd__clkbuf_1
Xinput100 sram_ro_data[16] VGND VGND VPWR VPWR _4840_/A sky130_fd_sc_hd__clkbuf_1
Xinput144 wb_adr_i[20] VGND VGND VPWR VPWR _7837_/B sky130_fd_sc_hd__buf_2
Xinput133 wb_adr_i[10] VGND VGND VPWR VPWR _7771_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_88_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput122 sram_ro_data[7] VGND VGND VPWR VPWR _6075_/A sky130_fd_sc_hd__clkbuf_1
Xinput177 wb_dat_i[20] VGND VGND VPWR VPWR _7744_/B sky130_fd_sc_hd__clkbuf_1
Xinput166 wb_dat_i[10] VGND VGND VPWR VPWR _7741_/B2 sky130_fd_sc_hd__clkbuf_1
Xinput155 wb_adr_i[30] VGND VGND VPWR VPWR _5931_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_76_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput199 wb_sel_i[1] VGND VGND VPWR VPWR _5058_/B sky130_fd_sc_hd__clkbuf_1
Xinput188 wb_dat_i[30] VGND VGND VPWR VPWR _7749_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7960_ _8193_/B VGND VGND VPWR VPWR _7960_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7891_ _7896_/A _8305_/B VGND VGND VPWR VPWR _8441_/A sky130_fd_sc_hd__or2_1
X_6911_ input62/X _4680_/Y _6910_/Y _5045_/B VGND VGND VPWR VPWR _6911_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_94_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9630_ _9639_/CLK _9630_/D _9757_/SET_B VGND VGND VPWR VPWR _9630_/Q sky130_fd_sc_hd__dfstp_1
X_6842_ _6837_/Y _5121_/B _6838_/Y _5110_/B _6841_/X VGND VGND VPWR VPWR _6878_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_62_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9561_ _9788_/CLK _9561_/D _9295_/SET_B VGND VGND VPWR VPWR _9561_/Q sky130_fd_sc_hd__dfrtp_1
X_6773_ _9648_/Q VGND VGND VPWR VPWR _6773_/Y sky130_fd_sc_hd__inv_2
X_8512_ _8603_/A _8512_/B _8603_/C _8512_/D VGND VGND VPWR VPWR _8513_/A sky130_fd_sc_hd__or4_1
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5724_ _5725_/B _5724_/B _7041_/A VGND VGND VPWR VPWR _5724_/Y sky130_fd_sc_hd__nor3_1
X_9492_ _9545_/CLK _9492_/D _4628_/A VGND VGND VPWR VPWR _9492_/Q sky130_fd_sc_hd__dfrtp_1
X_8443_ _7902_/B _8624_/B _7896_/X VGND VGND VPWR VPWR _8444_/B sky130_fd_sc_hd__o21ai_1
X_5655_ _5649_/B _5647_/X _5658_/A _5654_/X VGND VGND VPWR VPWR _9279_/D sky130_fd_sc_hd__o2bb2a_1
X_8374_ _8204_/A _8279_/C _8280_/C VGND VGND VPWR VPWR _8646_/A sky130_fd_sc_hd__o21ai_1
X_4606_ _9730_/Q _4604_/A _5963_/B1 _4604_/Y VGND VGND VPWR VPWR _9730_/D sky130_fd_sc_hd__a22o_1
X_5586_ _9319_/Q _5585_/A _8846_/X _5585_/Y VGND VGND VPWR VPWR _9319_/D sky130_fd_sc_hd__a22o_1
X_7325_ _6929_/Y _7059_/D _6801_/Y _7116_/X _7324_/X VGND VGND VPWR VPWR _7330_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_7_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4537_ _5259_/A _4537_/B VGND VGND VPWR VPWR _4540_/S sky130_fd_sc_hd__or2_2
XFILLER_171_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7256_ _6176_/Y _7112_/X _6212_/Y _7077_/B VGND VGND VPWR VPWR _7256_/X sky130_fd_sc_hd__o22a_1
XFILLER_116_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4468_ _8938_/X VGND VGND VPWR VPWR _4665_/B sky130_fd_sc_hd__inv_2
X_7187_ _8753_/A _7068_/A _8785_/A _7105_/X VGND VGND VPWR VPWR _7187_/X sky130_fd_sc_hd__o22a_1
X_6207_ _6207_/A VGND VGND VPWR VPWR _6207_/Y sky130_fd_sc_hd__inv_2
X_6138_ _9301_/Q VGND VGND VPWR VPWR _7282_/A sky130_fd_sc_hd__clkinv_2
XFILLER_131_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6069_ _6067_/Y _5621_/B _6068_/Y _5507_/B VGND VGND VPWR VPWR _6069_/X sky130_fd_sc_hd__o22a_1
XFILLER_85_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9759_ _4450_/A1 _9759_/D _6146_/A VGND VGND VPWR VPWR _9759_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5440_ _9417_/Q _5433_/A _8840_/X _5433_/Y VGND VGND VPWR VPWR _9417_/D sky130_fd_sc_hd__a22o_1
XFILLER_157_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5371_ _9465_/Q _5368_/A _5965_/B1 _5368_/Y VGND VGND VPWR VPWR _9465_/D sky130_fd_sc_hd__a22o_1
X_8090_ _8218_/A _8096_/B _7968_/A _8120_/A VGND VGND VPWR VPWR _8386_/A sky130_fd_sc_hd__or4bb_4
XFILLER_153_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7110_ _7110_/A VGND VGND VPWR VPWR _7110_/X sky130_fd_sc_hd__buf_8
X_7041_ _7041_/A _7073_/C VGND VGND VPWR VPWR _7392_/B sky130_fd_sc_hd__or2_4
XFILLER_113_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8992_ _8992_/A _8761_/A VGND VGND VPWR VPWR mgmt_gpio_out[15] sky130_fd_sc_hd__ebufn_8
XFILLER_82_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7943_ _8636_/A _7943_/B VGND VGND VPWR VPWR _7944_/A sky130_fd_sc_hd__or2_1
XFILLER_82_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7874_ _8238_/A _8226_/C VGND VGND VPWR VPWR _8239_/B sky130_fd_sc_hd__or2_2
Xclkbuf_3_7_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A VGND VGND VPWR VPWR _9664_/CLK sky130_fd_sc_hd__clkbuf_2
X_9613_ _9613_/CLK _9613_/D _9646_/SET_B VGND VGND VPWR VPWR _9613_/Q sky130_fd_sc_hd__dfrtp_1
X_6825_ _9495_/Q VGND VGND VPWR VPWR _6825_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_23_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6756_ _9356_/Q VGND VGND VPWR VPWR _6756_/Y sky130_fd_sc_hd__clkinv_2
X_9544_ _9768_/CLK _9544_/D _4628_/A VGND VGND VPWR VPWR _9544_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5707_ _9252_/Q VGND VGND VPWR VPWR _7476_/A sky130_fd_sc_hd__inv_2
XFILLER_50_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9475_ _9687_/CLK _9475_/D _9528_/SET_B VGND VGND VPWR VPWR _9475_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_164_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6687_ _9179_/Q VGND VGND VPWR VPWR _6687_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_12_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5638_ _9282_/Q _5634_/A _8840_/X _5634_/Y VGND VGND VPWR VPWR _9282_/D sky130_fd_sc_hd__a22o_1
X_8426_ _8476_/A _8539_/A VGND VGND VPWR VPWR _8601_/D sky130_fd_sc_hd__or2_2
XFILLER_12_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8357_ _8357_/A _8658_/B VGND VGND VPWR VPWR _8573_/C sky130_fd_sc_hd__or2_1
X_5569_ _9330_/Q _5566_/A _5965_/B1 _5566_/Y VGND VGND VPWR VPWR _9330_/D sky130_fd_sc_hd__a22o_1
X_7308_ _7308_/A _7308_/B _7308_/C _7308_/D VGND VGND VPWR VPWR _7309_/C sky130_fd_sc_hd__and4_1
X_8288_ _8340_/C _8390_/B _8340_/B _8287_/X VGND VGND VPWR VPWR _8288_/X sky130_fd_sc_hd__a31o_1
XFILLER_144_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7239_ _6246_/Y _5728_/X _6303_/Y _7040_/A _7238_/X VGND VGND VPWR VPWR _7242_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_77_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4940_ _9092_/Q VGND VGND VPWR VPWR _6022_/A sky130_fd_sc_hd__inv_2
X_4871_ _9756_/Q VGND VGND VPWR VPWR _4871_/Y sky130_fd_sc_hd__inv_2
XFILLER_177_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6610_ _9349_/Q VGND VGND VPWR VPWR _8765_/A sky130_fd_sc_hd__clkinv_8
X_7590_ _7590_/A _7590_/B _7590_/C _7590_/D VGND VGND VPWR VPWR _7590_/Y sky130_fd_sc_hd__nand4_4
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6541_ _7703_/A _5949_/B _6538_/Y _5178_/B _6540_/X VGND VGND VPWR VPWR _6541_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_20_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9260_ _9601_/CLK _9260_/D _9295_/SET_B VGND VGND VPWR VPWR _9260_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_145_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6472_ _6467_/Y _5829_/B _6468_/Y _5872_/B _6471_/X VGND VGND VPWR VPWR _6473_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_161_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5423_ _9431_/Q _5422_/A _8846_/X _5422_/Y VGND VGND VPWR VPWR _9431_/D sky130_fd_sc_hd__a22o_1
X_9191_ _9378_/CLK _9191_/D _9646_/SET_B VGND VGND VPWR VPWR _9191_/Q sky130_fd_sc_hd__dfstp_1
X_8211_ _8341_/B _8264_/B VGND VGND VPWR VPWR _8312_/D sky130_fd_sc_hd__or2_2
Xoutput234 _8798_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[33] sky130_fd_sc_hd__buf_2
Xoutput223 _8778_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[23] sky130_fd_sc_hd__buf_2
X_5354_ _9476_/Q _5346_/A _8916_/A1 _5346_/Y VGND VGND VPWR VPWR _9476_/D sky130_fd_sc_hd__a22o_1
Xoutput212 _8758_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[13] sky130_fd_sc_hd__buf_2
X_8142_ _8213_/A _8550_/A VGND VGND VPWR VPWR _8575_/A sky130_fd_sc_hd__nor2_1
Xoutput245 _8750_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[9] sky130_fd_sc_hd__buf_2
Xoutput267 _9722_/Q VGND VGND VPWR VPWR pll_div[1] sky130_fd_sc_hd__buf_2
Xoutput256 _7014_/A VGND VGND VPWR VPWR pad_flash_io0_ieb sky130_fd_sc_hd__buf_2
X_5285_ _9523_/Q _5280_/A _8842_/X _5280_/Y VGND VGND VPWR VPWR _9523_/D sky130_fd_sc_hd__a22o_1
X_8073_ _8713_/A _8540_/A VGND VGND VPWR VPWR _8704_/A sky130_fd_sc_hd__or2_1
XFILLER_141_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput278 _9744_/Q VGND VGND VPWR VPWR pll_trim[12] sky130_fd_sc_hd__buf_2
Xoutput289 _9754_/Q VGND VGND VPWR VPWR pll_trim[22] sky130_fd_sc_hd__buf_2
XFILLER_101_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7024_ _9246_/Q _9245_/Q _7111_/C _7075_/A VGND VGND VPWR VPWR _7025_/A sky130_fd_sc_hd__or4_1
XFILLER_114_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8975_ _8742_/X _8728_/X _8975_/S VGND VGND VPWR VPWR _8975_/X sky130_fd_sc_hd__mux2_2
XFILLER_82_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7926_ _8305_/A _8270_/B _7925_/Y VGND VGND VPWR VPWR _7927_/B sky130_fd_sc_hd__o21ai_1
XFILLER_36_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7857_ _8496_/A _8260_/A VGND VGND VPWR VPWR _7858_/A sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_4_csclk _9329_/CLK VGND VGND VPWR VPWR _9380_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_168_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6808_ _6808_/A VGND VGND VPWR VPWR _6808_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_168_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7788_ _7903_/C _7823_/A _7787_/X VGND VGND VPWR VPWR _8528_/B sky130_fd_sc_hd__o21ai_2
XFILLER_11_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9527_ _9527_/CLK _9527_/D _9528_/SET_B VGND VGND VPWR VPWR _9527_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_139_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6739_ _6737_/Y _5534_/B _6738_/Y _5583_/B VGND VGND VPWR VPWR _6739_/X sky130_fd_sc_hd__o22a_1
XFILLER_139_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9458_ _9789_/CLK _9458_/D _9647_/SET_B VGND VGND VPWR VPWR _9458_/Q sky130_fd_sc_hd__dfrtp_1
X_8409_ _8137_/B _8401_/B _8406_/X _8408_/Y VGND VGND VPWR VPWR _8409_/X sky130_fd_sc_hd__o211a_1
XFILLER_155_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9389_ _9775_/CLK _9389_/D _7011_/B VGND VGND VPWR VPWR _9389_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_155_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5070_ _8965_/X _9663_/Q _5078_/S VGND VGND VPWR VPWR _5071_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8760_ _8760_/A VGND VGND VPWR VPWR _8760_/X sky130_fd_sc_hd__clkbuf_1
X_5972_ _9099_/Q _5970_/A _8845_/X _5970_/Y VGND VGND VPWR VPWR _9099_/D sky130_fd_sc_hd__a22o_1
XFILLER_92_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4923_ _4914_/Y _5420_/B _4916_/Y _5382_/B _4922_/X VGND VGND VPWR VPWR _4934_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7711_ _7711_/A VGND VGND VPWR VPWR _7713_/B sky130_fd_sc_hd__inv_2
X_8691_ _8713_/A _8689_/X _8635_/Y _8690_/Y VGND VGND VPWR VPWR _8691_/Y sky130_fd_sc_hd__o211ai_2
X_7642_ _6896_/Y _7471_/X _7326_/A _7473_/X _7641_/X VGND VGND VPWR VPWR _7643_/D
+ sky130_fd_sc_hd__o221a_1
X_4854_ _4846_/Y _5267_/B _4848_/Y _5442_/B _4853_/X VGND VGND VPWR VPWR _4864_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_178_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7573_ _6196_/Y _7408_/X _6230_/Y _7410_/X VGND VGND VPWR VPWR _7573_/X sky130_fd_sc_hd__o22a_1
X_4785_ _4900_/B _4843_/B VGND VGND VPWR VPWR _5941_/B sky130_fd_sc_hd__or2_4
XFILLER_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9312_ _9534_/CLK _9312_/D _9647_/SET_B VGND VGND VPWR VPWR _9312_/Q sky130_fd_sc_hd__dfstp_1
X_6524_ _6522_/Y _5602_/B _8743_/A _5045_/B VGND VGND VPWR VPWR _6524_/X sky130_fd_sc_hd__o22a_1
X_9243_ _9789_/CLK _9243_/D _9647_/SET_B VGND VGND VPWR VPWR _9243_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6455_ _6455_/A VGND VGND VPWR VPWR _8808_/B sky130_fd_sc_hd__clkinv_4
XFILLER_118_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5406_ _5406_/A VGND VGND VPWR VPWR _5406_/Y sky130_fd_sc_hd__inv_2
X_9174_ _9280_/CLK _9174_/D _9757_/SET_B VGND VGND VPWR VPWR _9174_/Q sky130_fd_sc_hd__dfrtp_1
X_6386_ input7/X VGND VGND VPWR VPWR _6386_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8125_ _8213_/A _8401_/A VGND VGND VPWR VPWR _8571_/A sky130_fd_sc_hd__nor2_1
X_5337_ _5337_/A VGND VGND VPWR VPWR _5338_/A sky130_fd_sc_hd__clkbuf_2
X_5268_ _5268_/A VGND VGND VPWR VPWR _5269_/A sky130_fd_sc_hd__buf_2
X_8056_ _8389_/A _8168_/A VGND VGND VPWR VPWR _8536_/A sky130_fd_sc_hd__or2_1
XFILLER_102_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7007_ _4952_/Y _4953_/Y _6023_/Y _9051_/Q _7008_/A VGND VGND VPWR VPWR _9051_/D
+ sky130_fd_sc_hd__a32o_1
X_5199_ _9580_/Q _5193_/Y _8955_/X _5193_/A VGND VGND VPWR VPWR _9580_/D sky130_fd_sc_hd__o22a_1
XFILLER_141_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8958_ _9090_/Q _9092_/Q _9091_/Q VGND VGND VPWR VPWR _8958_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7909_ _8077_/A _8239_/B _7877_/X _7907_/X _8303_/A VGND VGND VPWR VPWR _7909_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8889_ _8888_/X _9145_/Q _9054_/Q VGND VGND VPWR VPWR _8889_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4570_ _9752_/Q _4566_/A _5963_/B1 _4566_/Y VGND VGND VPWR VPWR _9752_/D sky130_fd_sc_hd__a22o_1
XFILLER_162_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6240_ _9507_/Q VGND VGND VPWR VPWR _6240_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6171_ _9534_/Q VGND VGND VPWR VPWR _6171_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5122_ _5122_/A VGND VGND VPWR VPWR _5123_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_111_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_opt_6_0_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR clkbuf_opt_6_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_16
X_5053_ _9669_/Q _5047_/A _8955_/A1 _5047_/Y VGND VGND VPWR VPWR _9669_/D sky130_fd_sc_hd__a22o_1
X_8812_ _8812_/A _8813_/B VGND VGND VPWR VPWR _9061_/D sky130_fd_sc_hd__nor2_1
XFILLER_1_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5955_ _9110_/Q _5951_/A _8925_/A1 _5951_/Y VGND VGND VPWR VPWR _9110_/D sky130_fd_sc_hd__a22o_1
X_8743_ _8743_/A VGND VGND VPWR VPWR _8744_/A sky130_fd_sc_hd__clkbuf_1
X_8674_ _8674_/A _8674_/B VGND VGND VPWR VPWR _8675_/B sky130_fd_sc_hd__or2_1
X_5886_ _5849_/X _8891_/X _8924_/X _9147_/Q VGND VGND VPWR VPWR _9147_/D sky130_fd_sc_hd__o22a_1
X_4906_ _4906_/A VGND VGND VPWR VPWR _4906_/Y sky130_fd_sc_hd__inv_2
X_7625_ _7625_/A _7625_/B _7625_/C _7625_/D VGND VGND VPWR VPWR _7626_/D sky130_fd_sc_hd__and4_1
X_4837_ _4919_/A _4911_/A VGND VGND VPWR VPWR _5232_/B sky130_fd_sc_hd__or2_4
XFILLER_193_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7556_ _6276_/Y _7400_/X _6309_/Y _7405_/X _7555_/X VGND VGND VPWR VPWR _7572_/A
+ sky130_fd_sc_hd__o221a_1
X_4768_ _7121_/A _5610_/B _4761_/Y _5829_/B _4767_/X VGND VGND VPWR VPWR _4790_/B
+ sky130_fd_sc_hd__o221a_1
X_4699_ _9133_/Q VGND VGND VPWR VPWR _4699_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_119_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7487_ _6818_/Y _7427_/X _6895_/Y _5699_/X VGND VGND VPWR VPWR _7487_/X sky130_fd_sc_hd__o22a_1
X_6507_ _8755_/A _5757_/B _6503_/Y _5488_/B _6506_/X VGND VGND VPWR VPWR _6526_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_136_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9226_ _9440_/CLK _9226_/D _9685_/SET_B VGND VGND VPWR VPWR _9226_/Q sky130_fd_sc_hd__dfrtp_1
X_6438_ _6438_/A VGND VGND VPWR VPWR _6438_/Y sky130_fd_sc_hd__inv_2
XFILLER_161_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9157_ _9378_/CLK _9157_/D _9646_/SET_B VGND VGND VPWR VPWR _9157_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_22_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR _9601_/CLK sky130_fd_sc_hd__clkbuf_16
X_8108_ _8108_/A VGND VGND VPWR VPWR _8640_/A sky130_fd_sc_hd__buf_6
XFILLER_121_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6369_ _9202_/Q VGND VGND VPWR VPWR _6369_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9088_ _9089_/CLK _9088_/D _5998_/X VGND VGND VPWR VPWR _9088_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_152_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8039_ _8039_/A _8416_/A VGND VGND VPWR VPWR _8041_/A sky130_fd_sc_hd__nand2_1
XFILLER_75_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_37_csclk clkbuf_2_1_0_csclk/X VGND VGND VPWR VPWR _9639_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_44_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_mgmt_gpio_in[4] mgmt_gpio_in[4] VGND VGND VPWR VPWR clkbuf_0_mgmt_gpio_in[4]/X
+ sky130_fd_sc_hd__clkbuf_16
XPHY_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_8 _7287_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5740_ _5740_/A VGND VGND VPWR VPWR _9246_/D sky130_fd_sc_hd__inv_2
XFILLER_175_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5671_ _5671_/A _5671_/B VGND VGND VPWR VPWR _5672_/A sky130_fd_sc_hd__or2_1
X_7410_ _7410_/A VGND VGND VPWR VPWR _7410_/X sky130_fd_sc_hd__buf_6
XFILLER_30_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8390_ _8518_/B _8390_/B VGND VGND VPWR VPWR _8544_/C sky130_fd_sc_hd__or2_1
X_4622_ _6158_/A _4917_/A VGND VGND VPWR VPWR _4623_/B sky130_fd_sc_hd__or2_2
XFILLER_128_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7341_ _6640_/Y _7068_/A _6725_/Y _7105_/X VGND VGND VPWR VPWR _7341_/X sky130_fd_sc_hd__o22a_2
X_4553_ _4669_/A _8932_/X _8946_/X _4729_/B VGND VGND VPWR VPWR _4925_/A sky130_fd_sc_hd__or4_4
X_7272_ _6078_/Y _7095_/X _6122_/Y _7068_/D _7271_/X VGND VGND VPWR VPWR _7277_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_116_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4484_ _9787_/Q _4466_/A _8930_/A1 _4466_/Y VGND VGND VPWR VPWR _9787_/D sky130_fd_sc_hd__a22o_1
X_9011_ _9590_/Q _8799_/A VGND VGND VPWR VPWR mgmt_gpio_out[34] sky130_fd_sc_hd__ebufn_8
XFILLER_116_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6223_ _6218_/Y _5949_/B _6219_/Y _4841_/X _6222_/X VGND VGND VPWR VPWR _6236_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6154_ _9352_/Q VGND VGND VPWR VPWR _6154_/Y sky130_fd_sc_hd__clkinv_2
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6085_ _6085_/A VGND VGND VPWR VPWR _6085_/Y sky130_fd_sc_hd__inv_2
X_5105_ _9643_/Q _5102_/A _5965_/B1 _5102_/Y VGND VGND VPWR VPWR _9643_/D sky130_fd_sc_hd__a22o_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5036_ _5981_/B VGND VGND VPWR VPWR _5985_/B sky130_fd_sc_hd__inv_2
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater364 _8841_/X VGND VGND VPWR VPWR _5965_/B1 sky130_fd_sc_hd__buf_12
Xrepeater375 _4628_/A VGND VGND VPWR VPWR _9685_/SET_B sky130_fd_sc_hd__buf_12
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6987_ _8810_/A _8809_/A _6974_/A VGND VGND VPWR VPWR _9066_/D sky130_fd_sc_hd__o21ai_1
X_9775_ _9775_/CLK _9775_/D _7011_/B VGND VGND VPWR VPWR _9775_/Q sky130_fd_sc_hd__dfstp_1
X_5938_ _6147_/B _7001_/B VGND VGND VPWR VPWR _5938_/Y sky130_fd_sc_hd__nor2_1
X_8726_ _8077_/A _8246_/B _8243_/A _8314_/X _8504_/C VGND VGND VPWR VPWR _8727_/B
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_193_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5869_ _9161_/Q _5866_/A _8841_/X _5866_/Y VGND VGND VPWR VPWR _9161_/D sky130_fd_sc_hd__a22o_1
X_8657_ _8657_/A _8657_/B _8657_/C _8657_/D VGND VGND VPWR VPWR _8696_/C sky130_fd_sc_hd__or4_2
X_8588_ _8720_/B _8588_/B _8705_/A _8681_/A VGND VGND VPWR VPWR _8588_/X sky130_fd_sc_hd__or4_1
XFILLER_139_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7608_ _7608_/A _7608_/B _7608_/C _7608_/D VGND VGND VPWR VPWR _7608_/Y sky130_fd_sc_hd__nand4_4
XFILLER_193_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7539_ _6463_/Y _7419_/X _6403_/Y _7421_/X VGND VGND VPWR VPWR _7539_/X sky130_fd_sc_hd__o22a_1
XFILLER_193_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9209_ _9652_/CLK _9209_/D _9646_/SET_B VGND VGND VPWR VPWR _9209_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_134_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput101 sram_ro_data[17] VGND VGND VPWR VPWR _6806_/A sky130_fd_sc_hd__clkbuf_1
Xinput145 wb_adr_i[21] VGND VGND VPWR VPWR _7832_/A sky130_fd_sc_hd__buf_2
Xinput134 wb_adr_i[11] VGND VGND VPWR VPWR _7771_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_88_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput112 sram_ro_data[27] VGND VGND VPWR VPWR _6561_/A sky130_fd_sc_hd__clkbuf_1
Xinput123 sram_ro_data[8] VGND VGND VPWR VPWR _4892_/A sky130_fd_sc_hd__clkbuf_1
Xinput178 wb_dat_i[21] VGND VGND VPWR VPWR _7746_/B sky130_fd_sc_hd__clkbuf_1
Xinput167 wb_dat_i[11] VGND VGND VPWR VPWR _7743_/B2 sky130_fd_sc_hd__clkbuf_1
Xinput156 wb_adr_i[31] VGND VGND VPWR VPWR _5931_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_76_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput189 wb_dat_i[31] VGND VGND VPWR VPWR _7751_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_91_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7890_ _7890_/A VGND VGND VPWR VPWR _8305_/B sky130_fd_sc_hd__buf_4
X_6910_ _9668_/Q VGND VGND VPWR VPWR _6910_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6841_ _6839_/Y _4558_/B _6840_/Y _5450_/B VGND VGND VPWR VPWR _6841_/X sky130_fd_sc_hd__o22a_1
X_9560_ _9776_/CLK _9560_/D _4628_/A VGND VGND VPWR VPWR _9560_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8511_ _8282_/C _8566_/B _8587_/A _8673_/A VGND VGND VPWR VPWR _8512_/D sky130_fd_sc_hd__a211o_1
X_6772_ _9116_/Q VGND VGND VPWR VPWR _6772_/Y sky130_fd_sc_hd__inv_2
XFILLER_148_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5723_ _7104_/A _7098_/C VGND VGND VPWR VPWR _7041_/A sky130_fd_sc_hd__or2_2
X_9491_ _9493_/CLK _9491_/D _4628_/A VGND VGND VPWR VPWR _9491_/Q sky130_fd_sc_hd__dfstp_1
X_8442_ _7896_/A _8498_/A _8624_/B _8013_/B VGND VGND VPWR VPWR _8444_/A sky130_fd_sc_hd__o22ai_1
X_5654_ _5649_/B _5751_/C _5647_/A _5651_/B VGND VGND VPWR VPWR _5654_/X sky130_fd_sc_hd__o31a_1
X_8373_ _8373_/A _8693_/B VGND VGND VPWR VPWR _8582_/A sky130_fd_sc_hd__or2_2
X_4605_ _9731_/Q _4604_/A _8844_/X _4604_/Y VGND VGND VPWR VPWR _9731_/D sky130_fd_sc_hd__a22o_1
XFILLER_163_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5585_ _5585_/A VGND VGND VPWR VPWR _5585_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7324_ _6874_/Y _7118_/X _6892_/Y _7048_/C VGND VGND VPWR VPWR _7324_/X sky130_fd_sc_hd__o22a_1
XFILLER_190_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4536_ _6111_/A _4929_/A VGND VGND VPWR VPWR _4537_/B sky130_fd_sc_hd__or2_2
XFILLER_131_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7255_ _7255_/A _7255_/B _7255_/C _7255_/D VGND VGND VPWR VPWR _7265_/B sky130_fd_sc_hd__and4_1
XFILLER_116_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4467_ _9790_/Q _4466_/A _8845_/X _4466_/Y VGND VGND VPWR VPWR _9790_/D sky130_fd_sc_hd__a22o_1
X_7186_ _6582_/Y _7059_/B _8797_/A _7068_/C _7185_/X VGND VGND VPWR VPWR _7189_/C
+ sky130_fd_sc_hd__o221a_2
X_6206_ input9/X VGND VGND VPWR VPWR _6206_/Y sky130_fd_sc_hd__inv_2
X_6137_ _6132_/Y _6322_/A _6133_/Y _5545_/B _6136_/Y VGND VGND VPWR VPWR _6144_/C
+ sky130_fd_sc_hd__o221a_2
XFILLER_133_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6068_ _9371_/Q VGND VGND VPWR VPWR _6068_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_85_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5019_ _9692_/Q _5015_/A _8925_/A1 _5015_/Y VGND VGND VPWR VPWR _9692_/D sky130_fd_sc_hd__a22o_1
XFILLER_73_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9758_ _9758_/CLK _9758_/D _7011_/B VGND VGND VPWR VPWR _9758_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_41_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8709_ _8709_/A _8709_/B _8709_/C _8709_/D VGND VGND VPWR VPWR _8738_/A sky130_fd_sc_hd__or4_1
X_9689_ _9695_/CLK _9689_/D _9779_/SET_B VGND VGND VPWR VPWR _9689_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_21_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5370_ _9466_/Q _5368_/A _5964_/B1 _5368_/Y VGND VGND VPWR VPWR _9466_/D sky130_fd_sc_hd__a22o_1
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7040_ _7040_/A _7040_/B _7040_/C _7040_/D VGND VGND VPWR VPWR _7079_/C sky130_fd_sc_hd__and4_1
XFILLER_141_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8991_ _8991_/A _8759_/A VGND VGND VPWR VPWR mgmt_gpio_out[14] sky130_fd_sc_hd__ebufn_2
XFILLER_67_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7942_ _8651_/A _8562_/A _7942_/C VGND VGND VPWR VPWR _7943_/B sky130_fd_sc_hd__or3_1
XFILLER_94_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9612_ _9788_/CLK _9612_/D _9646_/SET_B VGND VGND VPWR VPWR _9612_/Q sky130_fd_sc_hd__dfrtp_1
X_7873_ _7873_/A VGND VGND VPWR VPWR _8238_/A sky130_fd_sc_hd__buf_2
XFILLER_168_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6824_ _9485_/Q VGND VGND VPWR VPWR _6824_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6755_ _9153_/Q VGND VGND VPWR VPWR _6755_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9543_ _9768_/CLK _9543_/D _4628_/A VGND VGND VPWR VPWR _9543_/Q sky130_fd_sc_hd__dfstp_1
X_9474_ _9687_/CLK _9474_/D _9528_/SET_B VGND VGND VPWR VPWR _9474_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_10_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5706_ _7406_/B _5704_/Y _9055_/Q _5705_/X VGND VGND VPWR VPWR _9253_/D sky130_fd_sc_hd__a31o_1
XFILLER_176_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6686_ _9366_/Q VGND VGND VPWR VPWR _6686_/Y sky130_fd_sc_hd__inv_2
XFILLER_148_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8425_ _8688_/A _8631_/A _8425_/C VGND VGND VPWR VPWR _8427_/A sky130_fd_sc_hd__or3_1
XFILLER_31_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5637_ _9283_/Q _5634_/A _8841_/X _5634_/Y VGND VGND VPWR VPWR _9283_/D sky130_fd_sc_hd__a22o_1
XFILLER_163_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8356_ _8356_/A _8356_/B _8571_/C _8677_/A VGND VGND VPWR VPWR _8360_/A sky130_fd_sc_hd__or4_1
X_5568_ _9331_/Q _5566_/A _5964_/B1 _5566_/Y VGND VGND VPWR VPWR _9331_/D sky130_fd_sc_hd__a22o_1
X_8287_ _8713_/A _8287_/B VGND VGND VPWR VPWR _8287_/X sky130_fd_sc_hd__or2_1
XFILLER_117_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4519_ _4931_/A _6158_/A _5259_/A VGND VGND VPWR VPWR _4520_/S sky130_fd_sc_hd__or3_1
X_7307_ _4918_/Y _7124_/X _4763_/Y _7068_/B _7306_/X VGND VGND VPWR VPWR _7308_/D
+ sky130_fd_sc_hd__o221a_1
X_7238_ _7238_/A _7392_/B VGND VGND VPWR VPWR _7238_/X sky130_fd_sc_hd__or2_1
X_5499_ _9379_/Q _5498_/A _8846_/X _5498_/Y VGND VGND VPWR VPWR _9379_/D sky130_fd_sc_hd__a22o_1
XFILLER_144_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7169_ _6687_/Y _7040_/D _6737_/Y _7110_/X _7168_/X VGND VGND VPWR VPWR _7176_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_58_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4870_ _6158_/A _4900_/B VGND VGND VPWR VPWR _4870_/X sky130_fd_sc_hd__or2_4
XFILLER_45_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6540_ _4629_/C _8955_/S _6539_/Y _5941_/B VGND VGND VPWR VPWR _6540_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_60_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6471_ _6469_/Y _4524_/B _6470_/Y _4870_/X VGND VGND VPWR VPWR _6471_/X sky130_fd_sc_hd__o22a_2
X_5422_ _5422_/A VGND VGND VPWR VPWR _5422_/Y sky130_fd_sc_hd__inv_2
XFILLER_145_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9190_ _9352_/CLK _9190_/D _9646_/SET_B VGND VGND VPWR VPWR _9190_/Q sky130_fd_sc_hd__dfstp_1
X_8210_ _8210_/A VGND VGND VPWR VPWR _8260_/B sky130_fd_sc_hd__buf_4
Xoutput235 _8800_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[34] sky130_fd_sc_hd__buf_2
Xoutput224 _8780_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[24] sky130_fd_sc_hd__buf_2
X_5353_ _9477_/Q _5346_/A _8840_/X _5346_/Y VGND VGND VPWR VPWR _9477_/D sky130_fd_sc_hd__a22o_1
Xoutput213 _8760_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[14] sky130_fd_sc_hd__buf_2
X_8141_ _8550_/A _8378_/B VGND VGND VPWR VPWR _8362_/A sky130_fd_sc_hd__nor2_1
XFILLER_99_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput268 _9723_/Q VGND VGND VPWR VPWR pll_div[2] sky130_fd_sc_hd__buf_2
Xoutput257 _7014_/Y VGND VGND VPWR VPWR pad_flash_io0_oeb sky130_fd_sc_hd__buf_2
Xoutput246 _8824_/X VGND VGND VPWR VPWR mgmt_gpio_out[0] sky130_fd_sc_hd__buf_2
X_5284_ _9524_/Q _5280_/A _8925_/A1 _5280_/Y VGND VGND VPWR VPWR _9524_/D sky130_fd_sc_hd__a22o_1
X_8072_ _8305_/A _8437_/B VGND VGND VPWR VPWR _8540_/A sky130_fd_sc_hd__nor2_1
XFILLER_114_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput279 _9745_/Q VGND VGND VPWR VPWR pll_trim[13] sky130_fd_sc_hd__buf_2
XFILLER_101_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7023_ _9248_/Q _9247_/Q VGND VGND VPWR VPWR _7111_/C sky130_fd_sc_hd__or2_2
XFILLER_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8974_ _8725_/Y _8697_/X _8975_/S VGND VGND VPWR VPWR _8974_/X sky130_fd_sc_hd__mux2_2
X_7925_ _8599_/A _7925_/B VGND VGND VPWR VPWR _7925_/Y sky130_fd_sc_hd__nor2_1
XFILLER_82_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7856_ _8525_/A _7894_/B _7959_/A _8528_/A VGND VGND VPWR VPWR _8260_/A sky130_fd_sc_hd__or4_4
XFILLER_70_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6807_ _9786_/Q VGND VGND VPWR VPWR _6807_/Y sky130_fd_sc_hd__inv_4
X_9526_ _9527_/CLK _9526_/D _9528_/SET_B VGND VGND VPWR VPWR _9526_/Q sky130_fd_sc_hd__dfrtp_1
X_7787_ _7959_/A _7787_/B VGND VGND VPWR VPWR _7787_/X sky130_fd_sc_hd__or2_1
X_4999_ _6040_/A VGND VGND VPWR VPWR _5000_/A sky130_fd_sc_hd__clkbuf_1
X_6738_ _9314_/Q VGND VGND VPWR VPWR _6738_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9457_ _9483_/CLK _9457_/D _9528_/SET_B VGND VGND VPWR VPWR _9457_/Q sky130_fd_sc_hd__dfrtp_1
X_6669_ _6669_/A VGND VGND VPWR VPWR _6669_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8408_ _8607_/B _8573_/A VGND VGND VPWR VPWR _8408_/Y sky130_fd_sc_hd__nor2_1
X_9388_ _9775_/CLK _9388_/D _7011_/B VGND VGND VPWR VPWR _9388_/Q sky130_fd_sc_hd__dfrtp_1
X_8339_ _8651_/A _8672_/C VGND VGND VPWR VPWR _8705_/A sky130_fd_sc_hd__or2_2
XFILLER_105_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5971_ _9100_/Q _5970_/A _8846_/X _5970_/Y VGND VGND VPWR VPWR _9100_/D sky130_fd_sc_hd__a22o_1
X_8690_ _8714_/C VGND VGND VPWR VPWR _8690_/Y sky130_fd_sc_hd__inv_2
X_4922_ _4918_/Y _5480_/B _4920_/Y _5518_/B VGND VGND VPWR VPWR _4922_/X sky130_fd_sc_hd__o22a_2
X_7710_ _9083_/Q _9082_/Q _7711_/A VGND VGND VPWR VPWR _7710_/X sky130_fd_sc_hd__o21a_1
XFILLER_178_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7641_ _6812_/Y _7475_/X _6928_/Y _7477_/X VGND VGND VPWR VPWR _7641_/X sky130_fd_sc_hd__o22a_1
X_4853_ _4850_/Y _5355_/B _4852_/Y _4524_/B VGND VGND VPWR VPWR _4853_/X sky130_fd_sc_hd__o22a_1
XFILLER_193_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7572_ _7572_/A _7572_/B _7572_/C _7572_/D VGND VGND VPWR VPWR _7572_/Y sky130_fd_sc_hd__nand4_4
X_4784_ _9114_/Q VGND VGND VPWR VPWR _4784_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9311_ _9789_/CLK _9311_/D _9685_/SET_B VGND VGND VPWR VPWR _9311_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_119_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_opt_2_0_csclk clkbuf_2_1_0_csclk/X VGND VGND VPWR VPWR clkbuf_opt_2_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_16
X_6523_ _9670_/Q VGND VGND VPWR VPWR _8743_/A sky130_fd_sc_hd__inv_4
X_9242_ _9789_/CLK _9242_/D _9647_/SET_B VGND VGND VPWR VPWR _9242_/Q sky130_fd_sc_hd__dfstp_1
X_6454_ _6449_/Y _4590_/B _6450_/Y _6135_/A _6453_/X VGND VGND VPWR VPWR _6473_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_106_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5405_ _5405_/A VGND VGND VPWR VPWR _5406_/A sky130_fd_sc_hd__clkbuf_2
X_6385_ _6385_/A VGND VGND VPWR VPWR _6385_/Y sky130_fd_sc_hd__inv_2
X_9173_ _9280_/CLK _9173_/D _9757_/SET_B VGND VGND VPWR VPWR _9173_/Q sky130_fd_sc_hd__dfrtp_1
X_8124_ _8114_/Y _8115_/Y _8115_/Y _8390_/B _8123_/X VGND VGND VPWR VPWR _8127_/B
+ sky130_fd_sc_hd__a221o_1
X_5336_ _5671_/A _5336_/B VGND VGND VPWR VPWR _5337_/A sky130_fd_sc_hd__or2_1
XFILLER_141_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5267_ _5545_/A _5267_/B VGND VGND VPWR VPWR _5268_/A sky130_fd_sc_hd__or2_1
X_8055_ _8055_/A _8708_/C VGND VGND VPWR VPWR _8057_/A sky130_fd_sc_hd__nor2_1
XFILLER_114_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7006_ _9708_/Q _5993_/B _9048_/Q _9052_/Q VGND VGND VPWR VPWR _9052_/D sky130_fd_sc_hd__a31o_1
X_5198_ _9581_/Q _5193_/Y _8923_/X _5193_/A VGND VGND VPWR VPWR _9581_/D sky130_fd_sc_hd__o22a_1
X_8957_ _5007_/S _6022_/B _8957_/S VGND VGND VPWR VPWR _8957_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7908_ _8521_/B _8232_/B VGND VGND VPWR VPWR _8303_/A sky130_fd_sc_hd__or2_1
XFILLER_43_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8888_ _7309_/Y _9627_/Q _8959_/S VGND VGND VPWR VPWR _8888_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7839_ _7839_/A VGND VGND VPWR VPWR _8195_/A sky130_fd_sc_hd__inv_2
XFILLER_34_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9509_ _9509_/CLK _9509_/D _9528_/SET_B VGND VGND VPWR VPWR _9509_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_149_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6170_ _9292_/Q VGND VGND VPWR VPWR _6170_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_130_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_3_csclk _9329_/CLK VGND VGND VPWR VPWR _9771_/CLK sky130_fd_sc_hd__clkbuf_16
X_5121_ _5259_/A _5121_/B VGND VGND VPWR VPWR _5122_/A sky130_fd_sc_hd__or2_1
XFILLER_111_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5052_ _9670_/Q _5047_/A _8929_/A1 _5047_/Y VGND VGND VPWR VPWR _9670_/D sky130_fd_sc_hd__a22o_1
X_8811_ _8811_/A _8813_/B VGND VGND VPWR VPWR _9062_/D sky130_fd_sc_hd__nor2_1
XFILLER_92_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9791_ _9791_/CLK _9791_/D _9633_/SET_B VGND VGND VPWR VPWR _9791_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_37_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8742_ _8729_/Y _8723_/Y _8731_/X _8741_/X VGND VGND VPWR VPWR _8742_/X sky130_fd_sc_hd__a31o_1
XFILLER_92_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5954_ _9111_/Q _5951_/A _8844_/X _5951_/Y VGND VGND VPWR VPWR _9111_/D sky130_fd_sc_hd__a22o_1
XFILLER_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8673_ _8673_/A _8706_/A _8673_/C _8707_/B VGND VGND VPWR VPWR _8673_/X sky130_fd_sc_hd__or4_2
X_4905_ _4897_/Y _5344_/B _4899_/Y _5404_/B _4904_/X VGND VGND VPWR VPWR _4934_/A
+ sky130_fd_sc_hd__o221a_1
X_5885_ _5849_/X _8893_/X _8924_/X _9148_/Q VGND VGND VPWR VPWR _9148_/D sky130_fd_sc_hd__o22a_1
XFILLER_33_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7624_ _4699_/Y _7471_/X _7304_/A _7473_/X _7623_/X VGND VGND VPWR VPWR _7625_/D
+ sky130_fd_sc_hd__o221a_1
X_4836_ _9554_/Q VGND VGND VPWR VPWR _4836_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7555_ _6290_/Y _7408_/X _6303_/Y _7410_/X VGND VGND VPWR VPWR _7555_/X sky130_fd_sc_hd__o22a_1
XFILLER_193_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6506_ _6504_/Y _5829_/B _6505_/Y _6134_/A VGND VGND VPWR VPWR _6506_/X sky130_fd_sc_hd__o22a_1
X_4767_ _4763_/Y _5564_/B _4765_/Y _5960_/B VGND VGND VPWR VPWR _4767_/X sky130_fd_sc_hd__o22a_1
XFILLER_146_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7486_ _6890_/Y _7415_/X _6921_/Y _7417_/X _7485_/X VGND VGND VPWR VPWR _7500_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4698_ _4698_/A VGND VGND VPWR VPWR _6165_/A sky130_fd_sc_hd__buf_12
X_9225_ _9695_/CLK _9225_/D _9779_/SET_B VGND VGND VPWR VPWR _9225_/Q sky130_fd_sc_hd__dfrtp_1
X_6437_ _6435_/Y _5110_/B _6436_/Y _5507_/B VGND VGND VPWR VPWR _6437_/X sky130_fd_sc_hd__o22a_1
XFILLER_20_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6368_ _9235_/Q VGND VGND VPWR VPWR _6368_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9156_ _9695_/CLK _9156_/D _9779_/SET_B VGND VGND VPWR VPWR _9156_/Q sky130_fd_sc_hd__dfrtp_1
X_8107_ _8218_/A _8200_/B _8218_/C VGND VGND VPWR VPWR _8108_/A sky130_fd_sc_hd__or3_1
X_5319_ _5319_/A VGND VGND VPWR VPWR _5319_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6299_ input49/X _8926_/S _6298_/Y _5818_/B VGND VGND VPWR VPWR _6299_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_29_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9087_ _9089_/CLK _9087_/D _6001_/X VGND VGND VPWR VPWR _9087_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_102_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8038_ _8521_/A _8552_/A VGND VGND VPWR VPWR _8416_/A sky130_fd_sc_hd__or2_1
XFILLER_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_9 _7287_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5670_ _9269_/Q _5662_/A _8839_/X _5662_/Y VGND VGND VPWR VPWR _9269_/D sky130_fd_sc_hd__a22o_1
XFILLER_148_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4621_ _4669_/A _8932_/X _8946_/X _8944_/X VGND VGND VPWR VPWR _4917_/A sky130_fd_sc_hd__or4_4
XFILLER_163_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4552_ _7731_/A _5062_/D _9759_/Q _8960_/X _4551_/X VGND VGND VPWR VPWR _9759_/D
+ sky130_fd_sc_hd__a32o_1
X_7340_ _6707_/Y _7059_/B _6719_/Y _7068_/C _7339_/X VGND VGND VPWR VPWR _7343_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_183_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4483_ _4483_/A VGND VGND VPWR VPWR _9788_/D sky130_fd_sc_hd__clkbuf_1
X_7271_ _6110_/Y _7097_/X _6079_/Y _7099_/X VGND VGND VPWR VPWR _7271_/X sky130_fd_sc_hd__o22a_1
X_9010_ _9010_/A _8797_/A VGND VGND VPWR VPWR mgmt_gpio_out[33] sky130_fd_sc_hd__ebufn_8
XFILLER_131_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6222_ _6220_/Y _4564_/B _6221_/Y _4893_/X VGND VGND VPWR VPWR _6222_/X sky130_fd_sc_hd__o22a_1
X_6153_ _6153_/A VGND VGND VPWR VPWR _6153_/Y sky130_fd_sc_hd__inv_2
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6084_ _9739_/Q VGND VGND VPWR VPWR _6084_/Y sky130_fd_sc_hd__inv_2
X_5104_ _9644_/Q _5102_/A _5964_/B1 _5102_/Y VGND VGND VPWR VPWR _9644_/D sky130_fd_sc_hd__a22o_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5035_ _9048_/Q _9050_/Q _9051_/Q VGND VGND VPWR VPWR _5981_/B sky130_fd_sc_hd__or3_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater365 _8841_/X VGND VGND VPWR VPWR _8955_/A1 sky130_fd_sc_hd__buf_12
Xrepeater376 _7011_/B VGND VGND VPWR VPWR _4628_/A sky130_fd_sc_hd__buf_12
XFILLER_65_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6986_ _8811_/A _8809_/A _5939_/X VGND VGND VPWR VPWR _9064_/D sky130_fd_sc_hd__o21ai_1
XFILLER_80_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9774_ _9774_/CLK _9774_/D _7011_/B VGND VGND VPWR VPWR _9774_/Q sky130_fd_sc_hd__dfrtp_1
X_5937_ _9059_/Q _5939_/B VGND VGND VPWR VPWR _7001_/B sky130_fd_sc_hd__and2_1
X_8725_ _8702_/Y _8733_/A _8712_/Y _8739_/A _8724_/Y VGND VGND VPWR VPWR _8725_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8656_ _7836_/B _7862_/Y _8518_/A _8367_/B VGND VGND VPWR VPWR _8657_/B sky130_fd_sc_hd__a31o_1
XFILLER_40_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5868_ _9162_/Q _5866_/A _8842_/X _5866_/Y VGND VGND VPWR VPWR _9162_/D sky130_fd_sc_hd__a22o_1
X_7607_ _7607_/A _7607_/B _7607_/C _7607_/D VGND VGND VPWR VPWR _7608_/D sky130_fd_sc_hd__and4_1
X_8587_ _8587_/A _8606_/B VGND VGND VPWR VPWR _8681_/A sky130_fd_sc_hd__or2_1
X_5799_ _5799_/A VGND VGND VPWR VPWR _5799_/Y sky130_fd_sc_hd__clkinv_2
X_4819_ _4816_/Y _5393_/B _4818_/Y _4623_/B VGND VGND VPWR VPWR _4819_/X sky130_fd_sc_hd__o22a_1
XFILLER_193_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7538_ _6421_/Y _7400_/X _6371_/Y _7405_/X _7537_/X VGND VGND VPWR VPWR _7554_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_31_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7469_ _4716_/Y _7461_/X _4910_/Y _7463_/X _7468_/X VGND VGND VPWR VPWR _7480_/C
+ sky130_fd_sc_hd__o221a_1
X_9208_ _9788_/CLK _9208_/D _9647_/SET_B VGND VGND VPWR VPWR _9208_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_107_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9139_ _9280_/CLK _9139_/D _9633_/SET_B VGND VGND VPWR VPWR _9139_/Q sky130_fd_sc_hd__dfrtp_1
Xinput102 sram_ro_data[18] VGND VGND VPWR VPWR _6744_/A sky130_fd_sc_hd__clkbuf_1
Xinput135 wb_adr_i[12] VGND VGND VPWR VPWR _7771_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput113 sram_ro_data[28] VGND VGND VPWR VPWR _6444_/A sky130_fd_sc_hd__clkbuf_1
Xinput124 sram_ro_data[9] VGND VGND VPWR VPWR _6808_/A sky130_fd_sc_hd__clkbuf_1
Xinput168 wb_dat_i[12] VGND VGND VPWR VPWR _7745_/B2 sky130_fd_sc_hd__clkbuf_1
Xinput146 wb_adr_i[22] VGND VGND VPWR VPWR _7781_/B sky130_fd_sc_hd__clkbuf_1
Xinput157 wb_adr_i[3] VGND VGND VPWR VPWR _8379_/D sky130_fd_sc_hd__buf_4
XFILLER_88_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput179 wb_dat_i[22] VGND VGND VPWR VPWR _7748_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_91_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6840_ _9407_/Q VGND VGND VPWR VPWR _6840_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6771_ _6766_/Y _4907_/X _6767_/Y _5458_/B _6770_/X VGND VGND VPWR VPWR _6783_/B
+ sky130_fd_sc_hd__o221a_1
X_8510_ _8510_/A _8660_/B _8660_/C VGND VGND VPWR VPWR _8603_/C sky130_fd_sc_hd__nor3_1
X_5722_ _7037_/A _7056_/B VGND VGND VPWR VPWR _7098_/C sky130_fd_sc_hd__or2_2
Xclkbuf_leaf_21_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR _9371_/CLK sky130_fd_sc_hd__clkbuf_16
X_9490_ _9545_/CLK _9490_/D _4628_/A VGND VGND VPWR VPWR _9490_/Q sky130_fd_sc_hd__dfrtp_1
X_8441_ _8441_/A _8441_/B VGND VGND VPWR VPWR _8449_/A sky130_fd_sc_hd__nand2_1
X_5653_ _5649_/B _5647_/X _5649_/A _5651_/X _5652_/Y VGND VGND VPWR VPWR _9280_/D
+ sky130_fd_sc_hd__o311a_1
X_5584_ _5584_/A VGND VGND VPWR VPWR _5585_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_136_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8372_ _8372_/A _8645_/C _8579_/C _8715_/C VGND VGND VPWR VPWR _8375_/A sky130_fd_sc_hd__or4_4
X_4604_ _4604_/A VGND VGND VPWR VPWR _4604_/Y sky130_fd_sc_hd__clkinv_2
X_7323_ _6909_/Y _7040_/D _6898_/Y _7110_/X _7322_/X VGND VGND VPWR VPWR _7330_/A
+ sky130_fd_sc_hd__o221a_2
Xclkbuf_leaf_36_csclk clkbuf_2_1_0_csclk/X VGND VGND VPWR VPWR _9791_/CLK sky130_fd_sc_hd__clkbuf_16
X_4535_ _8946_/X _8944_/X _8934_/X _4729_/D VGND VGND VPWR VPWR _4929_/A sky130_fd_sc_hd__or4_4
XFILLER_144_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7254_ _6184_/Y _7048_/D _6157_/Y _7040_/B _7253_/X VGND VGND VPWR VPWR _7255_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_104_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4466_ _4466_/A VGND VGND VPWR VPWR _4466_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_171_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6205_ _9370_/Q VGND VGND VPWR VPWR _6205_/Y sky130_fd_sc_hd__clkinv_4
X_7185_ _8795_/A _7079_/B _8759_/A _7059_/A VGND VGND VPWR VPWR _7185_/X sky130_fd_sc_hd__o22a_1
XFILLER_104_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6136_ input42/X _8930_/S input51/X _8926_/S VGND VGND VPWR VPWR _6136_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_131_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6067_ _9293_/Q VGND VGND VPWR VPWR _6067_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5018_ _9693_/Q _5015_/A _8844_/X _5015_/Y VGND VGND VPWR VPWR _9693_/D sky130_fd_sc_hd__a22o_1
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6969_ _6629_/Y _6964_/A _9023_/Q _6964_/Y VGND VGND VPWR VPWR _9023_/D sky130_fd_sc_hd__o22a_1
X_9757_ _9757_/CLK _9757_/D _9757_/SET_B VGND VGND VPWR VPWR _9757_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_53_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8708_ _8708_/A _8708_/B _8708_/C _8708_/D VGND VGND VPWR VPWR _8709_/B sky130_fd_sc_hd__or4_1
X_9688_ _9695_/CLK _9688_/D _9779_/SET_B VGND VGND VPWR VPWR _9688_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_166_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8639_ _8115_/Y _8390_/B _8595_/C _8356_/A _8572_/C VGND VGND VPWR VPWR _8677_/D
+ sky130_fd_sc_hd__a2111o_1
XFILLER_21_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8990_ _8990_/A _8757_/A VGND VGND VPWR VPWR mgmt_gpio_out[13] sky130_fd_sc_hd__ebufn_8
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7941_ _8587_/A _7941_/B VGND VGND VPWR VPWR _7942_/C sky130_fd_sc_hd__or2_1
X_7872_ _8583_/A _8189_/A _7959_/A _8528_/A VGND VGND VPWR VPWR _7873_/A sky130_fd_sc_hd__or4_4
X_9611_ _9613_/CLK _9611_/D _9646_/SET_B VGND VGND VPWR VPWR _9611_/Q sky130_fd_sc_hd__dfrtp_1
X_6823_ _9071_/Q VGND VGND VPWR VPWR _6823_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_168_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6754_ _9127_/Q VGND VGND VPWR VPWR _6754_/Y sky130_fd_sc_hd__clkinv_2
X_9542_ _9545_/CLK _9542_/D _4628_/A VGND VGND VPWR VPWR _9542_/Q sky130_fd_sc_hd__dfrtp_1
X_6685_ _9685_/Q VGND VGND VPWR VPWR _6685_/Y sky130_fd_sc_hd__clkinv_4
X_9473_ _9687_/CLK _9473_/D _9528_/SET_B VGND VGND VPWR VPWR _9473_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_148_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5705_ _5724_/B _7462_/A _5692_/A _9253_/Q VGND VGND VPWR VPWR _5705_/X sky130_fd_sc_hd__o211a_1
XFILLER_191_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5636_ _9284_/Q _5634_/A _8842_/X _5634_/Y VGND VGND VPWR VPWR _9284_/D sky130_fd_sc_hd__a22o_1
XFILLER_148_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8424_ _8168_/A _8401_/B _8423_/X VGND VGND VPWR VPWR _8425_/C sky130_fd_sc_hd__o21bai_1
XFILLER_163_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8355_ _8683_/B _8499_/B VGND VGND VPWR VPWR _8677_/A sky130_fd_sc_hd__or2_1
X_5567_ _9332_/Q _5566_/A _5963_/B1 _5566_/Y VGND VGND VPWR VPWR _9332_/D sky130_fd_sc_hd__a22o_1
X_8286_ _8585_/B _8721_/A _8286_/C VGND VGND VPWR VPWR _8287_/B sky130_fd_sc_hd__or3_1
XFILLER_117_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4518_ _9771_/Q _4517_/Y _5967_/B1 _4517_/A _8939_/X VGND VGND VPWR VPWR _9771_/D
+ sky130_fd_sc_hd__o221a_1
X_5498_ _5498_/A VGND VGND VPWR VPWR _5498_/Y sky130_fd_sc_hd__inv_2
X_7306_ _4882_/Y _7126_/X _4809_/Y _7128_/X VGND VGND VPWR VPWR _7306_/X sky130_fd_sc_hd__o22a_1
X_4449_ _9577_/Q _4449_/A1 _9786_/Q VGND VGND VPWR VPWR _8992_/A sky130_fd_sc_hd__mux2_1
XFILLER_132_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7237_ _6315_/Y _7059_/D _6276_/Y _7116_/X _7236_/X VGND VGND VPWR VPWR _7242_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_144_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7168_ _6661_/Y _7112_/X _6755_/Y _7077_/B VGND VGND VPWR VPWR _7168_/X sky130_fd_sc_hd__o22a_1
X_6119_ _6119_/A _6119_/B _6119_/C _6119_/D VGND VGND VPWR VPWR _6145_/C sky130_fd_sc_hd__and4_1
X_7099_ _7099_/A VGND VGND VPWR VPWR _7099_/X sky130_fd_sc_hd__buf_8
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6470_ _6470_/A VGND VGND VPWR VPWR _6470_/Y sky130_fd_sc_hd__inv_2
XFILLER_161_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5421_ _5421_/A VGND VGND VPWR VPWR _5422_/A sky130_fd_sc_hd__clkbuf_4
Xoutput225 _8782_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[25] sky130_fd_sc_hd__buf_2
X_5352_ _9478_/Q _5346_/A _8841_/X _5346_/Y VGND VGND VPWR VPWR _9478_/D sky130_fd_sc_hd__a22o_1
XFILLER_173_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput214 _8762_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[15] sky130_fd_sc_hd__buf_2
X_8140_ _8140_/A _8574_/A _8361_/A _8730_/A VGND VGND VPWR VPWR _8144_/A sky130_fd_sc_hd__or4_1
Xoutput236 _8833_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[35] sky130_fd_sc_hd__buf_2
X_8071_ _8202_/A _8077_/A VGND VGND VPWR VPWR _8713_/A sky130_fd_sc_hd__nor2_4
Xoutput258 _8816_/X VGND VGND VPWR VPWR pad_flash_io1_do sky130_fd_sc_hd__buf_2
Xoutput247 _8827_/X VGND VGND VPWR VPWR mgmt_gpio_out[1] sky130_fd_sc_hd__buf_2
X_5283_ _9525_/Q _5280_/A _8844_/X _5280_/Y VGND VGND VPWR VPWR _9525_/D sky130_fd_sc_hd__a22o_1
XFILLER_141_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7022_ _7022_/A _7022_/B VGND VGND VPWR VPWR _7022_/Y sky130_fd_sc_hd__nor2_2
Xoutput269 _9724_/Q VGND VGND VPWR VPWR pll_div[3] sky130_fd_sc_hd__buf_2
XFILLER_87_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8973_ _8692_/Y _8664_/X _8975_/S VGND VGND VPWR VPWR _8973_/X sky130_fd_sc_hd__mux2_2
XFILLER_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7924_ _8463_/A _7924_/B VGND VGND VPWR VPWR _7925_/B sky130_fd_sc_hd__or2_1
X_7855_ _8077_/A _8270_/B VGND VGND VPWR VPWR _8599_/A sky130_fd_sc_hd__nor2_1
XFILLER_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6806_ _6806_/A VGND VGND VPWR VPWR _6806_/Y sky130_fd_sc_hd__clkinv_2
X_9525_ _9684_/CLK _9525_/D _9685_/SET_B VGND VGND VPWR VPWR _9525_/Q sky130_fd_sc_hd__dfrtp_1
X_7786_ _7787_/B VGND VGND VPWR VPWR _7823_/A sky130_fd_sc_hd__inv_2
X_4998_ _6050_/A VGND VGND VPWR VPWR _6040_/A sky130_fd_sc_hd__buf_8
XFILLER_23_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6737_ _9348_/Q VGND VGND VPWR VPWR _6737_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9456_ _9509_/CLK _9456_/D _9528_/SET_B VGND VGND VPWR VPWR _9456_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_128_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6668_ _9382_/Q VGND VGND VPWR VPWR _6668_/Y sky130_fd_sc_hd__inv_2
X_5619_ _9295_/Q _5612_/A _8840_/X _5612_/Y VGND VGND VPWR VPWR _9295_/D sky130_fd_sc_hd__a22o_1
X_8407_ _8407_/A VGND VGND VPWR VPWR _8607_/B sky130_fd_sc_hd__inv_2
X_6599_ _9729_/Q VGND VGND VPWR VPWR _6599_/Y sky130_fd_sc_hd__inv_2
X_9387_ _9775_/CLK _9387_/D _7011_/B VGND VGND VPWR VPWR _9387_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_164_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8338_ _8338_/A VGND VGND VPWR VPWR _8338_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8269_ _8269_/A _8579_/B VGND VGND VPWR VPWR _8271_/A sky130_fd_sc_hd__or2_1
XFILLER_120_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5970_ _5970_/A VGND VGND VPWR VPWR _5970_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4921_ _4921_/A _4931_/B VGND VGND VPWR VPWR _5518_/B sky130_fd_sc_hd__or2_4
XFILLER_52_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7640_ _6909_/Y _7461_/X _6845_/Y _7463_/X _7639_/X VGND VGND VPWR VPWR _7643_/C
+ sky130_fd_sc_hd__o221a_1
X_4852_ _9762_/Q VGND VGND VPWR VPWR _4852_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7571_ _7571_/A _7571_/B _7571_/C _7571_/D VGND VGND VPWR VPWR _7572_/D sky130_fd_sc_hd__and4_2
X_4783_ _4783_/A VGND VGND VPWR VPWR _6322_/A sky130_fd_sc_hd__buf_12
X_9310_ _9789_/CLK _9310_/D _9647_/SET_B VGND VGND VPWR VPWR _9310_/Q sky130_fd_sc_hd__dfrtp_1
X_6522_ _9305_/Q VGND VGND VPWR VPWR _6522_/Y sky130_fd_sc_hd__clkinv_2
X_9241_ _9789_/CLK _9241_/D _9647_/SET_B VGND VGND VPWR VPWR _9241_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6453_ _6451_/Y _4861_/X _6452_/Y _4602_/B VGND VGND VPWR VPWR _6453_/X sky130_fd_sc_hd__o22a_2
XFILLER_133_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5404_ _5671_/A _5404_/B VGND VGND VPWR VPWR _5405_/A sky130_fd_sc_hd__or2_1
X_9172_ _9203_/CLK _9172_/D _9757_/SET_B VGND VGND VPWR VPWR _9172_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_161_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8123_ _8394_/C _7839_/A _8393_/A _8118_/X _8122_/X VGND VGND VPWR VPWR _8123_/X
+ sky130_fd_sc_hd__a41o_2
XFILLER_133_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6384_ _9752_/Q VGND VGND VPWR VPWR _6384_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5335_ _9489_/Q _5330_/A _5967_/B1 _5330_/Y VGND VGND VPWR VPWR _9489_/D sky130_fd_sc_hd__a22o_1
X_8054_ _8624_/B _8168_/A VGND VGND VPWR VPWR _8708_/C sky130_fd_sc_hd__nor2_1
XFILLER_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5266_ _9536_/Q _5261_/A _5967_/B1 _5261_/Y VGND VGND VPWR VPWR _9536_/D sky130_fd_sc_hd__a22o_1
X_7005_ _7005_/A VGND VGND VPWR VPWR _9048_/D sky130_fd_sc_hd__inv_2
XFILLER_18_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5197_ _9582_/Q _5193_/Y _8920_/X _5193_/A VGND VGND VPWR VPWR _9582_/D sky130_fd_sc_hd__o22a_1
XFILLER_141_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8956_ _8955_/S _6322_/Y _8977_/S VGND VGND VPWR VPWR _8956_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7907_ _7864_/X _8230_/A _7887_/Y _7893_/X _7906_/X VGND VGND VPWR VPWR _7907_/X
+ sky130_fd_sc_hd__o2111a_2
XFILLER_169_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8887_ _8886_/X _9144_/Q _9054_/Q VGND VGND VPWR VPWR _8887_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7838_ _8379_/D _7838_/B _8394_/D _7879_/A VGND VGND VPWR VPWR _8298_/A sky130_fd_sc_hd__or4_1
XFILLER_51_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7769_ _8528_/A VGND VGND VPWR VPWR _8193_/A sky130_fd_sc_hd__clkinv_4
X_9508_ _9508_/CLK _9508_/D _9528_/SET_B VGND VGND VPWR VPWR _9508_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_109_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9439_ _9440_/CLK _9439_/D _9685_/SET_B VGND VGND VPWR VPWR _9439_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_137_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5120_ _9632_/Q _5112_/A _5967_/B1 _5112_/Y VGND VGND VPWR VPWR _9632_/D sky130_fd_sc_hd__a22o_1
XFILLER_151_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5051_ _9671_/Q _5047_/A _8925_/A1 _5047_/Y VGND VGND VPWR VPWR _9671_/D sky130_fd_sc_hd__a22o_1
XFILLER_111_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8810_ _8810_/A _8813_/B VGND VGND VPWR VPWR _9063_/D sky130_fd_sc_hd__nor2_1
X_9790_ _9790_/CLK _9790_/D _9757_/SET_B VGND VGND VPWR VPWR _9790_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_53_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8741_ _8732_/Y _8733_/Y _8735_/X _8740_/X VGND VGND VPWR VPWR _8741_/X sky130_fd_sc_hd__a31o_1
XFILLER_92_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5953_ _9112_/Q _5951_/A _8845_/X _5951_/Y VGND VGND VPWR VPWR _9112_/D sky130_fd_sc_hd__a22o_1
XFILLER_80_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8672_ _8703_/B _8672_/B _8672_/C VGND VGND VPWR VPWR _8673_/C sky130_fd_sc_hd__or3_1
X_4904_ _6158_/A _4927_/A _4901_/Y _4902_/Y _5412_/B VGND VGND VPWR VPWR _4904_/X
+ sky130_fd_sc_hd__o32a_1
X_5884_ _5849_/X _8895_/X _8924_/X _9149_/Q VGND VGND VPWR VPWR _9149_/D sky130_fd_sc_hd__o22a_1
XFILLER_33_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4835_ _9081_/Q VGND VGND VPWR VPWR _4835_/Y sky130_fd_sc_hd__clkinv_4
X_7623_ _4882_/Y _7475_/X _4706_/Y _7477_/X VGND VGND VPWR VPWR _7623_/X sky130_fd_sc_hd__o22a_1
X_7554_ _7554_/A _7554_/B _7554_/C _7554_/D VGND VGND VPWR VPWR _7554_/Y sky130_fd_sc_hd__nand4_4
X_4766_ _6111_/B _4843_/B VGND VGND VPWR VPWR _5960_/B sky130_fd_sc_hd__or2_4
X_6505_ _6505_/A VGND VGND VPWR VPWR _6505_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7485_ _6910_/Y _7419_/X _6844_/Y _7421_/X VGND VGND VPWR VPWR _7485_/X sky130_fd_sc_hd__o22a_1
X_4697_ _4787_/A _4903_/B VGND VGND VPWR VPWR _4698_/A sky130_fd_sc_hd__or2_1
XFILLER_161_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6436_ _9368_/Q VGND VGND VPWR VPWR _6436_/Y sky130_fd_sc_hd__inv_2
X_9224_ _9695_/CLK _9224_/D _9779_/SET_B VGND VGND VPWR VPWR _9224_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6367_ _9208_/Q VGND VGND VPWR VPWR _6367_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_136_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9155_ _9695_/CLK _9155_/D _9646_/SET_B VGND VGND VPWR VPWR _9155_/Q sky130_fd_sc_hd__dfrtp_1
X_8106_ _8200_/C VGND VGND VPWR VPWR _8218_/C sky130_fd_sc_hd__inv_2
X_5318_ _5318_/A VGND VGND VPWR VPWR _5319_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6298_ _9195_/Q VGND VGND VPWR VPWR _6298_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9086_ _9089_/CLK _9086_/D _6004_/X VGND VGND VPWR VPWR _9086_/Q sky130_fd_sc_hd__dfrtp_2
X_8037_ _8544_/A _7987_/Y _8036_/Y VGND VGND VPWR VPWR _8039_/A sky130_fd_sc_hd__a21oi_1
X_5249_ _9547_/Q _5242_/A _5966_/B1 _5242_/Y VGND VGND VPWR VPWR _9547_/D sky130_fd_sc_hd__a22o_1
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8939_ _9710_/Q _9759_/Q _9587_/Q VGND VGND VPWR VPWR _8939_/X sky130_fd_sc_hd__mux2_8
XFILLER_169_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4620_ _9721_/Q _4615_/A _5967_/B1 _4615_/Y VGND VGND VPWR VPWR _9721_/D sky130_fd_sc_hd__a22o_1
XFILLER_187_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4551_ _9065_/Q _4551_/B VGND VGND VPWR VPWR _4551_/X sky130_fd_sc_hd__or2_1
X_4482_ _8955_/A1 _9788_/Q _6018_/S VGND VGND VPWR VPWR _4483_/A sky130_fd_sc_hd__mux2_1
X_7270_ _6140_/Y _7048_/B _6120_/Y _7077_/A _7269_/X VGND VGND VPWR VPWR _7277_/A
+ sky130_fd_sc_hd__o221a_1
X_6221_ _6221_/A VGND VGND VPWR VPWR _6221_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_131_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6152_ _9378_/Q VGND VGND VPWR VPWR _6152_/Y sky130_fd_sc_hd__inv_2
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5103_ _9645_/Q _5102_/A _5963_/B1 _5102_/Y VGND VGND VPWR VPWR _9645_/D sky130_fd_sc_hd__a22o_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6083_ _9553_/Q VGND VGND VPWR VPWR _6083_/Y sky130_fd_sc_hd__clkinv_4
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ _9052_/Q VGND VGND VPWR VPWR _5034_/Y sky130_fd_sc_hd__inv_2
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater366 _8840_/X VGND VGND VPWR VPWR _5966_/B1 sky130_fd_sc_hd__buf_12
XFILLER_72_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater377 _9757_/SET_B VGND VGND VPWR VPWR _9633_/SET_B sky130_fd_sc_hd__buf_12
X_9773_ _9775_/CLK _9773_/D _7011_/B VGND VGND VPWR VPWR _9773_/Q sky130_fd_sc_hd__dfrtp_1
X_6985_ _9710_/Q _9569_/Q _8977_/S VGND VGND VPWR VPWR _8809_/A sky130_fd_sc_hd__o21ai_4
X_5936_ _5936_/A _5936_/B _5936_/C _5936_/D VGND VGND VPWR VPWR _5939_/B sky130_fd_sc_hd__or4_2
X_8724_ _8729_/A _8731_/C _8723_/Y VGND VGND VPWR VPWR _8724_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_80_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8655_ _8655_/A VGND VGND VPWR VPWR _8655_/Y sky130_fd_sc_hd__inv_2
X_5867_ _9163_/Q _5866_/A _8843_/X _5866_/Y VGND VGND VPWR VPWR _9163_/D sky130_fd_sc_hd__a22o_1
X_7606_ _6128_/Y _7471_/X _7282_/A _7473_/X _7605_/X VGND VGND VPWR VPWR _7607_/D
+ sky130_fd_sc_hd__o221a_1
X_8586_ _8586_/A _8646_/B _8678_/B _8721_/B VGND VGND VPWR VPWR _8588_/B sky130_fd_sc_hd__or4_1
XFILLER_166_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5798_ _5798_/A VGND VGND VPWR VPWR _5799_/A sky130_fd_sc_hd__clkbuf_4
X_4818_ _9719_/Q VGND VGND VPWR VPWR _4818_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_21_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4749_ _9302_/Q VGND VGND VPWR VPWR _4749_/Y sky130_fd_sc_hd__clkinv_2
X_7537_ _6396_/Y _7408_/X _6334_/Y _7410_/X VGND VGND VPWR VPWR _7537_/X sky130_fd_sc_hd__o22a_1
X_7468_ _4734_/Y _7465_/X _4855_/Y _7467_/X VGND VGND VPWR VPWR _7468_/X sky130_fd_sc_hd__o22a_1
XFILLER_110_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9207_ _9788_/CLK _9207_/D _9647_/SET_B VGND VGND VPWR VPWR _9207_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_134_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6419_ _6417_/Y _5412_/B _6418_/Y _5024_/B VGND VGND VPWR VPWR _6419_/X sky130_fd_sc_hd__o22a_2
XFILLER_134_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7399_ _7476_/A _9251_/Q _7456_/A _7474_/D VGND VGND VPWR VPWR _7400_/A sky130_fd_sc_hd__or4_1
XFILLER_163_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9138_ _9203_/CLK _9138_/D _9633_/SET_B VGND VGND VPWR VPWR _9138_/Q sky130_fd_sc_hd__dfrtp_1
Xinput136 wb_adr_i[13] VGND VGND VPWR VPWR _7771_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_163_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput125 trap VGND VGND VPWR VPWR _4901_/A sky130_fd_sc_hd__buf_6
Xinput114 sram_ro_data[29] VGND VGND VPWR VPWR _6249_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9069_ _9790_/CLK _9069_/D _9757_/SET_B VGND VGND VPWR VPWR _9069_/Q sky130_fd_sc_hd__dfrtp_4
Xinput103 sram_ro_data[19] VGND VGND VPWR VPWR _6558_/A sky130_fd_sc_hd__clkbuf_1
Xinput169 wb_dat_i[13] VGND VGND VPWR VPWR _7747_/B2 sky130_fd_sc_hd__clkbuf_1
Xinput147 wb_adr_i[23] VGND VGND VPWR VPWR _7781_/A sky130_fd_sc_hd__clkbuf_1
Xinput158 wb_adr_i[4] VGND VGND VPWR VPWR _7894_/B sky130_fd_sc_hd__buf_4
XFILLER_48_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_2_csclk clkbuf_leaf_2_csclk/A VGND VGND VPWR VPWR _9514_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6770_ _6768_/Y _4564_/B _6769_/Y _6086_/X VGND VGND VPWR VPWR _6770_/X sky130_fd_sc_hd__o22a_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5721_ _9247_/Q VGND VGND VPWR VPWR _7056_/B sky130_fd_sc_hd__inv_2
XFILLER_176_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8440_ _7864_/X _8230_/A _8544_/A _8115_/Y VGND VGND VPWR VPWR _8665_/A sky130_fd_sc_hd__a2bb2o_1
X_5652_ _5649_/B _5647_/X _5649_/A VGND VGND VPWR VPWR _5652_/Y sky130_fd_sc_hd__o21ai_1
X_5583_ _6052_/A _5583_/B VGND VGND VPWR VPWR _5584_/A sky130_fd_sc_hd__or2_1
XFILLER_129_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8371_ _8708_/D _8506_/B VGND VGND VPWR VPWR _8715_/C sky130_fd_sc_hd__or2_1
X_4603_ _4603_/A VGND VGND VPWR VPWR _4604_/A sky130_fd_sc_hd__buf_2
X_7322_ _6938_/Y _7112_/X _6896_/Y _7077_/B VGND VGND VPWR VPWR _7322_/X sky130_fd_sc_hd__o22a_1
X_4534_ _9762_/Q _4526_/A _5967_/B1 _4526_/Y VGND VGND VPWR VPWR _9762_/D sky130_fd_sc_hd__a22o_1
XFILLER_144_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7253_ _6182_/Y _7068_/A _6199_/Y _7105_/X VGND VGND VPWR VPWR _7253_/X sky130_fd_sc_hd__o22a_1
X_4465_ _4465_/A VGND VGND VPWR VPWR _4466_/A sky130_fd_sc_hd__buf_2
XFILLER_131_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7184_ _8775_/A _7095_/X _8755_/A _7068_/D _7183_/X VGND VGND VPWR VPWR _7189_/B
+ sky130_fd_sc_hd__o221a_1
X_6204_ _6199_/Y _5240_/B _6200_/Y _5393_/B _6203_/X VGND VGND VPWR VPWR _6211_/C
+ sky130_fd_sc_hd__o221a_1
X_6135_ _6135_/A VGND VGND VPWR VPWR _8926_/S sky130_fd_sc_hd__clkinv_8
XFILLER_112_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6066_ _9276_/Q VGND VGND VPWR VPWR _6066_/Y sky130_fd_sc_hd__clkinv_2
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5017_ _9694_/Q _5015_/A _8845_/X _5015_/Y VGND VGND VPWR VPWR _9694_/D sky130_fd_sc_hd__a22o_1
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9756_ _9757_/CLK _9756_/D _9757_/SET_B VGND VGND VPWR VPWR _9756_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_26_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8707_ _8707_/A _8707_/B _8707_/C VGND VGND VPWR VPWR _8733_/A sky130_fd_sc_hd__or3_2
X_6968_ _6475_/Y _6964_/A _9024_/Q _6964_/Y VGND VGND VPWR VPWR _9024_/D sky130_fd_sc_hd__o22a_2
X_9687_ _9687_/CLK _9687_/D _9685_/SET_B VGND VGND VPWR VPWR _9687_/Q sky130_fd_sc_hd__dfrtp_1
X_6899_ _6897_/Y _5810_/B _6898_/Y _5556_/B VGND VGND VPWR VPWR _6899_/X sky130_fd_sc_hd__o22a_1
X_5919_ _9124_/Q _5918_/A _5963_/B1 _5918_/Y VGND VGND VPWR VPWR _9124_/D sky130_fd_sc_hd__a22o_1
X_8638_ _8721_/B VGND VGND VPWR VPWR _8638_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8569_ _8640_/A _8568_/X _8223_/A _8352_/C VGND VGND VPWR VPWR _8719_/A sky130_fd_sc_hd__o211ai_4
XFILLER_181_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7940_ _8202_/A _8341_/A _7939_/X VGND VGND VPWR VPWR _7941_/B sky130_fd_sc_hd__o21ai_1
XFILLER_103_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7871_ _8515_/B _8246_/B VGND VGND VPWR VPWR _8734_/A sky130_fd_sc_hd__nor2_2
X_9610_ _9613_/CLK _9610_/D _9646_/SET_B VGND VGND VPWR VPWR _9610_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6822_ _6817_/Y _4832_/X _6818_/Y _5393_/B _6821_/X VGND VGND VPWR VPWR _6829_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_35_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6753_ _9392_/Q VGND VGND VPWR VPWR _6753_/Y sky130_fd_sc_hd__inv_2
X_9541_ _9545_/CLK _9541_/D _4628_/A VGND VGND VPWR VPWR _9541_/Q sky130_fd_sc_hd__dfrtp_1
X_9472_ _9684_/CLK _9472_/D _9685_/SET_B VGND VGND VPWR VPWR _9472_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_148_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6684_ _6679_/Y _4861_/X _6680_/Y _6322_/A _6683_/X VGND VGND VPWR VPWR _6690_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_31_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5704_ _7462_/A VGND VGND VPWR VPWR _5704_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5635_ _9285_/Q _5634_/A _8843_/X _5634_/Y VGND VGND VPWR VPWR _9285_/D sky130_fd_sc_hd__a22o_1
X_8423_ _8708_/A _8708_/B _8422_/X VGND VGND VPWR VPWR _8423_/X sky130_fd_sc_hd__or3b_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8354_ _8354_/A _8595_/B VGND VGND VPWR VPWR _8571_/C sky130_fd_sc_hd__or2_1
X_5566_ _5566_/A VGND VGND VPWR VPWR _5566_/Y sky130_fd_sc_hd__inv_2
X_8285_ _8476_/B _8285_/B VGND VGND VPWR VPWR _8286_/C sky130_fd_sc_hd__or2_1
XFILLER_132_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7305_ _4858_/Y _5728_/X _4692_/A _7040_/A _7304_/X VGND VGND VPWR VPWR _7308_/C
+ sky130_fd_sc_hd__o221a_2
XFILLER_104_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4517_ _4517_/A VGND VGND VPWR VPWR _4517_/Y sky130_fd_sc_hd__inv_2
X_5497_ _5497_/A VGND VGND VPWR VPWR _5498_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_132_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7236_ _6275_/Y _7118_/X _6321_/Y _7048_/C VGND VGND VPWR VPWR _7236_/X sky130_fd_sc_hd__o22a_1
X_4448_ _9584_/Q input77/X _8801_/B VGND VGND VPWR VPWR _8983_/A sky130_fd_sc_hd__mux2_1
X_7167_ _7167_/A _7167_/B _7167_/C _7167_/D VGND VGND VPWR VPWR _7177_/B sky130_fd_sc_hd__and4_1
XFILLER_86_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6118_ _6113_/Y _5382_/B _6114_/Y _5355_/B _6117_/X VGND VGND VPWR VPWR _6119_/D
+ sky130_fd_sc_hd__o221a_1
X_7098_ _9246_/Q _9245_/Q _7098_/C _7127_/C VGND VGND VPWR VPWR _7099_/A sky130_fd_sc_hd__or4_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6049_ _6049_/A VGND VGND VPWR VPWR _6049_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9739_ _9774_/CLK _9739_/D _9757_/SET_B VGND VGND VPWR VPWR _9739_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_41_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_20_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR _9596_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_110_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_35_csclk clkbuf_opt_4_0_csclk/X VGND VGND VPWR VPWR _9790_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_60_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5420_ _5545_/A _5420_/B VGND VGND VPWR VPWR _5421_/A sky130_fd_sc_hd__or2_1
XFILLER_145_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput226 _8784_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[26] sky130_fd_sc_hd__buf_2
X_5351_ _9479_/Q _5346_/A _8842_/X _5346_/Y VGND VGND VPWR VPWR _9479_/D sky130_fd_sc_hd__a22o_1
XFILLER_173_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput215 _8764_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[16] sky130_fd_sc_hd__buf_2
XFILLER_145_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput204 _8806_/X VGND VGND VPWR VPWR debug_in sky130_fd_sc_hd__buf_2
Xoutput237 _8834_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[36] sky130_fd_sc_hd__buf_2
Xoutput248 _8828_/X VGND VGND VPWR VPWR mgmt_gpio_out[35] sky130_fd_sc_hd__buf_2
X_5282_ _9526_/Q _5280_/A _8845_/X _5280_/Y VGND VGND VPWR VPWR _9526_/D sky130_fd_sc_hd__a22o_1
XFILLER_160_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8070_ _8515_/A _8305_/A _8069_/Y VGND VGND VPWR VPWR _8074_/A sky130_fd_sc_hd__o21bai_1
Xoutput259 _7017_/Y VGND VGND VPWR VPWR pad_flash_io1_ieb sky130_fd_sc_hd__buf_2
X_7021_ _7021_/A VGND VGND VPWR VPWR _7021_/X sky130_fd_sc_hd__buf_4
XFILLER_141_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8972_ _8655_/Y _8604_/X _8975_/S VGND VGND VPWR VPWR _8972_/X sky130_fd_sc_hd__mux2_2
XFILLER_83_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7923_ _8667_/A _7923_/B VGND VGND VPWR VPWR _7924_/B sky130_fd_sc_hd__or2_1
XFILLER_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7854_ _8515_/B _8270_/B VGND VGND VPWR VPWR _8615_/A sky130_fd_sc_hd__nor2_1
XFILLER_51_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7785_ _8583_/A _8189_/A _7791_/B VGND VGND VPWR VPWR _7787_/B sky130_fd_sc_hd__or3_1
X_6805_ _9555_/Q VGND VGND VPWR VPWR _6805_/Y sky130_fd_sc_hd__clkinv_2
X_6736_ _9478_/Q VGND VGND VPWR VPWR _6736_/Y sky130_fd_sc_hd__clkinv_4
X_9524_ _9527_/CLK _9524_/D _9528_/SET_B VGND VGND VPWR VPWR _9524_/Q sky130_fd_sc_hd__dfrtp_1
X_4997_ _4997_/A VGND VGND VPWR VPWR _9699_/D sky130_fd_sc_hd__clkbuf_1
X_9455_ _9483_/CLK _9455_/D _9528_/SET_B VGND VGND VPWR VPWR _9455_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_176_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6667_ _9669_/Q VGND VGND VPWR VPWR _6667_/Y sky130_fd_sc_hd__inv_2
X_5618_ _9296_/Q _5612_/A _8955_/A1 _5612_/Y VGND VGND VPWR VPWR _9296_/D sky130_fd_sc_hd__a22o_1
X_8406_ _8130_/B _8401_/B _8402_/X _8405_/Y VGND VGND VPWR VPWR _8406_/X sky130_fd_sc_hd__o211a_1
X_6598_ _9549_/Q VGND VGND VPWR VPWR _8785_/A sky130_fd_sc_hd__inv_8
X_9386_ _9777_/CLK _9386_/D _7011_/B VGND VGND VPWR VPWR _9386_/Q sky130_fd_sc_hd__dfrtp_1
X_5549_ _9344_/Q _5547_/A _8845_/X _5547_/Y VGND VGND VPWR VPWR _9344_/D sky130_fd_sc_hd__a22o_1
X_8337_ _8636_/A _8650_/B _8337_/C VGND VGND VPWR VPWR _8338_/A sky130_fd_sc_hd__or3_1
XFILLER_124_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8268_ _8660_/A _8270_/B VGND VGND VPWR VPWR _8579_/B sky130_fd_sc_hd__nor2_1
X_8199_ _8213_/B VGND VGND VPWR VPWR _8340_/B sky130_fd_sc_hd__clkinvlp_2
X_7219_ _6328_/Y _7124_/X _6410_/Y _7068_/B _7218_/X VGND VGND VPWR VPWR _7220_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_171_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_6_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A VGND VGND VPWR VPWR _4450_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_89_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4920_ _9359_/Q VGND VGND VPWR VPWR _4920_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_18_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4851_ _4911_/A _4898_/A VGND VGND VPWR VPWR _5355_/B sky130_fd_sc_hd__or2_4
X_7570_ _6302_/Y _7471_/X _7238_/A _7473_/X _7569_/X VGND VGND VPWR VPWR _7571_/D
+ sky130_fd_sc_hd__o221a_1
X_4782_ _4787_/A _4898_/A VGND VGND VPWR VPWR _4783_/A sky130_fd_sc_hd__or2_1
XFILLER_60_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6521_ _6521_/A VGND VGND VPWR VPWR _6521_/Y sky130_fd_sc_hd__inv_4
XFILLER_158_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9240_ _9789_/CLK _9240_/D _9647_/SET_B VGND VGND VPWR VPWR _9240_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6452_ _9730_/Q VGND VGND VPWR VPWR _6452_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9171_ _9280_/CLK _9171_/D _9757_/SET_B VGND VGND VPWR VPWR _9171_/Q sky130_fd_sc_hd__dfrtp_1
X_5403_ _9442_/Q _5395_/A _8916_/A1 _5395_/Y VGND VGND VPWR VPWR _9442_/D sky130_fd_sc_hd__a22o_1
X_8122_ _7886_/B _8566_/A _8546_/A _8121_/Y VGND VGND VPWR VPWR _8122_/X sky130_fd_sc_hd__o31a_1
X_6383_ _6367_/Y _5797_/B _6370_/X _6376_/X _6382_/X VGND VGND VPWR VPWR _6475_/C
+ sky130_fd_sc_hd__o2111a_1
X_5334_ _9490_/Q _5330_/A _5966_/B1 _5330_/Y VGND VGND VPWR VPWR _9490_/D sky130_fd_sc_hd__a22o_1
X_8053_ _8053_/A _8392_/A VGND VGND VPWR VPWR _8055_/A sky130_fd_sc_hd__nand2_1
X_5265_ _9537_/Q _5261_/A _5966_/B1 _5261_/Y VGND VGND VPWR VPWR _9537_/D sky130_fd_sc_hd__a22o_1
XFILLER_87_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5196_ _9583_/Q _5193_/Y _8915_/X _5193_/A VGND VGND VPWR VPWR _9583_/D sky130_fd_sc_hd__o22a_1
X_7004_ _4964_/B _7008_/A _7008_/B _6022_/B _7003_/X VGND VGND VPWR VPWR _7005_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_28_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8955_ _9620_/Q _8955_/A1 _8955_/S VGND VGND VPWR VPWR _8955_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7906_ _7864_/X _7885_/B _7896_/X _7902_/X _7905_/X VGND VGND VPWR VPWR _7906_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_83_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8886_ _7287_/Y _9639_/Q _8959_/S VGND VGND VPWR VPWR _8886_/X sky130_fd_sc_hd__mux2_1
X_7837_ _7837_/A _7837_/B _7837_/C VGND VGND VPWR VPWR _7879_/A sky130_fd_sc_hd__or3_4
XFILLER_70_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7768_ _7768_/A _7768_/B _7768_/C _7768_/D VGND VGND VPWR VPWR _7966_/A sky130_fd_sc_hd__nand4_1
XFILLER_51_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9507_ _9509_/CLK _9507_/D _9528_/SET_B VGND VGND VPWR VPWR _9507_/Q sky130_fd_sc_hd__dfrtp_1
X_7699_ _7699_/A VGND VGND VPWR VPWR _7700_/A sky130_fd_sc_hd__clkbuf_1
X_6719_ _9408_/Q VGND VGND VPWR VPWR _6719_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_50_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9438_ _9514_/CLK _9438_/D _9685_/SET_B VGND VGND VPWR VPWR _9438_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9369_ _9371_/CLK _9369_/D _9295_/SET_B VGND VGND VPWR VPWR _9369_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5050_ _9672_/Q _5047_/A _8844_/X _5047_/Y VGND VGND VPWR VPWR _9672_/D sky130_fd_sc_hd__a22o_1
XFILLER_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8740_ _8712_/B _8737_/Y _8689_/A _8738_/Y _8739_/Y VGND VGND VPWR VPWR _8740_/X
+ sky130_fd_sc_hd__o311a_1
X_5952_ _9113_/Q _5951_/A _8846_/X _5951_/Y VGND VGND VPWR VPWR _9113_/D sky130_fd_sc_hd__a22o_1
XFILLER_1_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4903_ _4911_/A _4903_/B VGND VGND VPWR VPWR _5412_/B sky130_fd_sc_hd__or2_4
X_8671_ _8735_/D _8699_/D _8671_/C _8703_/A VGND VGND VPWR VPWR _8671_/Y sky130_fd_sc_hd__nor4_2
X_5883_ _5849_/X _8897_/X _8924_/X _9150_/Q VGND VGND VPWR VPWR _9150_/D sky130_fd_sc_hd__o22a_1
X_7622_ _4694_/Y _7461_/X _4883_/Y _7463_/X _7621_/X VGND VGND VPWR VPWR _7625_/C
+ sky130_fd_sc_hd__o221a_1
X_4834_ _4911_/A _4876_/B VGND VGND VPWR VPWR _5431_/B sky130_fd_sc_hd__or2_4
XFILLER_60_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7553_ _7553_/A _7553_/B _7553_/C _7553_/D VGND VGND VPWR VPWR _7554_/D sky130_fd_sc_hd__and4_1
X_4765_ _9101_/Q VGND VGND VPWR VPWR _4765_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_193_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6504_ _9188_/Q VGND VGND VPWR VPWR _6504_/Y sky130_fd_sc_hd__clkinv_4
X_4696_ _8805_/A VGND VGND VPWR VPWR _4696_/Y sky130_fd_sc_hd__inv_2
X_7484_ _6859_/Y _7400_/X _6891_/Y _7405_/X _7483_/X VGND VGND VPWR VPWR _7500_/A
+ sky130_fd_sc_hd__o221a_1
X_9223_ _9695_/CLK _9223_/D _9646_/SET_B VGND VGND VPWR VPWR _9223_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_174_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6435_ _9636_/Q VGND VGND VPWR VPWR _6435_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9154_ _9695_/CLK _9154_/D _9779_/SET_B VGND VGND VPWR VPWR _9154_/Q sky130_fd_sc_hd__dfrtp_1
X_6366_ _6353_/Y _5818_/B _6355_/X _6359_/X _6365_/X VGND VGND VPWR VPWR _6475_/B
+ sky130_fd_sc_hd__o2111a_2
X_8105_ _7756_/B _8103_/Y _7837_/B _8103_/A VGND VGND VPWR VPWR _8200_/C sky130_fd_sc_hd__o22a_1
X_5317_ _5545_/A _5317_/B VGND VGND VPWR VPWR _5318_/A sky130_fd_sc_hd__or2_1
XFILLER_0_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9085_ _9089_/CLK _9085_/D _6007_/X VGND VGND VPWR VPWR _9085_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_102_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8036_ _8389_/A _8551_/A _8035_/X VGND VGND VPWR VPWR _8036_/Y sky130_fd_sc_hd__o21ai_1
X_6297_ _9693_/Q VGND VGND VPWR VPWR _6297_/Y sky130_fd_sc_hd__clkinv_2
X_5248_ _9548_/Q _5242_/A _5965_/B1 _5242_/Y VGND VGND VPWR VPWR _9548_/D sky130_fd_sc_hd__a22o_1
XFILLER_29_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5179_ _5179_/A VGND VGND VPWR VPWR _5180_/A sky130_fd_sc_hd__buf_2
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8938_ _8937_/X _9680_/Q _9587_/Q VGND VGND VPWR VPWR _8938_/X sky130_fd_sc_hd__mux2_2
XFILLER_71_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8869_ _8868_/X _9173_/Q _9054_/Q VGND VGND VPWR VPWR _8869_/X sky130_fd_sc_hd__mux2_1
XPHY_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4550_ _4551_/B VGND VGND VPWR VPWR _5062_/D sky130_fd_sc_hd__inv_6
XFILLER_128_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4481_ _5259_/A _4481_/B VGND VGND VPWR VPWR _6018_/S sky130_fd_sc_hd__or2_2
XFILLER_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6220_ _9754_/Q VGND VGND VPWR VPWR _6220_/Y sky130_fd_sc_hd__inv_2
X_6151_ _9344_/Q VGND VGND VPWR VPWR _6151_/Y sky130_fd_sc_hd__clkinv_2
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ _5102_/A VGND VGND VPWR VPWR _5102_/Y sky130_fd_sc_hd__inv_2
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6082_ _6078_/Y _5344_/B _6079_/Y _5278_/B _6081_/X VGND VGND VPWR VPWR _6096_/B
+ sky130_fd_sc_hd__o221a_2
XFILLER_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5033_ _5033_/A VGND VGND VPWR VPWR _5033_/X sky130_fd_sc_hd__clkbuf_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater367 _8840_/X VGND VGND VPWR VPWR _8930_/A1 sky130_fd_sc_hd__buf_12
XFILLER_122_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater378 _7011_/B VGND VGND VPWR VPWR _9757_/SET_B sky130_fd_sc_hd__buf_12
X_6984_ _4936_/Y _6976_/A _9012_/Q _6976_/Y VGND VGND VPWR VPWR _9012_/D sky130_fd_sc_hd__o22a_1
X_9772_ _9790_/CLK _9772_/D _9757_/SET_B VGND VGND VPWR VPWR _9772_/Q sky130_fd_sc_hd__dfrtp_4
X_5935_ _7837_/C _5935_/B _5935_/C _5934_/X VGND VGND VPWR VPWR _5936_/D sky130_fd_sc_hd__or4b_1
X_8723_ _8723_/A _8723_/B _8723_/C VGND VGND VPWR VPWR _8723_/Y sky130_fd_sc_hd__nor3_4
X_5866_ _5866_/A VGND VGND VPWR VPWR _5866_/Y sky130_fd_sc_hd__inv_2
X_8654_ _8705_/A _8707_/B _8620_/Y _8637_/X _8653_/X VGND VGND VPWR VPWR _8655_/A
+ sky130_fd_sc_hd__o311a_1
XFILLER_33_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7605_ _6104_/Y _7475_/X _6066_/Y _7477_/X VGND VGND VPWR VPWR _7605_/X sky130_fd_sc_hd__o22a_1
X_4817_ _4911_/A _4927_/A VGND VGND VPWR VPWR _5393_/B sky130_fd_sc_hd__or2_4
XFILLER_166_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8585_ _8585_/A _8585_/B VGND VGND VPWR VPWR _8721_/B sky130_fd_sc_hd__or2_1
X_5797_ _6052_/A _5797_/B VGND VGND VPWR VPWR _5798_/A sky130_fd_sc_hd__or2_1
XFILLER_21_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4748_ _4726_/Y _5660_/B _4731_/X _4736_/X _4747_/X VGND VGND VPWR VPWR _4791_/C
+ sky130_fd_sc_hd__o2111a_1
X_7536_ _7536_/A _7536_/B _7536_/C _7536_/D VGND VGND VPWR VPWR _7536_/Y sky130_fd_sc_hd__nand4_4
X_4679_ _4787_/A _4925_/A VGND VGND VPWR VPWR _5178_/B sky130_fd_sc_hd__or2_4
X_7467_ _7467_/A VGND VGND VPWR VPWR _7467_/X sky130_fd_sc_hd__buf_8
X_6418_ _9687_/Q VGND VGND VPWR VPWR _6418_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_162_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9206_ _9652_/CLK _9206_/D _9647_/SET_B VGND VGND VPWR VPWR _9206_/Q sky130_fd_sc_hd__dfrtp_1
X_9137_ _9354_/CLK _9137_/D _9685_/SET_B VGND VGND VPWR VPWR _9137_/Q sky130_fd_sc_hd__dfrtp_1
X_7398_ _7456_/A _7462_/A _9255_/Q VGND VGND VPWR VPWR _8978_/S sky130_fd_sc_hd__nor3_4
X_6349_ _9524_/Q VGND VGND VPWR VPWR _6349_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9068_ _4450_/A1 _9068_/D _6146_/A VGND VGND VPWR VPWR _9068_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_163_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput126 uart_enabled VGND VGND VPWR VPWR _8801_/B sky130_fd_sc_hd__buf_4
XFILLER_0_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput104 sram_ro_data[1] VGND VGND VPWR VPWR _6820_/A sky130_fd_sc_hd__clkbuf_1
Xinput115 sram_ro_data[2] VGND VGND VPWR VPWR _6679_/A sky130_fd_sc_hd__clkbuf_1
Xinput148 wb_adr_i[24] VGND VGND VPWR VPWR _5925_/C sky130_fd_sc_hd__clkbuf_1
Xinput137 wb_adr_i[14] VGND VGND VPWR VPWR _7770_/B sky130_fd_sc_hd__clkbuf_1
Xinput159 wb_adr_i[5] VGND VGND VPWR VPWR _8525_/A sky130_fd_sc_hd__buf_6
X_8019_ _8612_/A _8016_/X _8019_/C _8441_/B VGND VGND VPWR VPWR _8019_/X sky130_fd_sc_hd__and4bb_1
XFILLER_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5720_ _9248_/Q VGND VGND VPWR VPWR _7037_/A sky130_fd_sc_hd__inv_2
XFILLER_176_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5651_ _5658_/A _5651_/B VGND VGND VPWR VPWR _5651_/X sky130_fd_sc_hd__or2_1
XFILLER_175_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5582_ _9320_/Q _5574_/A _8916_/A1 _5574_/Y VGND VGND VPWR VPWR _9320_/D sky130_fd_sc_hd__a22o_1
X_8370_ _8370_/A _8599_/B VGND VGND VPWR VPWR _8579_/C sky130_fd_sc_hd__or2_1
X_4602_ _5960_/A _4602_/B VGND VGND VPWR VPWR _4603_/A sky130_fd_sc_hd__or2_1
XFILLER_129_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7321_ _7321_/A _7321_/B _7321_/C _7321_/D VGND VGND VPWR VPWR _7331_/B sky130_fd_sc_hd__and4_1
X_4533_ _9763_/Q _4526_/A _5966_/B1 _4526_/Y VGND VGND VPWR VPWR _9763_/D sky130_fd_sc_hd__a22o_1
XFILLER_7_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7252_ _6170_/Y _7059_/B _6201_/Y _7068_/C _7251_/X VGND VGND VPWR VPWR _7255_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6203_ _6201_/Y _6081_/B _6202_/Y _4590_/B VGND VGND VPWR VPWR _6203_/X sky130_fd_sc_hd__o22a_1
X_4464_ _5960_/A _6251_/A VGND VGND VPWR VPWR _4465_/A sky130_fd_sc_hd__or2_1
X_7183_ _8777_/A _7097_/X _8787_/A _7099_/X VGND VGND VPWR VPWR _7183_/X sky130_fd_sc_hd__o22a_1
X_6134_ _6134_/A VGND VGND VPWR VPWR _8930_/S sky130_fd_sc_hd__clkinv_8
XFILLER_112_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6065_ _9184_/Q VGND VGND VPWR VPWR _6065_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_133_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5016_ _9695_/Q _5015_/A _8846_/X _5015_/Y VGND VGND VPWR VPWR _9695_/D sky130_fd_sc_hd__a22o_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6967_ _6326_/Y _6964_/A _9025_/Q _6964_/Y VGND VGND VPWR VPWR _9025_/D sky130_fd_sc_hd__o22a_1
X_9755_ _9755_/CLK _9755_/D _9757_/SET_B VGND VGND VPWR VPWR _9755_/Q sky130_fd_sc_hd__dfstp_1
X_8706_ _8706_/A _8706_/B _8706_/C _8706_/D VGND VGND VPWR VPWR _8707_/C sky130_fd_sc_hd__or4_1
XFILLER_81_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5918_ _5918_/A VGND VGND VPWR VPWR _5918_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9686_ _9687_/CLK _9686_/D _9685_/SET_B VGND VGND VPWR VPWR _9686_/Q sky130_fd_sc_hd__dfrtp_1
X_6898_ _9334_/Q VGND VGND VPWR VPWR _6898_/Y sky130_fd_sc_hd__inv_2
XFILLER_139_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8637_ _8621_/Y _8633_/Y _8635_/Y _8714_/C VGND VGND VPWR VPWR _8637_/X sky130_fd_sc_hd__a31o_1
X_5849_ _5849_/A VGND VGND VPWR VPWR _5849_/X sky130_fd_sc_hd__buf_6
XFILLER_166_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8568_ _8213_/A _8640_/C _8215_/X VGND VGND VPWR VPWR _8568_/X sky130_fd_sc_hd__o21a_1
XFILLER_107_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7519_ _8767_/A _7400_/X _8757_/A _7405_/X VGND VGND VPWR VPWR _7519_/X sky130_fd_sc_hd__o22a_1
XFILLER_5_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8499_ _8571_/B _8499_/B VGND VGND VPWR VPWR _8659_/A sky130_fd_sc_hd__or2_1
XFILLER_135_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7870_ _7870_/A VGND VGND VPWR VPWR _8246_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_23_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6821_ _6819_/Y _5431_/B _6820_/Y _4861_/X VGND VGND VPWR VPWR _6821_/X sky130_fd_sc_hd__o22a_1
XFILLER_90_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9540_ _9768_/CLK _9540_/D _4628_/A VGND VGND VPWR VPWR _9540_/Q sky130_fd_sc_hd__dfrtp_1
X_6752_ _6748_/Y _5621_/B _6749_/Y _6052_/C _6751_/X VGND VGND VPWR VPWR _6759_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_16_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9471_ _9687_/CLK _9471_/D _9685_/SET_B VGND VGND VPWR VPWR _9471_/Q sky130_fd_sc_hd__dfrtp_4
X_6683_ _6681_/Y _5013_/B _6682_/Y _5829_/B VGND VGND VPWR VPWR _6683_/X sky130_fd_sc_hd__o22a_1
X_5703_ _9253_/Q VGND VGND VPWR VPWR _7406_/B sky130_fd_sc_hd__inv_2
X_5634_ _5634_/A VGND VGND VPWR VPWR _5634_/Y sky130_fd_sc_hd__inv_2
X_8422_ _8554_/A _8401_/B _8419_/X _8421_/Y VGND VGND VPWR VPWR _8422_/X sky130_fd_sc_hd__o211a_1
XFILLER_31_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8353_ _8164_/A _8117_/A _8343_/Y _8223_/X _8352_/X VGND VGND VPWR VPWR _8356_/B
+ sky130_fd_sc_hd__o2111ai_4
X_7304_ _7304_/A _7392_/B VGND VGND VPWR VPWR _7304_/X sky130_fd_sc_hd__or2_1
X_5565_ _5565_/A VGND VGND VPWR VPWR _5566_/A sky130_fd_sc_hd__clkbuf_2
X_8284_ _8539_/A _8284_/B VGND VGND VPWR VPWR _8285_/B sky130_fd_sc_hd__or2_1
XFILLER_132_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4516_ _4898_/A _6158_/A VGND VGND VPWR VPWR _4517_/A sky130_fd_sc_hd__or2_2
X_5496_ _5545_/A _5496_/B VGND VGND VPWR VPWR _5497_/A sky130_fd_sc_hd__or2_1
XFILLER_171_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7235_ _6284_/Y _7040_/D _6277_/Y _7110_/X _7234_/X VGND VGND VPWR VPWR _7242_/A
+ sky130_fd_sc_hd__o221a_1
X_4447_ _9570_/Q _4629_/C _9080_/Q VGND VGND VPWR VPWR _8985_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7166_ _6637_/Y _7048_/D _6773_/Y _7040_/B _7165_/X VGND VGND VPWR VPWR _7167_/D
+ sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_1_csclk _9329_/CLK VGND VGND VPWR VPWR _9493_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6117_ _6115_/Y _4564_/B _6116_/Y _4491_/B VGND VGND VPWR VPWR _6117_/X sky130_fd_sc_hd__o22a_2
XFILLER_100_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7097_ _7097_/A VGND VGND VPWR VPWR _7097_/X sky130_fd_sc_hd__buf_8
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6048_ _6050_/A VGND VGND VPWR VPWR _6049_/A sky130_fd_sc_hd__clkbuf_1
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7999_ _8116_/B _8050_/B VGND VGND VPWR VPWR _8000_/A sky130_fd_sc_hd__or2_1
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9738_ _9774_/CLK _9738_/D _9757_/SET_B VGND VGND VPWR VPWR _9738_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_179_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9669_ _9674_/CLK _9669_/D _9633_/SET_B VGND VGND VPWR VPWR _9669_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_10_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_0_0_mgmt_gpio_in[4] clkbuf_2_1_0_mgmt_gpio_in[4]/A VGND VGND VPWR VPWR _8837_/A1
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_110_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5350_ _9480_/Q _5346_/A _8925_/A1 _5346_/Y VGND VGND VPWR VPWR _9480_/D sky130_fd_sc_hd__a22o_1
Xoutput216 _8766_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[17] sky130_fd_sc_hd__buf_2
Xoutput205 _9771_/Q VGND VGND VPWR VPWR irq[0] sky130_fd_sc_hd__buf_2
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput227 _8786_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[27] sky130_fd_sc_hd__buf_2
Xoutput249 _8829_/X VGND VGND VPWR VPWR mgmt_gpio_out[36] sky130_fd_sc_hd__buf_2
Xoutput238 _8835_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[37] sky130_fd_sc_hd__buf_2
X_5281_ _9527_/Q _5280_/A _8846_/X _5280_/Y VGND VGND VPWR VPWR _9527_/D sky130_fd_sc_hd__a22o_1
XFILLER_99_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7020_ _9586_/Q _7020_/B VGND VGND VPWR VPWR _7021_/A sky130_fd_sc_hd__and2b_1
XFILLER_68_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8971_ _8590_/Y _8513_/X _8975_/S VGND VGND VPWR VPWR _8971_/X sky130_fd_sc_hd__mux2_4
XFILLER_83_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7922_ _7836_/B _8299_/B _7862_/Y _7921_/Y VGND VGND VPWR VPWR _7923_/B sky130_fd_sc_hd__a31o_1
XFILLER_36_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7853_ _8521_/B _8270_/B VGND VGND VPWR VPWR _8325_/A sky130_fd_sc_hd__or2_1
XFILLER_23_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7784_ _7897_/A _7898_/B VGND VGND VPWR VPWR _8084_/A sky130_fd_sc_hd__or2_1
XFILLER_168_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6804_ _6799_/Y _5905_/B _6800_/Y _5941_/B _6803_/X VGND VGND VPWR VPWR _6830_/C
+ sky130_fd_sc_hd__o221a_1
X_4996_ _8901_/X _9699_/Q _5001_/S VGND VGND VPWR VPWR _4997_/A sky130_fd_sc_hd__mux2_1
X_9523_ _9684_/CLK _9523_/D _9685_/SET_B VGND VGND VPWR VPWR _9523_/Q sky130_fd_sc_hd__dfrtp_2
X_6735_ _9522_/Q VGND VGND VPWR VPWR _6735_/Y sky130_fd_sc_hd__clkinv_2
X_9454_ _9483_/CLK _9454_/D _9528_/SET_B VGND VGND VPWR VPWR _9454_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_139_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6666_ _6661_/Y _5572_/B _6662_/Y _5556_/B _6665_/X VGND VGND VPWR VPWR _6691_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_164_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5617_ _9297_/Q _5612_/A _8842_/X _5612_/Y VGND VGND VPWR VPWR _9297_/D sky130_fd_sc_hd__a22o_1
X_8405_ _8405_/A VGND VGND VPWR VPWR _8405_/Y sky130_fd_sc_hd__inv_2
X_6597_ _9557_/Q VGND VGND VPWR VPWR _6597_/Y sky130_fd_sc_hd__clkinv_2
X_9385_ _9775_/CLK _9385_/D _7011_/B VGND VGND VPWR VPWR _9385_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_155_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5548_ _9345_/Q _5547_/A _8846_/X _5547_/Y VGND VGND VPWR VPWR _9345_/D sky130_fd_sc_hd__a22o_1
X_8336_ _8673_/A _8336_/B VGND VGND VPWR VPWR _8337_/C sky130_fd_sc_hd__or2_1
X_8267_ _8267_/A _8599_/B VGND VGND VPWR VPWR _8269_/A sky130_fd_sc_hd__or2_1
X_5479_ _9390_/Q _5471_/A _8916_/A1 _5471_/Y VGND VGND VPWR VPWR _9390_/D sky130_fd_sc_hd__a22o_1
XFILLER_132_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7218_ _6430_/Y _7126_/X _6403_/Y _7128_/X VGND VGND VPWR VPWR _7218_/X sky130_fd_sc_hd__o22a_1
XFILLER_78_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8198_ _8525_/A _8583_/B _8583_/C VGND VGND VPWR VPWR _8213_/B sky130_fd_sc_hd__or3_1
XFILLER_132_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7149_ _6919_/Y _7059_/D _6859_/Y _7116_/X _7148_/X VGND VGND VPWR VPWR _7154_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_58_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4850_ _9468_/Q VGND VGND VPWR VPWR _4850_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4781_ _4781_/A VGND VGND VPWR VPWR _4781_/Y sky130_fd_sc_hd__clkinv_2
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6520_ _9180_/Q VGND VGND VPWR VPWR _8747_/A sky130_fd_sc_hd__clkinv_4
XFILLER_33_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6451_ _6451_/A VGND VGND VPWR VPWR _6451_/Y sky130_fd_sc_hd__inv_2
XFILLER_161_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6382_ _6377_/Y _5660_/B _7392_/A _5632_/B _6381_/X VGND VGND VPWR VPWR _6382_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_118_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9170_ _9203_/CLK _9170_/D _9633_/SET_B VGND VGND VPWR VPWR _9170_/Q sky130_fd_sc_hd__dfrtp_1
X_5402_ _9443_/Q _5395_/A _8930_/A1 _5395_/Y VGND VGND VPWR VPWR _9443_/D sky130_fd_sc_hd__a22o_1
XFILLER_173_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8121_ _8397_/A _8397_/B _8098_/A VGND VGND VPWR VPWR _8121_/Y sky130_fd_sc_hd__o21ai_1
X_5333_ _9491_/Q _5330_/A _5965_/B1 _5330_/Y VGND VGND VPWR VPWR _9491_/D sky130_fd_sc_hd__a22o_1
XFILLER_114_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8052_ _8521_/A _8168_/A VGND VGND VPWR VPWR _8392_/A sky130_fd_sc_hd__or2_1
X_5264_ _9538_/Q _5261_/A _5965_/B1 _5261_/Y VGND VGND VPWR VPWR _9538_/D sky130_fd_sc_hd__a22o_1
XFILLER_114_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7003_ _4951_/B _4958_/Y _7003_/C _8958_/X VGND VGND VPWR VPWR _7003_/X sky130_fd_sc_hd__and4bb_1
X_5195_ _9584_/Q _5193_/Y _8904_/X _5193_/A VGND VGND VPWR VPWR _9584_/D sky130_fd_sc_hd__o22a_1
XFILLER_68_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8954_ _7707_/Y _5214_/A _9050_/Q VGND VGND VPWR VPWR _9058_/D sky130_fd_sc_hd__mux2_1
X_7905_ _8496_/A _8077_/A _8341_/B _7896_/A _8498_/A VGND VGND VPWR VPWR _7905_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_83_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8885_ _8884_/X _9143_/Q _9054_/Q VGND VGND VPWR VPWR _8885_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7836_ _7836_/A _7836_/B _7836_/C VGND VGND VPWR VPWR _8662_/A sky130_fd_sc_hd__and3_1
XFILLER_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4979_ _9703_/Q _4966_/A _9702_/Q _4966_/Y VGND VGND VPWR VPWR _9703_/D sky130_fd_sc_hd__a22o_1
X_7767_ _8394_/A _8394_/B _7767_/C VGND VGND VPWR VPWR _7791_/B sky130_fd_sc_hd__or3_2
XFILLER_149_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9506_ _9527_/CLK _9506_/D _9528_/SET_B VGND VGND VPWR VPWR _9506_/Q sky130_fd_sc_hd__dfrtp_1
X_7698_ _7698_/A _7698_/B _7698_/C _7698_/D VGND VGND VPWR VPWR _7698_/Y sky130_fd_sc_hd__nand4_4
X_6718_ _9361_/Q VGND VGND VPWR VPWR _6718_/Y sky130_fd_sc_hd__inv_2
XFILLER_192_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6649_ _6649_/A _6649_/B _6649_/C VGND VGND VPWR VPWR _6785_/A sky130_fd_sc_hd__and3_1
X_9437_ _9514_/CLK _9437_/D _4628_/A VGND VGND VPWR VPWR _9437_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9368_ _9508_/CLK _9368_/D _9295_/SET_B VGND VGND VPWR VPWR _9368_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_124_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_34_csclk clkbuf_2_1_0_csclk/X VGND VGND VPWR VPWR _9620_/CLK sky130_fd_sc_hd__clkbuf_16
X_9299_ _9371_/CLK _9299_/D _9295_/SET_B VGND VGND VPWR VPWR _9299_/Q sky130_fd_sc_hd__dfrtp_1
X_8319_ _8319_/A _8498_/B VGND VGND VPWR VPWR _8493_/C sky130_fd_sc_hd__nor2_1
XFILLER_182_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_49_csclk _9329_/CLK VGND VGND VPWR VPWR _9769_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_115_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5951_ _5951_/A VGND VGND VPWR VPWR _5951_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_1_0_1_mgmt_gpio_in[4] clkbuf_1_0_1_mgmt_gpio_in[4]/A VGND VGND VPWR VPWR clkbuf_2_1_0_mgmt_gpio_in[4]/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_65_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8670_ _8703_/C _8705_/D _8670_/C _8707_/A VGND VGND VPWR VPWR _8671_/C sky130_fd_sc_hd__or4_1
X_4902_ _9432_/Q VGND VGND VPWR VPWR _4902_/Y sky130_fd_sc_hd__inv_2
XFILLER_178_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5882_ _9151_/Q _5874_/A _8916_/A1 _5874_/Y VGND VGND VPWR VPWR _9151_/D sky130_fd_sc_hd__a22o_1
X_4833_ _9416_/Q VGND VGND VPWR VPWR _4833_/Y sky130_fd_sc_hd__inv_4
X_7621_ _4685_/Y _7465_/X _4888_/Y _7467_/X VGND VGND VPWR VPWR _7621_/X sky130_fd_sc_hd__o22a_1
XFILLER_119_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7552_ _6468_/Y _7471_/X _7216_/A _7473_/X _7551_/X VGND VGND VPWR VPWR _7553_/D
+ sky130_fd_sc_hd__o221a_1
X_4764_ _4787_/A _6111_/B VGND VGND VPWR VPWR _5564_/B sky130_fd_sc_hd__or2_2
XFILLER_60_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7483_ _6865_/Y _7408_/X _6913_/Y _7410_/X VGND VGND VPWR VPWR _7483_/X sky130_fd_sc_hd__o22a_1
X_6503_ _9383_/Q VGND VGND VPWR VPWR _6503_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6434_ _9163_/Q VGND VGND VPWR VPWR _6434_/Y sky130_fd_sc_hd__inv_2
X_4695_ _4903_/B _4843_/B VGND VGND VPWR VPWR _5864_/B sky130_fd_sc_hd__or2_4
X_9222_ _9695_/CLK _9222_/D _9779_/SET_B VGND VGND VPWR VPWR _9222_/Q sky130_fd_sc_hd__dfrtp_1
X_6365_ _6360_/Y _5572_/B _6361_/Y _5594_/B _6364_/X VGND VGND VPWR VPWR _6365_/X
+ sky130_fd_sc_hd__o221a_2
X_9153_ _9352_/CLK _9153_/D _9646_/SET_B VGND VGND VPWR VPWR _9153_/Q sky130_fd_sc_hd__dfrtp_1
X_8104_ _7832_/A _8103_/A _7969_/A _8103_/Y VGND VGND VPWR VPWR _8200_/B sky130_fd_sc_hd__a22o_1
X_6296_ _9291_/Q VGND VGND VPWR VPWR _6296_/Y sky130_fd_sc_hd__inv_2
X_5316_ _9502_/Q _5308_/A _8916_/A1 _5308_/Y VGND VGND VPWR VPWR _9502_/D sky130_fd_sc_hd__a22o_1
XFILLER_161_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9084_ _8837_/A1 _9084_/D _6010_/X VGND VGND VPWR VPWR _9084_/Q sky130_fd_sc_hd__dfrtp_2
X_8035_ _8035_/A _8460_/A VGND VGND VPWR VPWR _8035_/X sky130_fd_sc_hd__and2_1
X_5247_ _9549_/Q _5242_/A _5964_/B1 _5242_/Y VGND VGND VPWR VPWR _9549_/D sky130_fd_sc_hd__a22o_1
XFILLER_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5178_ _5960_/A _5178_/B VGND VGND VPWR VPWR _5179_/A sky130_fd_sc_hd__or2_2
XFILLER_68_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8937_ _9087_/Q _9086_/Q _9051_/Q VGND VGND VPWR VPWR _8937_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8868_ _7662_/Y _9629_/Q _8978_/S VGND VGND VPWR VPWR _8868_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8799_ _8799_/A VGND VGND VPWR VPWR _8800_/A sky130_fd_sc_hd__clkbuf_1
XPHY_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7819_ _7819_/A VGND VGND VPWR VPWR _8660_/B sky130_fd_sc_hd__clkbuf_4
XPHY_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4480_ _6111_/A _4931_/A VGND VGND VPWR VPWR _4481_/B sky130_fd_sc_hd__or2_4
X_6150_ _6145_/Y _6149_/A _9043_/Q _6149_/Y VGND VGND VPWR VPWR _9043_/D sky130_fd_sc_hd__o22a_1
XFILLER_143_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5101_ _5101_/A VGND VGND VPWR VPWR _5102_/A sky130_fd_sc_hd__clkbuf_2
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6081_ _6081_/A _6081_/B VGND VGND VPWR VPWR _6081_/X sky130_fd_sc_hd__or2_1
XFILLER_111_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5032_ _6040_/A VGND VGND VPWR VPWR _5033_/A sky130_fd_sc_hd__clkbuf_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater368 _8839_/X VGND VGND VPWR VPWR _5967_/B1 sky130_fd_sc_hd__buf_12
XFILLER_26_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6983_ _6946_/Y _6976_/A _9013_/Q _6976_/Y VGND VGND VPWR VPWR _9013_/D sky130_fd_sc_hd__o22a_1
X_9771_ _9771_/CLK _9771_/D _4628_/A VGND VGND VPWR VPWR _9771_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5934_ _7837_/A _7756_/B VGND VGND VPWR VPWR _5934_/X sky130_fd_sc_hd__or2_1
X_8722_ _8722_/A _8722_/B _8722_/C VGND VGND VPWR VPWR _8723_/B sky130_fd_sc_hd__or3_1
X_8653_ _8638_/Y _8647_/Y _8649_/Y _8652_/X VGND VGND VPWR VPWR _8653_/X sky130_fd_sc_hd__a31o_1
X_5865_ _5865_/A VGND VGND VPWR VPWR _5866_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_80_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7604_ _6065_/Y _7461_/X _6079_/Y _7463_/X _7603_/X VGND VGND VPWR VPWR _7607_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_21_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4816_ _9442_/Q VGND VGND VPWR VPWR _4816_/Y sky130_fd_sc_hd__inv_4
XFILLER_193_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8584_ _8340_/C _8544_/B _8583_/Y _8330_/B _8380_/B VGND VGND VPWR VPWR _8678_/B
+ sky130_fd_sc_hd__a311o_1
X_5796_ _9212_/Q _5791_/A _5967_/B1 _5791_/Y VGND VGND VPWR VPWR _9212_/D sky130_fd_sc_hd__a22o_1
XFILLER_147_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4747_ _4737_/Y _6134_/A _4740_/Y _5818_/B _4746_/X VGND VGND VPWR VPWR _4747_/X
+ sky130_fd_sc_hd__o221a_1
X_7535_ _7535_/A _7535_/B _7535_/C _7535_/D VGND VGND VPWR VPWR _7536_/D sky130_fd_sc_hd__and4_1
XFILLER_181_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7466_ _7466_/A _7476_/C _7474_/D VGND VGND VPWR VPWR _7467_/A sky130_fd_sc_hd__or3_1
X_4678_ _4921_/A _4843_/B VGND VGND VPWR VPWR _5080_/B sky130_fd_sc_hd__or2_4
X_9205_ _9613_/CLK _9205_/D _9646_/SET_B VGND VGND VPWR VPWR _9205_/Q sky130_fd_sc_hd__dfstp_1
X_6417_ _9436_/Q VGND VGND VPWR VPWR _6417_/Y sky130_fd_sc_hd__inv_2
X_7397_ _7397_/A _7397_/B _7397_/C VGND VGND VPWR VPWR _7397_/Y sky130_fd_sc_hd__nand3_4
X_9136_ _9354_/CLK _9136_/D _9685_/SET_B VGND VGND VPWR VPWR _9136_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_122_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6348_ _9441_/Q VGND VGND VPWR VPWR _6348_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_163_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput127 user_clock VGND VGND VPWR VPWR _4449_/A1 sky130_fd_sc_hd__buf_2
X_9067_ _4450_/A1 _9067_/D _6146_/A VGND VGND VPWR VPWR _9067_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_142_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6279_ _6274_/Y _5382_/B _6275_/Y _5267_/B _6278_/X VGND VGND VPWR VPWR _6280_/D
+ sky130_fd_sc_hd__o221a_2
Xinput116 sram_ro_data[30] VGND VGND VPWR VPWR _6227_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_48_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput105 sram_ro_data[20] VGND VGND VPWR VPWR _6438_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput149 wb_adr_i[25] VGND VGND VPWR VPWR input149/X sky130_fd_sc_hd__clkbuf_1
Xinput138 wb_adr_i[15] VGND VGND VPWR VPWR _7770_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_130_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8018_ _8624_/B _8401_/A VGND VGND VPWR VPWR _8441_/B sky130_fd_sc_hd__or2_1
XFILLER_29_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5650_ _9054_/Q _6997_/C _9056_/Q VGND VGND VPWR VPWR _5651_/B sky130_fd_sc_hd__a21o_1
XFILLER_175_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4601_ _6111_/A _4921_/A VGND VGND VPWR VPWR _4602_/B sky130_fd_sc_hd__or2_4
XFILLER_191_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5581_ _9321_/Q _5574_/A _8930_/A1 _5574_/Y VGND VGND VPWR VPWR _9321_/D sky130_fd_sc_hd__a22o_1
XFILLER_156_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7320_ _6897_/Y _7048_/D _6833_/Y _7040_/B _7319_/X VGND VGND VPWR VPWR _7321_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4532_ _9764_/Q _4526_/A _5965_/B1 _4526_/Y VGND VGND VPWR VPWR _9764_/D sky130_fd_sc_hd__a22o_1
XFILLER_183_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7251_ _6190_/Y _7079_/B _6179_/Y _7059_/A VGND VGND VPWR VPWR _7251_/X sky130_fd_sc_hd__o22a_1
X_4463_ _6111_/A _4919_/A VGND VGND VPWR VPWR _6251_/A sky130_fd_sc_hd__or2_4
XFILLER_117_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6202_ _9738_/Q VGND VGND VPWR VPWR _6202_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7182_ _8749_/A _7048_/B _8745_/A _7077_/A _7181_/X VGND VGND VPWR VPWR _7189_/A
+ sky130_fd_sc_hd__o221a_1
X_6133_ _9345_/Q VGND VGND VPWR VPWR _6133_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6064_ _6059_/Y _5968_/B _8807_/B _6165_/A _6063_/X VGND VGND VPWR VPWR _6071_/A
+ sky130_fd_sc_hd__o221a_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5015_ _5015_/A VGND VGND VPWR VPWR _5015_/Y sky130_fd_sc_hd__inv_2
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6966_ _6237_/Y _6964_/A _9026_/Q _6964_/Y VGND VGND VPWR VPWR _9026_/D sky130_fd_sc_hd__o22a_1
XFILLER_81_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9754_ _9755_/CLK _9754_/D _9757_/SET_B VGND VGND VPWR VPWR _9754_/Q sky130_fd_sc_hd__dfstp_1
X_8705_ _8705_/A _8705_/B _8705_/C _8705_/D VGND VGND VPWR VPWR _8706_/D sky130_fd_sc_hd__or4_1
X_5917_ _5917_/A VGND VGND VPWR VPWR _5918_/A sky130_fd_sc_hd__clkbuf_2
X_9685_ _9687_/CLK _9685_/D _9685_/SET_B VGND VGND VPWR VPWR _9685_/Q sky130_fd_sc_hd__dfstp_1
X_6897_ _9199_/Q VGND VGND VPWR VPWR _6897_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_42_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8636_ _8636_/A _8636_/B _8636_/C _8636_/D VGND VGND VPWR VPWR _8714_/C sky130_fd_sc_hd__or4_2
X_5848_ _8924_/X VGND VGND VPWR VPWR _5849_/A sky130_fd_sc_hd__clkinv_4
XFILLER_139_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8567_ _8640_/A _8566_/Y _8352_/A VGND VGND VPWR VPWR _8641_/B sky130_fd_sc_hd__o21ai_2
X_5779_ _9225_/Q _5778_/A _8846_/X _5778_/Y VGND VGND VPWR VPWR _9225_/D sky130_fd_sc_hd__a22o_1
XFILLER_166_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7518_ _7518_/A _7518_/B _7518_/C _7518_/D VGND VGND VPWR VPWR _7518_/Y sky130_fd_sc_hd__nand4_4
XFILLER_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8498_ _8498_/A _8498_/B VGND VGND VPWR VPWR _8695_/A sky130_fd_sc_hd__nor2_1
XFILLER_162_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7449_ _4779_/Y _7441_/X _4850_/Y _7443_/X _7448_/X VGND VGND VPWR VPWR _7480_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_107_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9119_ _4450_/A1 _9119_/D _6146_/A VGND VGND VPWR VPWR _9119_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6820_ _6820_/A VGND VGND VPWR VPWR _6820_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6751_ input37/X _8930_/S _6750_/Y _5897_/B VGND VGND VPWR VPWR _6751_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_176_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9470_ _9687_/CLK _9470_/D _9528_/SET_B VGND VGND VPWR VPWR _9470_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_1_1_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
X_6682_ _9187_/Q VGND VGND VPWR VPWR _6682_/Y sky130_fd_sc_hd__clkinv_4
X_5702_ _5696_/Y _5701_/X _5692_/A VGND VGND VPWR VPWR _9254_/D sky130_fd_sc_hd__o21a_1
X_5633_ _5633_/A VGND VGND VPWR VPWR _5634_/A sky130_fd_sc_hd__clkbuf_2
X_8421_ _8630_/C VGND VGND VPWR VPWR _8421_/Y sky130_fd_sc_hd__inv_2
X_8352_ _8352_/A _8352_/B _8352_/C VGND VGND VPWR VPWR _8352_/X sky130_fd_sc_hd__and3_1
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5564_ _5671_/A _5564_/B VGND VGND VPWR VPWR _5565_/A sky130_fd_sc_hd__or2_1
XFILLER_191_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7303_ _4765_/Y _7059_/D _4920_/Y _7116_/X _7302_/X VGND VGND VPWR VPWR _7308_/B
+ sky130_fd_sc_hd__o221a_1
X_4515_ _4515_/A VGND VGND VPWR VPWR _6158_/A sky130_fd_sc_hd__buf_8
X_8283_ _8283_/A _8330_/B VGND VGND VPWR VPWR _8284_/B sky130_fd_sc_hd__or2_1
X_5495_ _9380_/Q _5490_/A _5967_/B1 _5490_/Y VGND VGND VPWR VPWR _9380_/D sky130_fd_sc_hd__a22o_1
XFILLER_132_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7234_ _6320_/Y _7112_/X _6302_/Y _7077_/B VGND VGND VPWR VPWR _7234_/X sky130_fd_sc_hd__o22a_1
X_4446_ _9571_/Q _4446_/A1 _9682_/Q VGND VGND VPWR VPWR _8986_/A sky130_fd_sc_hd__mux2_1
X_7165_ _6639_/Y _7068_/A _6761_/Y _7105_/X VGND VGND VPWR VPWR _7165_/X sky130_fd_sc_hd__o22a_1
XFILLER_98_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6116_ _9785_/Q VGND VGND VPWR VPWR _6116_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7096_ _7127_/C _7096_/B VGND VGND VPWR VPWR _7097_/A sky130_fd_sc_hd__or2_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6047_ _6047_/A VGND VGND VPWR VPWR _6047_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_39_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7998_ _7998_/A VGND VGND VPWR VPWR _8401_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6949_ _9063_/Q VGND VGND VPWR VPWR _6950_/B sky130_fd_sc_hd__inv_2
X_9737_ _9774_/CLK _9737_/D _9757_/SET_B VGND VGND VPWR VPWR _9737_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9668_ _9674_/CLK _9668_/D _9779_/SET_B VGND VGND VPWR VPWR _9668_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_179_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8619_ _8619_/A _8707_/A _8706_/B _8619_/D VGND VGND VPWR VPWR _8620_/D sky130_fd_sc_hd__or4_1
X_9599_ _9601_/CLK _9599_/D _9528_/SET_B VGND VGND VPWR VPWR _9599_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_155_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput217 _8768_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[18] sky130_fd_sc_hd__buf_2
Xoutput206 _8807_/Y VGND VGND VPWR VPWR irq[1] sky130_fd_sc_hd__buf_2
Xoutput228 _8788_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[28] sky130_fd_sc_hd__buf_2
X_5280_ _5280_/A VGND VGND VPWR VPWR _5280_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput239 _7706_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[3] sky130_fd_sc_hd__buf_2
XFILLER_141_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8970_ _8488_/X _8338_/X _8975_/S VGND VGND VPWR VPWR _8970_/X sky130_fd_sc_hd__mux2_4
XFILLER_95_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7921_ _8077_/A _8262_/B _7920_/X VGND VGND VPWR VPWR _7921_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7852_ _7852_/A VGND VGND VPWR VPWR _8270_/B sky130_fd_sc_hd__clkbuf_2
X_7783_ _7969_/A _7777_/Y _7832_/A _7777_/A _8218_/A VGND VGND VPWR VPWR _7898_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_90_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6803_ _6801_/Y _5518_/B _6802_/Y _5602_/B _6158_/X VGND VGND VPWR VPWR _6803_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4995_ _4995_/A VGND VGND VPWR VPWR _4995_/X sky130_fd_sc_hd__clkbuf_1
X_9522_ _9527_/CLK _9522_/D _9528_/SET_B VGND VGND VPWR VPWR _9522_/Q sky130_fd_sc_hd__dfrtp_1
X_6734_ _6729_/Y _5366_/B _6730_/Y _5298_/B _6733_/X VGND VGND VPWR VPWR _6741_/C
+ sky130_fd_sc_hd__o221a_1
X_9453_ _9483_/CLK _9453_/D _9528_/SET_B VGND VGND VPWR VPWR _9453_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_164_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6665_ _7348_/A _5632_/B _6664_/Y _5679_/B VGND VGND VPWR VPWR _6665_/X sky130_fd_sc_hd__o22a_1
X_8404_ _8665_/B _8571_/A VGND VGND VPWR VPWR _8405_/A sky130_fd_sc_hd__or2_1
XFILLER_191_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5616_ _9298_/Q _5612_/A _8925_/A1 _5612_/Y VGND VGND VPWR VPWR _9298_/D sky130_fd_sc_hd__a22o_1
X_9384_ _9771_/CLK _9384_/D _4628_/A VGND VGND VPWR VPWR _9384_/Q sky130_fd_sc_hd__dfrtp_1
X_6596_ _6591_/Y _4564_/B _6592_/Y _6086_/X _6595_/X VGND VGND VPWR VPWR _6596_/X
+ sky130_fd_sc_hd__o221a_1
X_5547_ _5547_/A VGND VGND VPWR VPWR _5547_/Y sky130_fd_sc_hd__inv_2
X_8335_ _8335_/A _8334_/X VGND VGND VPWR VPWR _8336_/B sky130_fd_sc_hd__or2b_1
XFILLER_105_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5478_ _9391_/Q _5471_/A _8840_/X _5471_/Y VGND VGND VPWR VPWR _9391_/D sky130_fd_sc_hd__a22o_1
XFILLER_155_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8266_ _8510_/A _8270_/B VGND VGND VPWR VPWR _8599_/B sky130_fd_sc_hd__nor2_1
XFILLER_132_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7217_ _6422_/Y _5728_/X _6334_/Y _7040_/A _7216_/X VGND VGND VPWR VPWR _7220_/C
+ sky130_fd_sc_hd__o221a_1
X_8197_ _8346_/A _8346_/B _8196_/X VGND VGND VPWR VPWR _8583_/C sky130_fd_sc_hd__o21ai_2
XFILLER_132_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7148_ _6788_/Y _7118_/X _6915_/Y _7048_/C VGND VGND VPWR VPWR _7148_/X sky130_fd_sc_hd__o22a_1
XFILLER_100_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7079_ _7127_/C _7079_/B _7079_/C _7079_/D VGND VGND VPWR VPWR _7080_/A sky130_fd_sc_hd__and4_1
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4780_ _6086_/B _4780_/B VGND VGND VPWR VPWR _5757_/B sky130_fd_sc_hd__or2_4
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_0_csclk _9329_/CLK VGND VGND VPWR VPWR _9545_/CLK sky130_fd_sc_hd__clkbuf_16
X_6450_ _6450_/A VGND VGND VPWR VPWR _6450_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_146_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6381_ _6379_/Y _5671_/B _7216_/A _5610_/B VGND VGND VPWR VPWR _6381_/X sky130_fd_sc_hd__o22a_1
X_5401_ _9444_/Q _5395_/A _5965_/B1 _5395_/Y VGND VGND VPWR VPWR _9444_/D sky130_fd_sc_hd__a22o_1
X_8120_ _8120_/A _8120_/B VGND VGND VPWR VPWR _8397_/B sky130_fd_sc_hd__or2_4
XFILLER_173_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5332_ _9492_/Q _5330_/A _5964_/B1 _5330_/Y VGND VGND VPWR VPWR _9492_/D sky130_fd_sc_hd__a22o_1
XFILLER_141_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8051_ _8051_/A VGND VGND VPWR VPWR _8168_/A sky130_fd_sc_hd__buf_2
XFILLER_114_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5263_ _9539_/Q _5261_/A _5964_/B1 _5261_/Y VGND VGND VPWR VPWR _9539_/D sky130_fd_sc_hd__a22o_1
X_7002_ _7002_/A VGND VGND VPWR VPWR _9059_/D sky130_fd_sc_hd__clkbuf_1
X_5194_ _9585_/Q _5193_/Y _8914_/X _5193_/A VGND VGND VPWR VPWR _9585_/D sky130_fd_sc_hd__o22a_1
XFILLER_83_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8953_ _9717_/Q _6145_/Y _8957_/S VGND VGND VPWR VPWR _8953_/X sky130_fd_sc_hd__mux2_1
X_7904_ _7904_/A VGND VGND VPWR VPWR _8498_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_70_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8884_ _7265_/Y _9638_/Q _8959_/S VGND VGND VPWR VPWR _8884_/X sky130_fd_sc_hd__mux2_1
X_7835_ _8496_/A VGND VGND VPWR VPWR _7836_/B sky130_fd_sc_hd__inv_4
XFILLER_24_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4978_ _4978_/A VGND VGND VPWR VPWR _4978_/X sky130_fd_sc_hd__clkbuf_1
X_9505_ _9527_/CLK _9505_/D _9528_/SET_B VGND VGND VPWR VPWR _9505_/Q sky130_fd_sc_hd__dfrtp_1
X_7766_ _7838_/B VGND VGND VPWR VPWR _7767_/C sky130_fd_sc_hd__inv_2
XFILLER_24_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6717_ _9496_/Q VGND VGND VPWR VPWR _6717_/Y sky130_fd_sc_hd__clkinv_2
X_7697_ _7697_/A _7697_/B _7697_/C _7697_/D VGND VGND VPWR VPWR _7698_/D sky130_fd_sc_hd__and4_1
XFILLER_192_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6648_ _6643_/Y _5757_/B _6644_/Y _5818_/B _6647_/X VGND VGND VPWR VPWR _6649_/C
+ sky130_fd_sc_hd__o221a_1
X_9436_ _9440_/CLK _9436_/D _4628_/A VGND VGND VPWR VPWR _9436_/Q sky130_fd_sc_hd__dfrtp_1
X_9367_ _9371_/CLK _9367_/D _9295_/SET_B VGND VGND VPWR VPWR _9367_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_125_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6579_ _6574_/Y _5298_/B _8767_/A _5496_/B _6578_/X VGND VGND VPWR VPWR _6586_/B
+ sky130_fd_sc_hd__o221a_1
X_8318_ _8318_/A _8490_/C _8597_/C VGND VGND VPWR VPWR _8318_/X sky130_fd_sc_hd__or3_1
X_9298_ _9788_/CLK _9298_/D _9295_/SET_B VGND VGND VPWR VPWR _9298_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_182_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8249_ _8510_/A _8254_/B VGND VGND VPWR VPWR _8250_/A sky130_fd_sc_hd__or2_1
XFILLER_120_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5950_ _5950_/A VGND VGND VPWR VPWR _5951_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_80_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4901_ _4901_/A VGND VGND VPWR VPWR _4901_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5881_ _9152_/Q _5874_/A _8930_/A1 _5874_/Y VGND VGND VPWR VPWR _9152_/D sky130_fd_sc_hd__a22o_1
X_7620_ _4761_/Y _7451_/X _4899_/Y _7453_/X _7619_/X VGND VGND VPWR VPWR _7625_/B
+ sky130_fd_sc_hd__o221a_1
XANTENNA_190 _6271_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4832_ _6111_/A _6086_/B VGND VGND VPWR VPWR _4832_/X sky130_fd_sc_hd__or2_4
XFILLER_193_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7551_ _6430_/Y _7475_/X _6377_/Y _7477_/X VGND VGND VPWR VPWR _7551_/X sky130_fd_sc_hd__o22a_1
X_4763_ _9328_/Q VGND VGND VPWR VPWR _4763_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6502_ _9234_/Q VGND VGND VPWR VPWR _8755_/A sky130_fd_sc_hd__inv_6
X_4694_ _9159_/Q VGND VGND VPWR VPWR _4694_/Y sky130_fd_sc_hd__clkinv_4
X_7482_ _7482_/A VGND VGND VPWR VPWR _7482_/X sky130_fd_sc_hd__clkbuf_1
X_6433_ _6433_/A _6433_/B _6433_/C _6433_/D VGND VGND VPWR VPWR _6474_/B sky130_fd_sc_hd__and4_1
X_9221_ _9695_/CLK _9221_/D _9779_/SET_B VGND VGND VPWR VPWR _9221_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6364_ _6362_/Y _5742_/B _6363_/Y _5556_/B VGND VGND VPWR VPWR _6364_/X sky130_fd_sc_hd__o22a_1
X_9152_ _9352_/CLK _9152_/D _9646_/SET_B VGND VGND VPWR VPWR _9152_/Q sky130_fd_sc_hd__dfstp_1
X_8103_ _8103_/A VGND VGND VPWR VPWR _8103_/Y sky130_fd_sc_hd__inv_2
X_5315_ _9503_/Q _5308_/A _8840_/X _5308_/Y VGND VGND VPWR VPWR _9503_/D sky130_fd_sc_hd__a22o_1
XFILLER_130_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6295_ _6287_/Y _5545_/B _6288_/Y _5797_/B _6294_/X VGND VGND VPWR VPWR _6307_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_114_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9083_ _9709_/CLK _9083_/D _6013_/X VGND VGND VPWR VPWR _9083_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_114_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8034_ _8624_/B _8551_/A VGND VGND VPWR VPWR _8460_/A sky130_fd_sc_hd__or2_1
X_5246_ _9550_/Q _5242_/A _5963_/B1 _5242_/Y VGND VGND VPWR VPWR _9550_/D sky130_fd_sc_hd__a22o_1
XFILLER_102_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5177_ _9594_/Q _5169_/A _8916_/A1 _5169_/Y VGND VGND VPWR VPWR _9594_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8936_ _8935_/X _9679_/Q _9587_/Q VGND VGND VPWR VPWR _8936_/X sky130_fd_sc_hd__mux2_2
XFILLER_169_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8867_ _8866_/X _9172_/Q _9054_/Q VGND VGND VPWR VPWR _8867_/X sky130_fd_sc_hd__mux2_1
X_8798_ _8798_/A VGND VGND VPWR VPWR _8798_/X sky130_fd_sc_hd__clkbuf_1
XPHY_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7818_ _7903_/C _8528_/A _8583_/A _7894_/B VGND VGND VPWR VPWR _7819_/A sky130_fd_sc_hd__or4_1
X_7749_ _9068_/Q _7749_/A2 _9067_/Q _7749_/B2 _7748_/X VGND VGND VPWR VPWR _7749_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_184_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9419_ _9684_/CLK _9419_/D _9685_/SET_B VGND VGND VPWR VPWR _9419_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_165_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6080_ _9397_/Q VGND VGND VPWR VPWR _6081_/A sky130_fd_sc_hd__clkinv_2
X_5100_ _5259_/A _5100_/B VGND VGND VPWR VPWR _5101_/A sky130_fd_sc_hd__or2_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5031_ _9683_/Q _5026_/A _8839_/X _5026_/Y VGND VGND VPWR VPWR _9683_/D sky130_fd_sc_hd__a22o_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater369 _8839_/X VGND VGND VPWR VPWR _8916_/A1 sky130_fd_sc_hd__buf_12
X_9770_ _9770_/CLK _9770_/D _7011_/B VGND VGND VPWR VPWR _9770_/Q sky130_fd_sc_hd__dfrtp_1
X_8721_ _8721_/A _8721_/B _8721_/C _8721_/D VGND VGND VPWR VPWR _8722_/C sky130_fd_sc_hd__or4_1
X_6982_ _6785_/Y _6976_/A _9014_/Q _6976_/Y VGND VGND VPWR VPWR _9014_/D sky130_fd_sc_hd__o22a_1
XFILLER_65_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5933_ _7837_/B VGND VGND VPWR VPWR _7756_/B sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_33_csclk clkbuf_2_1_0_csclk/X VGND VGND VPWR VPWR _9674_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_178_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8652_ _8681_/A _8722_/B _8681_/C VGND VGND VPWR VPWR _8652_/X sky130_fd_sc_hd__or3_1
X_5864_ _5960_/A _5864_/B VGND VGND VPWR VPWR _5865_/A sky130_fd_sc_hd__or2_1
X_8583_ _8583_/A _8583_/B _8583_/C VGND VGND VPWR VPWR _8583_/Y sky130_fd_sc_hd__nor3_1
X_7603_ _6121_/Y _7465_/X _6073_/Y _7467_/X VGND VGND VPWR VPWR _7603_/X sky130_fd_sc_hd__o22a_1
X_4815_ _4911_/A _6158_/B VGND VGND VPWR VPWR _6027_/B sky130_fd_sc_hd__or2_4
XFILLER_193_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7534_ _7699_/A _7471_/X _8761_/A _7473_/X _7533_/X VGND VGND VPWR VPWR _7535_/D
+ sky130_fd_sc_hd__o221a_1
X_5795_ _9213_/Q _5791_/A _8930_/A1 _5791_/Y VGND VGND VPWR VPWR _9213_/D sky130_fd_sc_hd__a22o_1
X_4746_ _4742_/Y _5572_/B _4744_/Y _6081_/B VGND VGND VPWR VPWR _4746_/X sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_48_csclk _9329_/CLK VGND VGND VPWR VPWR _9774_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_174_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7465_ _7465_/A VGND VGND VPWR VPWR _7465_/X sky130_fd_sc_hd__buf_8
X_4677_ _9654_/Q VGND VGND VPWR VPWR _4677_/Y sky130_fd_sc_hd__clkinv_2
X_9204_ _9652_/CLK _9204_/D _9647_/SET_B VGND VGND VPWR VPWR _9204_/Q sky130_fd_sc_hd__dfstp_1
X_7396_ _7396_/A _7396_/B _7396_/C _7396_/D VGND VGND VPWR VPWR _7397_/C sky130_fd_sc_hd__and4_1
X_6416_ _9118_/Q VGND VGND VPWR VPWR _6416_/Y sky130_fd_sc_hd__inv_2
XFILLER_162_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9135_ _9354_/CLK _9135_/D _9685_/SET_B VGND VGND VPWR VPWR _9135_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_115_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6347_ _9493_/Q VGND VGND VPWR VPWR _6347_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_163_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9066_ _4450_/A1 _9066_/D _6146_/A VGND VGND VPWR VPWR _9066_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_102_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6278_ _6276_/Y _5496_/B _6277_/Y _5534_/B VGND VGND VPWR VPWR _6278_/X sky130_fd_sc_hd__o22a_1
Xinput117 sram_ro_data[31] VGND VGND VPWR VPWR _6097_/A sky130_fd_sc_hd__clkbuf_1
Xinput106 sram_ro_data[21] VGND VGND VPWR VPWR _6252_/A sky130_fd_sc_hd__clkbuf_1
Xinput128 usr1_vcc_pwrgood VGND VGND VPWR VPWR _6593_/A sky130_fd_sc_hd__clkbuf_1
Xinput139 wb_adr_i[16] VGND VGND VPWR VPWR _7768_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_130_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8017_ _8521_/A _8401_/A VGND VGND VPWR VPWR _8019_/C sky130_fd_sc_hd__or2_1
XFILLER_29_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5229_ _5229_/A VGND VGND VPWR VPWR _9560_/D sky130_fd_sc_hd__clkbuf_1
X_8919_ _9603_/Q _8840_/X _8926_/S VGND VGND VPWR VPWR _8919_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_90 _8817_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_3_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_121_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4600_ _9732_/Q _4592_/A _5967_/B1 _4592_/Y VGND VGND VPWR VPWR _9732_/D sky130_fd_sc_hd__a22o_1
X_5580_ _9322_/Q _5574_/A _8955_/A1 _5574_/Y VGND VGND VPWR VPWR _9322_/D sky130_fd_sc_hd__a22o_1
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4531_ _9765_/Q _4526_/A _5964_/B1 _4526_/Y VGND VGND VPWR VPWR _9765_/D sky130_fd_sc_hd__a22o_1
X_7250_ _6196_/Y _7095_/X _6183_/Y _7068_/D _7249_/X VGND VGND VPWR VPWR _7255_/B
+ sky130_fd_sc_hd__o221a_1
X_4462_ _4729_/A _4729_/B _8934_/X _8932_/X VGND VGND VPWR VPWR _4919_/A sky130_fd_sc_hd__or4_4
X_6201_ _9396_/Q VGND VGND VPWR VPWR _6201_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_144_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7181_ _8743_/A _7040_/C _7701_/A _7059_/C VGND VGND VPWR VPWR _7181_/X sky130_fd_sc_hd__o22a_1
X_6132_ _6132_/A VGND VGND VPWR VPWR _6132_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6063_ _6061_/Y _5583_/B _6062_/Y _5089_/B VGND VGND VPWR VPWR _6063_/X sky130_fd_sc_hd__o22a_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5014_ _5014_/A VGND VGND VPWR VPWR _5015_/A sky130_fd_sc_hd__buf_2
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6965_ _6145_/Y _6964_/A _9027_/Q _6964_/Y VGND VGND VPWR VPWR _9027_/D sky130_fd_sc_hd__o22a_1
X_9753_ _9755_/CLK _9753_/D _9757_/SET_B VGND VGND VPWR VPWR _9753_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_26_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9684_ _9684_/CLK _9684_/D _9685_/SET_B VGND VGND VPWR VPWR _9684_/Q sky130_fd_sc_hd__dfrtp_1
X_8704_ _8704_/A _8704_/B VGND VGND VPWR VPWR _8705_/C sky130_fd_sc_hd__or2_1
X_5916_ _5960_/A _5916_/B VGND VGND VPWR VPWR _5917_/A sky130_fd_sc_hd__or2_1
XFILLER_167_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6896_ _9134_/Q VGND VGND VPWR VPWR _6896_/Y sky130_fd_sc_hd__clkinv_2
X_8635_ _8713_/B _8714_/A VGND VGND VPWR VPWR _8635_/Y sky130_fd_sc_hd__nor2_1
XFILLER_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5847_ _9177_/Q _5839_/A _8916_/A1 _5839_/Y VGND VGND VPWR VPWR _9177_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8566_ _8566_/A _8566_/B VGND VGND VPWR VPWR _8566_/Y sky130_fd_sc_hd__nor2_1
X_5778_ _5778_/A VGND VGND VPWR VPWR _5778_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_21_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8497_ _8497_/A _8395_/X VGND VGND VPWR VPWR _8501_/C sky130_fd_sc_hd__or2b_1
X_7517_ _7517_/A _7517_/B _7517_/C _7517_/D VGND VGND VPWR VPWR _7518_/D sky130_fd_sc_hd__and4_2
X_4729_ _4729_/A _4729_/B _8934_/X _4729_/D VGND VGND VPWR VPWR _4900_/B sky130_fd_sc_hd__or4_4
X_7448_ _4914_/Y _7445_/X _4928_/Y _7447_/X VGND VGND VPWR VPWR _7448_/X sky130_fd_sc_hd__o22a_1
XFILLER_107_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7379_ _6464_/Y _7040_/C _6331_/Y _7059_/C VGND VGND VPWR VPWR _7379_/X sky130_fd_sc_hd__o22a_1
X_9118_ _9779_/CLK _9118_/D _9779_/SET_B VGND VGND VPWR VPWR _9118_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9049_ _9709_/CLK _9049_/D _6049_/X VGND VGND VPWR VPWR _9049_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_49_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6750_ _9135_/Q VGND VGND VPWR VPWR _6750_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5701_ _9253_/Q _7462_/A _5724_/B _9254_/Q VGND VGND VPWR VPWR _5701_/X sky130_fd_sc_hd__o31a_1
X_6681_ _9690_/Q VGND VGND VPWR VPWR _6681_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5632_ _5671_/A _5632_/B VGND VGND VPWR VPWR _5633_/A sky130_fd_sc_hd__or2_1
X_8420_ _8615_/B _8578_/A VGND VGND VPWR VPWR _8630_/C sky130_fd_sc_hd__or2_1
X_5563_ _9333_/Q _5558_/A _8839_/X _5558_/Y VGND VGND VPWR VPWR _9333_/D sky130_fd_sc_hd__a22o_1
XFILLER_136_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8351_ _8640_/A _8378_/B _8640_/C VGND VGND VPWR VPWR _8352_/C sky130_fd_sc_hd__or3_1
XFILLER_129_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7302_ _4800_/Y _7118_/X _4786_/Y _7048_/C VGND VGND VPWR VPWR _7302_/X sky130_fd_sc_hd__o22a_1
X_4514_ _8936_/X _8938_/X _4665_/C VGND VGND VPWR VPWR _4515_/A sky130_fd_sc_hd__or3_1
X_8282_ _8625_/A _8282_/B _8282_/C VGND VGND VPWR VPWR _8330_/B sky130_fd_sc_hd__and3_1
X_5494_ _9381_/Q _5490_/A _5966_/B1 _5490_/Y VGND VGND VPWR VPWR _9381_/D sky130_fd_sc_hd__a22o_1
X_7233_ _7233_/A _7233_/B _7233_/C _7233_/D VGND VGND VPWR VPWR _7243_/B sky130_fd_sc_hd__and4_1
X_4445_ _9572_/Q _4949_/A _9682_/Q VGND VGND VPWR VPWR _8987_/A sky130_fd_sc_hd__mux2_1
X_7164_ _6748_/Y _7059_/B _6753_/Y _7068_/C _7163_/X VGND VGND VPWR VPWR _7167_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_98_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6115_ _9755_/Q VGND VGND VPWR VPWR _6115_/Y sky130_fd_sc_hd__inv_2
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7095_ _7095_/A VGND VGND VPWR VPWR _7095_/X sky130_fd_sc_hd__buf_8
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6046_ _6050_/A VGND VGND VPWR VPWR _6047_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7997_ _8116_/B _7997_/B VGND VGND VPWR VPWR _7998_/A sky130_fd_sc_hd__or2_1
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6948_ _4936_/Y _6149_/A _9036_/Q _6149_/Y VGND VGND VPWR VPWR _9036_/D sky130_fd_sc_hd__o22a_1
XFILLER_169_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9736_ _9774_/CLK _9736_/D _9757_/SET_B VGND VGND VPWR VPWR _9736_/Q sky130_fd_sc_hd__dfstp_1
X_6879_ _9205_/Q VGND VGND VPWR VPWR _6879_/Y sky130_fd_sc_hd__inv_2
X_9667_ _9674_/CLK _9667_/D _9779_/SET_B VGND VGND VPWR VPWR _9667_/Q sky130_fd_sc_hd__dfstp_1
X_9598_ _9601_/CLK _9598_/D _9528_/SET_B VGND VGND VPWR VPWR _9598_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8618_ _8515_/A _8305_/A _8521_/A _8515_/A VGND VGND VPWR VPWR _8706_/B sky130_fd_sc_hd__o22ai_2
XFILLER_139_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8549_ _8130_/B _8554_/B _8137_/B _8554_/B _8548_/X VGND VGND VPWR VPWR _8553_/A
+ sky130_fd_sc_hd__o221ai_1
XFILLER_185_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput207 _8808_/Y VGND VGND VPWR VPWR irq[2] sky130_fd_sc_hd__buf_2
Xoutput218 _8770_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[19] sky130_fd_sc_hd__buf_2
Xoutput229 _8790_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[29] sky130_fd_sc_hd__buf_2
XFILLER_181_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7920_ _7864_/X _8319_/A _7917_/Y _8492_/A _8320_/A VGND VGND VPWR VPWR _7920_/X
+ sky130_fd_sc_hd__o2111a_1
X_7851_ _8324_/A _8496_/A VGND VGND VPWR VPWR _7852_/A sky130_fd_sc_hd__or2_1
X_6802_ _9303_/Q VGND VGND VPWR VPWR _6802_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_36_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7782_ _7832_/A _7837_/B _7781_/Y _7837_/C _5934_/X VGND VGND VPWR VPWR _8218_/A
+ sky130_fd_sc_hd__a32o_2
X_4994_ _4994_/A VGND VGND VPWR VPWR _4995_/A sky130_fd_sc_hd__clkbuf_1
X_9521_ _9684_/CLK _9521_/D _9685_/SET_B VGND VGND VPWR VPWR _9521_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_51_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6733_ _6731_/Y _5960_/B _6732_/Y _5080_/B VGND VGND VPWR VPWR _6733_/X sky130_fd_sc_hd__o22a_1
X_9452_ _9483_/CLK _9452_/D _9685_/SET_B VGND VGND VPWR VPWR _9452_/Q sky130_fd_sc_hd__dfrtp_1
X_6664_ _9258_/Q VGND VGND VPWR VPWR _6664_/Y sky130_fd_sc_hd__clkinv_4
X_5615_ _9299_/Q _5612_/A _8844_/X _5612_/Y VGND VGND VPWR VPWR _9299_/D sky130_fd_sc_hd__a22o_1
X_8403_ _8403_/A VGND VGND VPWR VPWR _8665_/B sky130_fd_sc_hd__inv_2
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6595_ _6593_/Y _4868_/X _8795_/A _5431_/B VGND VGND VPWR VPWR _6595_/X sky130_fd_sc_hd__o22a_4
X_9383_ _9771_/CLK _9383_/D _4628_/A VGND VGND VPWR VPWR _9383_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_191_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5546_ _5546_/A VGND VGND VPWR VPWR _5547_/A sky130_fd_sc_hd__clkbuf_4
X_8334_ _8202_/A _8510_/A _8660_/A _8202_/A VGND VGND VPWR VPWR _8334_/X sky130_fd_sc_hd__o22a_1
X_5477_ _9392_/Q _5471_/A _8841_/X _5471_/Y VGND VGND VPWR VPWR _9392_/D sky130_fd_sc_hd__a22o_1
XFILLER_155_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8265_ _8265_/A _8645_/B VGND VGND VPWR VPWR _8267_/A sky130_fd_sc_hd__or2_1
XFILLER_2_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7216_ _7216_/A _7392_/B VGND VGND VPWR VPWR _7216_/X sky130_fd_sc_hd__or2_1
X_8196_ _7903_/C _8195_/Y _7839_/A _7960_/Y VGND VGND VPWR VPWR _8196_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_132_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7147_ _6920_/Y _7040_/D _6793_/Y _7110_/X _7146_/X VGND VGND VPWR VPWR _7154_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_86_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7078_ _7078_/A _7078_/B _7078_/C _7078_/D VGND VGND VPWR VPWR _7079_/D sky130_fd_sc_hd__and4_1
XFILLER_58_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6029_ _6029_/A VGND VGND VPWR VPWR _6029_/Y sky130_fd_sc_hd__inv_2
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9719_ _9770_/CLK _9719_/D _7011_/B VGND VGND VPWR VPWR _9719_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_42_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6380_ _9298_/Q VGND VGND VPWR VPWR _7216_/A sky130_fd_sc_hd__inv_4
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5400_ _9445_/Q _5395_/A _5964_/B1 _5395_/Y VGND VGND VPWR VPWR _9445_/D sky130_fd_sc_hd__a22o_1
XFILLER_173_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5331_ _9493_/Q _5330_/A _5963_/B1 _5330_/Y VGND VGND VPWR VPWR _9493_/D sky130_fd_sc_hd__a22o_1
XFILLER_154_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8050_ _8096_/B _8050_/B VGND VGND VPWR VPWR _8051_/A sky130_fd_sc_hd__or2_1
X_7001_ _9065_/Q _7001_/B VGND VGND VPWR VPWR _7002_/A sky130_fd_sc_hd__or2_1
X_5262_ _9540_/Q _5261_/A _5963_/B1 _5261_/Y VGND VGND VPWR VPWR _9540_/D sky130_fd_sc_hd__a22o_1
X_5193_ _5193_/A VGND VGND VPWR VPWR _5193_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8952_ _9711_/Q _6946_/Y _8957_/S VGND VGND VPWR VPWR _8952_/X sky130_fd_sc_hd__mux2_1
X_7903_ _8583_/A _8189_/A _7903_/C _8193_/A VGND VGND VPWR VPWR _7904_/A sky130_fd_sc_hd__or4_1
X_8883_ _8882_/X _9142_/Q _9054_/Q VGND VGND VPWR VPWR _8883_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7834_ _8226_/C VGND VGND VPWR VPWR _8496_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_70_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7765_ _7894_/B VGND VGND VPWR VPWR _8189_/A sky130_fd_sc_hd__inv_6
XFILLER_169_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4977_ _4994_/A VGND VGND VPWR VPWR _4978_/A sky130_fd_sc_hd__clkbuf_1
X_9504_ _9508_/CLK _9504_/D _9528_/SET_B VGND VGND VPWR VPWR _9504_/Q sky130_fd_sc_hd__dfrtp_1
X_6716_ _6716_/A _6716_/B _6716_/C _6716_/D VGND VGND VPWR VPWR _6784_/A sky130_fd_sc_hd__and4_1
XFILLER_149_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7696_ _6441_/Y _7471_/X _7392_/A _7473_/X _7695_/X VGND VGND VPWR VPWR _7697_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_177_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6647_ _6645_/Y _5742_/B _6646_/Y _5810_/B VGND VGND VPWR VPWR _6647_/X sky130_fd_sc_hd__o22a_1
X_9435_ _9440_/CLK _9435_/D _4628_/A VGND VGND VPWR VPWR _9435_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_166_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9366_ _9508_/CLK _9366_/D _9647_/SET_B VGND VGND VPWR VPWR _9366_/Q sky130_fd_sc_hd__dfrtp_1
X_6578_ _8779_/A _5267_/B _6577_/Y _5412_/B VGND VGND VPWR VPWR _6578_/X sky130_fd_sc_hd__o22a_1
XFILLER_192_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5529_ _9358_/Q _5528_/A _8843_/X _5528_/Y VGND VGND VPWR VPWR _9358_/D sky130_fd_sc_hd__a22o_1
XFILLER_117_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8317_ _8317_/A _8317_/B VGND VGND VPWR VPWR _8597_/C sky130_fd_sc_hd__or2_1
X_9297_ _9788_/CLK _9297_/D _9295_/SET_B VGND VGND VPWR VPWR _9297_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_117_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8248_ _8248_/A _8490_/B _8317_/B VGND VGND VPWR VPWR _8251_/A sky130_fd_sc_hd__or3_1
X_8179_ _8379_/B _8431_/A _8178_/X VGND VGND VPWR VPWR _8179_/X sky130_fd_sc_hd__a21o_1
XFILLER_132_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5880_ _9153_/Q _5874_/A _8955_/A1 _5874_/Y VGND VGND VPWR VPWR _9153_/D sky130_fd_sc_hd__a22o_1
X_4900_ _4931_/B _4900_/B VGND VGND VPWR VPWR _5404_/B sky130_fd_sc_hd__or2_4
XFILLER_65_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4831_ _4831_/A VGND VGND VPWR VPWR _4831_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_191 _6677_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_180 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7550_ _6457_/Y _7461_/X _6349_/Y _7463_/X _7549_/X VGND VGND VPWR VPWR _7553_/C
+ sky130_fd_sc_hd__o221a_1
X_4762_ _4891_/A _4843_/B VGND VGND VPWR VPWR _5829_/B sky130_fd_sc_hd__or2_4
X_4693_ _4685_/Y _5810_/B _4687_/Y _5949_/B _4692_/X VGND VGND VPWR VPWR _4705_/C
+ sky130_fd_sc_hd__o221a_1
X_7481_ _7481_/A _7481_/B _7481_/C _7481_/D VGND VGND VPWR VPWR _7482_/A sky130_fd_sc_hd__and4_2
X_6501_ _6501_/A _6501_/B _6501_/C _6501_/D VGND VGND VPWR VPWR _6629_/A sky130_fd_sc_hd__and4_1
XFILLER_146_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6432_ _6427_/Y _5317_/B _6428_/Y _5431_/B _6431_/X VGND VGND VPWR VPWR _6433_/D
+ sky130_fd_sc_hd__o221a_1
X_9220_ _9695_/CLK _9220_/D _9779_/SET_B VGND VGND VPWR VPWR _9220_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9151_ _9378_/CLK _9151_/D _9646_/SET_B VGND VGND VPWR VPWR _9151_/Q sky130_fd_sc_hd__dfstp_1
X_8102_ _8195_/A _8102_/B VGND VGND VPWR VPWR _8103_/A sky130_fd_sc_hd__or2_1
XFILLER_161_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6363_ _9337_/Q VGND VGND VPWR VPWR _6363_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5314_ _9504_/Q _5308_/A _8955_/A1 _5308_/Y VGND VGND VPWR VPWR _9504_/D sky130_fd_sc_hd__a22o_1
X_9082_ _9709_/CLK _9082_/D _6016_/X VGND VGND VPWR VPWR _9082_/Q sky130_fd_sc_hd__dfrtp_2
X_6294_ _6289_/Y _4564_/B _6290_/Y _5344_/B _6293_/X VGND VGND VPWR VPWR _6294_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_130_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8033_ _8033_/A _8614_/B VGND VGND VPWR VPWR _8035_/A sky130_fd_sc_hd__nor2_1
X_5245_ _9551_/Q _5242_/A _8844_/X _5242_/Y VGND VGND VPWR VPWR _9551_/D sky130_fd_sc_hd__a22o_1
XFILLER_114_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5176_ _9595_/Q _5169_/A _8840_/X _5169_/Y VGND VGND VPWR VPWR _9595_/D sky130_fd_sc_hd__a22o_1
XFILLER_152_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8935_ _9086_/Q _9085_/Q _9051_/Q VGND VGND VPWR VPWR _8935_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_5_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A VGND VGND VPWR VPWR _9039_/CLK sky130_fd_sc_hd__clkbuf_2
X_8866_ _7644_/Y _9628_/Q _8978_/S VGND VGND VPWR VPWR _8866_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8797_ _8797_/A VGND VGND VPWR VPWR _8798_/A sky130_fd_sc_hd__clkbuf_1
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7817_ _8341_/A VGND VGND VPWR VPWR _7836_/C sky130_fd_sc_hd__inv_2
XFILLER_51_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7748_ _9066_/Q _7748_/B VGND VGND VPWR VPWR _7748_/X sky130_fd_sc_hd__and2_1
XFILLER_101_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7679_ _7679_/A _7679_/B _7679_/C _7679_/D VGND VGND VPWR VPWR _7680_/D sky130_fd_sc_hd__and4_2
X_9418_ _9687_/CLK _9418_/D _9685_/SET_B VGND VGND VPWR VPWR _9418_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_152_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9349_ _9613_/CLK _9349_/D _9646_/SET_B VGND VGND VPWR VPWR _9349_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5030_ _9684_/Q _5026_/A _8840_/X _5026_/Y VGND VGND VPWR VPWR _9684_/D sky130_fd_sc_hd__a22o_1
XFILLER_97_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6981_ _6629_/Y _6976_/A _9015_/Q _6976_/Y VGND VGND VPWR VPWR _9015_/D sky130_fd_sc_hd__o22a_1
XFILLER_93_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5932_ _7832_/A VGND VGND VPWR VPWR _7837_/A sky130_fd_sc_hd__inv_2
X_8720_ _8720_/A _8720_/B _8720_/C VGND VGND VPWR VPWR _8721_/D sky130_fd_sc_hd__or3_1
XFILLER_18_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8651_ _8651_/A _8651_/B VGND VGND VPWR VPWR _8681_/C sky130_fd_sc_hd__or2_1
X_5863_ _8924_/X _6997_/A _5862_/Y _5849_/A _9164_/Q VGND VGND VPWR VPWR _9164_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_178_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4814_ _9070_/Q VGND VGND VPWR VPWR _4814_/Y sky130_fd_sc_hd__inv_6
X_8582_ _8582_/A _8582_/B VGND VGND VPWR VPWR _8646_/B sky130_fd_sc_hd__or2_1
X_7602_ _6140_/Y _7451_/X _6113_/Y _7453_/X _7601_/X VGND VGND VPWR VPWR _7607_/B
+ sky130_fd_sc_hd__o221a_1
X_5794_ _9214_/Q _5791_/A _5965_/B1 _5791_/Y VGND VGND VPWR VPWR _9214_/D sky130_fd_sc_hd__a22o_1
XFILLER_178_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7533_ _8783_/A _7475_/X _8759_/A _7477_/X VGND VGND VPWR VPWR _7533_/X sky130_fd_sc_hd__o22a_1
X_4745_ _4787_/A _4805_/A VGND VGND VPWR VPWR _6081_/B sky130_fd_sc_hd__or2_4
XFILLER_119_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7464_ _7476_/A _9251_/Q _7474_/C _9255_/Q VGND VGND VPWR VPWR _7465_/A sky130_fd_sc_hd__or4_1
X_4676_ _4787_/A _6158_/B VGND VGND VPWR VPWR _5507_/B sky130_fd_sc_hd__or2_4
X_6415_ _9454_/Q VGND VGND VPWR VPWR _6415_/Y sky130_fd_sc_hd__clkinv_4
X_9203_ _9203_/CLK _9203_/D _9633_/SET_B VGND VGND VPWR VPWR _9203_/Q sky130_fd_sc_hd__dfrtp_1
X_7395_ _6404_/Y _7124_/X _6343_/Y _7068_/B _7394_/X VGND VGND VPWR VPWR _7396_/D
+ sky130_fd_sc_hd__o221a_1
X_9134_ _9358_/CLK _9134_/D _9685_/SET_B VGND VGND VPWR VPWR _9134_/Q sky130_fd_sc_hd__dfrtp_1
X_6346_ _9532_/Q VGND VGND VPWR VPWR _6346_/Y sky130_fd_sc_hd__inv_2
X_9065_ _9664_/CLK _9065_/D _6146_/A VGND VGND VPWR VPWR _9065_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_130_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8016_ _8016_/A _8016_/B _8016_/C _8016_/D VGND VGND VPWR VPWR _8016_/X sky130_fd_sc_hd__or4_1
X_6277_ _9351_/Q VGND VGND VPWR VPWR _6277_/Y sky130_fd_sc_hd__inv_2
Xinput118 sram_ro_data[3] VGND VGND VPWR VPWR _6564_/A sky130_fd_sc_hd__clkbuf_1
Xinput107 sram_ro_data[22] VGND VGND VPWR VPWR _6219_/A sky130_fd_sc_hd__clkbuf_1
Xinput129 usr1_vdd_pwrgood VGND VGND VPWR VPWR _6847_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_102_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5228_ _5966_/B1 _9560_/Q _5230_/S VGND VGND VPWR VPWR _5229_/A sky130_fd_sc_hd__mux2_1
X_5159_ _9609_/Q _5158_/A _8846_/X _5158_/Y VGND VGND VPWR VPWR _9609_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8918_ _9608_/Q _8845_/X _8926_/S VGND VGND VPWR VPWR _8918_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8849_ _9618_/Q _8916_/A1 _8955_/S VGND VGND VPWR VPWR _8849_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_2_1_0_csclk clkbuf_2_1_0_csclk/A VGND VGND VPWR VPWR clkbuf_2_1_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_2
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_91 input77/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_80 _8824_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4530_ _9766_/Q _4526_/A _5963_/B1 _4526_/Y VGND VGND VPWR VPWR _9766_/D sky130_fd_sc_hd__a22o_1
XFILLER_116_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4461_ _8944_/X VGND VGND VPWR VPWR _4729_/B sky130_fd_sc_hd__clkinv_2
X_7180_ _8789_/A _7082_/X _8791_/A _7084_/X _7179_/X VGND VGND VPWR VPWR _7199_/A
+ sky130_fd_sc_hd__o221a_2
X_6200_ _9448_/Q VGND VGND VPWR VPWR _6200_/Y sky130_fd_sc_hd__inv_2
X_6131_ _6126_/Y _5776_/B _6127_/Y _5949_/B _6130_/X VGND VGND VPWR VPWR _6144_/B
+ sky130_fd_sc_hd__o221a_1
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6062_ _9653_/Q VGND VGND VPWR VPWR _6062_/Y sky130_fd_sc_hd__inv_2
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ _5960_/A _5013_/B VGND VGND VPWR VPWR _5014_/A sky130_fd_sc_hd__or2_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6964_ _6964_/A VGND VGND VPWR VPWR _6964_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9752_ _9755_/CLK _9752_/D _9757_/SET_B VGND VGND VPWR VPWR _9752_/Q sky130_fd_sc_hd__dfstp_1
X_9683_ _9684_/CLK _9683_/D _9685_/SET_B VGND VGND VPWR VPWR _9683_/Q sky130_fd_sc_hd__dfrtp_1
X_8703_ _8703_/A _8703_/B _8703_/C _8703_/D VGND VGND VPWR VPWR _8706_/C sky130_fd_sc_hd__or4_1
X_6895_ _9321_/Q VGND VGND VPWR VPWR _6895_/Y sky130_fd_sc_hd__clkinv_2
X_5915_ _9125_/Q _5907_/A _8916_/A1 _5907_/Y VGND VGND VPWR VPWR _9125_/D sky130_fd_sc_hd__a22o_1
XFILLER_81_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8634_ _8544_/A _8092_/Y _8587_/A _8431_/A VGND VGND VPWR VPWR _8714_/A sky130_fd_sc_hd__a211o_1
X_5846_ _9178_/Q _5839_/A _8930_/A1 _5839_/Y VGND VGND VPWR VPWR _9178_/D sky130_fd_sc_hd__a22o_1
XFILLER_166_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8565_ _8565_/A _8640_/B VGND VGND VPWR VPWR _8720_/B sky130_fd_sc_hd__nor2_1
XFILLER_166_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5777_ _5777_/A VGND VGND VPWR VPWR _5778_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_181_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8496_ _8496_/A _8496_/B VGND VGND VPWR VPWR _8695_/C sky130_fd_sc_hd__nor2_2
X_4728_ _9240_/Q VGND VGND VPWR VPWR _4731_/A sky130_fd_sc_hd__inv_2
X_7516_ _6755_/Y _7471_/X _7172_/A _7473_/X _7515_/X VGND VGND VPWR VPWR _7517_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_174_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7447_ _7447_/A VGND VGND VPWR VPWR _7447_/X sky130_fd_sc_hd__buf_8
X_4659_ _7003_/C VGND VGND VPWR VPWR _8957_/S sky130_fd_sc_hd__clkinv_4
XFILLER_162_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7378_ _6397_/Y _7082_/X _6387_/Y _7084_/X _7377_/X VGND VGND VPWR VPWR _7397_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_1_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6329_ _9506_/Q VGND VGND VPWR VPWR _6329_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_143_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9117_ _9785_/CLK _9117_/D _9779_/SET_B VGND VGND VPWR VPWR _9117_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9048_ _9709_/CLK _9048_/D _6051_/X VGND VGND VPWR VPWR _9048_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_190_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_32_csclk clkbuf_opt_3_0_csclk/X VGND VGND VPWR VPWR _9695_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_79_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_47_csclk _9329_/CLK VGND VGND VPWR VPWR _9776_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_57_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5700_ _9255_/Q _5692_/Y _5696_/Y _5724_/B _5699_/X VGND VGND VPWR VPWR _9255_/D
+ sky130_fd_sc_hd__o32a_1
X_6680_ _6680_/A VGND VGND VPWR VPWR _6680_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_188_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5631_ _9286_/Q _5623_/A _8916_/A1 _5623_/Y VGND VGND VPWR VPWR _9286_/D sky130_fd_sc_hd__a22o_1
X_8350_ _8583_/A _8583_/B _8350_/C VGND VGND VPWR VPWR _8640_/C sky130_fd_sc_hd__or3_4
XFILLER_148_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5562_ _9334_/Q _5558_/A _8930_/A1 _5558_/Y VGND VGND VPWR VPWR _9334_/D sky130_fd_sc_hd__a22o_1
X_8281_ _8678_/A _8281_/B VGND VGND VPWR VPWR _8283_/A sky130_fd_sc_hd__or2_1
XFILLER_129_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7301_ _4694_/Y _7040_/D _4660_/Y _7110_/X _7300_/X VGND VGND VPWR VPWR _7308_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_117_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4513_ _4669_/A _8932_/X _4729_/A _8944_/X VGND VGND VPWR VPWR _4898_/A sky130_fd_sc_hd__or4_4
X_7232_ _6288_/Y _7048_/D _6314_/Y _7040_/B _7231_/X VGND VGND VPWR VPWR _7233_/D
+ sky130_fd_sc_hd__o221a_1
X_5493_ _9382_/Q _5490_/A _5965_/B1 _5490_/Y VGND VGND VPWR VPWR _9382_/D sky130_fd_sc_hd__a22o_1
X_4444_ _9589_/Q input78/X _8833_/S VGND VGND VPWR VPWR _9010_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7163_ _6720_/Y _7079_/B _6633_/Y _7059_/A VGND VGND VPWR VPWR _7163_/X sky130_fd_sc_hd__o22a_1
X_6114_ _9475_/Q VGND VGND VPWR VPWR _6114_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_112_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7094_ _7127_/C _7094_/B VGND VGND VPWR VPWR _7095_/A sky130_fd_sc_hd__or2_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6045_ _6045_/A VGND VGND VPWR VPWR _6045_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_58_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7996_ _7996_/A VGND VGND VPWR VPWR _8130_/B sky130_fd_sc_hd__clkbuf_4
X_9735_ _9774_/CLK _9735_/D _9757_/SET_B VGND VGND VPWR VPWR _9735_/Q sky130_fd_sc_hd__dfstp_1
X_6947_ _6149_/A _6946_/Y _9037_/Q _6149_/Y VGND VGND VPWR VPWR _9037_/D sky130_fd_sc_hd__o22a_1
XFILLER_81_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9666_ _4450_/A1 _9666_/D _6146_/A VGND VGND VPWR VPWR _9666_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_149_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6878_ _6878_/A _6878_/B _6878_/C _6878_/D VGND VGND VPWR VPWR _6946_/B sky130_fd_sc_hd__and4_1
X_9597_ _9601_/CLK _9597_/D _9528_/SET_B VGND VGND VPWR VPWR _9597_/Q sky130_fd_sc_hd__dfrtp_1
X_8617_ _8617_/A _8617_/B VGND VGND VPWR VPWR _8707_/A sky130_fd_sc_hd__or2_1
X_5829_ _5960_/A _5829_/B VGND VGND VPWR VPWR _5830_/A sky130_fd_sc_hd__or2_1
X_8548_ _8393_/Y _8554_/B _8401_/A _8554_/B _8547_/X VGND VGND VPWR VPWR _8548_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_5_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8479_ _8704_/B _8479_/B VGND VGND VPWR VPWR _8481_/A sky130_fd_sc_hd__or2_1
XFILLER_190_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput208 _8831_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[0] sky130_fd_sc_hd__buf_2
XFILLER_126_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput219 _8832_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[1] sky130_fd_sc_hd__buf_2
XFILLER_181_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7850_ _7850_/A VGND VGND VPWR VPWR _8521_/B sky130_fd_sc_hd__buf_12
XFILLER_36_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6801_ _9360_/Q VGND VGND VPWR VPWR _6801_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7781_ _7781_/A _7781_/B VGND VGND VPWR VPWR _7781_/Y sky130_fd_sc_hd__nand2_1
XFILLER_63_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4993_ _4993_/A VGND VGND VPWR VPWR _9700_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9520_ _9527_/CLK _9520_/D _9528_/SET_B VGND VGND VPWR VPWR _9520_/Q sky130_fd_sc_hd__dfstp_1
X_6732_ _9656_/Q VGND VGND VPWR VPWR _6732_/Y sky130_fd_sc_hd__inv_2
X_9451_ _9483_/CLK _9451_/D _9685_/SET_B VGND VGND VPWR VPWR _9451_/Q sky130_fd_sc_hd__dfstp_1
X_6663_ _9283_/Q VGND VGND VPWR VPWR _7348_/A sky130_fd_sc_hd__inv_2
XFILLER_139_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5614_ _9300_/Q _5612_/A _8845_/X _5612_/Y VGND VGND VPWR VPWR _9300_/D sky130_fd_sc_hd__a22o_1
X_8402_ _8213_/A _8117_/A _8019_/C _8400_/X _8401_/X VGND VGND VPWR VPWR _8402_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_31_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6594_ _9419_/Q VGND VGND VPWR VPWR _8795_/A sky130_fd_sc_hd__inv_6
XFILLER_176_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9382_ _9771_/CLK _9382_/D _4628_/A VGND VGND VPWR VPWR _9382_/Q sky130_fd_sc_hd__dfstp_1
X_5545_ _5545_/A _5545_/B VGND VGND VPWR VPWR _5546_/A sky130_fd_sc_hd__or2_1
X_8333_ _8720_/A _8713_/A _8333_/C VGND VGND VPWR VPWR _8335_/A sky130_fd_sc_hd__or3_1
X_5476_ _9393_/Q _5471_/A _8842_/X _5471_/Y VGND VGND VPWR VPWR _9393_/D sky130_fd_sc_hd__a22o_1
X_8264_ _8324_/A _8264_/B VGND VGND VPWR VPWR _8645_/B sky130_fd_sc_hd__nor2_1
X_8195_ _8195_/A _8195_/B VGND VGND VPWR VPWR _8195_/Y sky130_fd_sc_hd__nor2_1
XFILLER_144_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7215_ _6456_/Y _7059_/D _6421_/Y _7116_/X _7214_/X VGND VGND VPWR VPWR _7220_/B
+ sky130_fd_sc_hd__o221a_1
X_7146_ _6895_/Y _7112_/X _6889_/Y _7077_/B VGND VGND VPWR VPWR _7146_/X sky130_fd_sc_hd__o22a_1
XFILLER_59_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7077_ _7077_/A _7077_/B _7077_/C _7077_/D VGND VGND VPWR VPWR _7078_/D sky130_fd_sc_hd__and4_1
X_6028_ _6028_/A VGND VGND VPWR VPWR _6029_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_100_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7979_ _7979_/A VGND VGND VPWR VPWR _7994_/A sky130_fd_sc_hd__inv_2
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9718_ _8837_/A1 _9718_/D _4994_/A VGND VGND VPWR VPWR _9718_/Q sky130_fd_sc_hd__dfrtn_1
X_9649_ _9652_/CLK _9649_/D _9646_/SET_B VGND VGND VPWR VPWR _9649_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5330_ _5330_/A VGND VGND VPWR VPWR _5330_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5261_ _5261_/A VGND VGND VPWR VPWR _5261_/Y sky130_fd_sc_hd__inv_2
X_7000_ _9056_/Q _5753_/B _6996_/Y _6999_/Y VGND VGND VPWR VPWR _9056_/D sky130_fd_sc_hd__a22o_1
X_5192_ _6322_/A _6165_/A _5259_/A _8956_/X VGND VGND VPWR VPWR _5193_/A sky130_fd_sc_hd__a211o_4
XFILLER_68_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8951_ _9712_/Q _6785_/Y _8957_/S VGND VGND VPWR VPWR _8951_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7902_ _8077_/A _7902_/B VGND VGND VPWR VPWR _7902_/X sky130_fd_sc_hd__or2_1
XFILLER_110_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8882_ _7243_/Y _9637_/Q _8959_/S VGND VGND VPWR VPWR _8882_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7833_ _7833_/A VGND VGND VPWR VPWR _8226_/C sky130_fd_sc_hd__buf_8
X_7764_ _7764_/A VGND VGND VPWR VPWR _8510_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_24_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4976_ _9704_/Q _4966_/A _9703_/Q _4966_/Y VGND VGND VPWR VPWR _9704_/D sky130_fd_sc_hd__a22o_1
X_9503_ _9527_/CLK _9503_/D _9528_/SET_B VGND VGND VPWR VPWR _9503_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_149_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6715_ _6710_/Y _5420_/B _6711_/Y _5259_/B _6714_/X VGND VGND VPWR VPWR _6716_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_51_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7695_ _6429_/Y _7475_/X _6379_/Y _7477_/X VGND VGND VPWR VPWR _7695_/X sky130_fd_sc_hd__o22a_1
XFILLER_192_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6646_ _9200_/Q VGND VGND VPWR VPWR _6646_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9434_ _9440_/CLK _9434_/D _4628_/A VGND VGND VPWR VPWR _9434_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_192_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9365_ _9508_/CLK _9365_/D _9647_/SET_B VGND VGND VPWR VPWR _9365_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_137_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6577_ _9435_/Q VGND VGND VPWR VPWR _6577_/Y sky130_fd_sc_hd__inv_2
X_5528_ _5528_/A VGND VGND VPWR VPWR _5528_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8316_ _8316_/A _8498_/B VGND VGND VPWR VPWR _8490_/C sky130_fd_sc_hd__nor2_1
XFILLER_3_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9296_ _9788_/CLK _9296_/D _9295_/SET_B VGND VGND VPWR VPWR _9296_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_132_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8247_ _8319_/A _8264_/B VGND VGND VPWR VPWR _8317_/B sky130_fd_sc_hd__nor2_1
X_5459_ _5459_/A VGND VGND VPWR VPWR _5460_/A sky130_fd_sc_hd__clkbuf_4
X_8178_ _8703_/A _8178_/B VGND VGND VPWR VPWR _8178_/X sky130_fd_sc_hd__or2_1
XFILLER_113_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7129_ _4814_/Y _7126_/X _4857_/Y _7128_/X VGND VGND VPWR VPWR _7129_/X sky130_fd_sc_hd__o22a_1
XFILLER_115_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_170 _7021_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4830_ _4830_/A _4830_/B _4830_/C _4830_/D VGND VGND VPWR VPWR _4935_/A sky130_fd_sc_hd__and4_1
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_181 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_192 _8765_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4761_ _9185_/Q VGND VGND VPWR VPWR _4761_/Y sky130_fd_sc_hd__inv_2
X_7480_ _7480_/A _7480_/B _7480_/C _7480_/D VGND VGND VPWR VPWR _7481_/D sky130_fd_sc_hd__and4_1
X_4692_ _4692_/A _5024_/B VGND VGND VPWR VPWR _4692_/X sky130_fd_sc_hd__or2_1
X_6500_ _7370_/A _5632_/B _7701_/A _5905_/B _6499_/X VGND VGND VPWR VPWR _6501_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_174_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6431_ _6429_/Y _4504_/B _6430_/Y _6027_/B VGND VGND VPWR VPWR _6431_/X sky130_fd_sc_hd__o22a_1
X_6362_ _9244_/Q VGND VGND VPWR VPWR _6362_/Y sky130_fd_sc_hd__inv_2
X_9150_ _9279_/CLK _9150_/D _9757_/SET_B VGND VGND VPWR VPWR _9150_/Q sky130_fd_sc_hd__dfrtp_1
X_5313_ _9505_/Q _5308_/A _8842_/X _5308_/Y VGND VGND VPWR VPWR _9505_/D sky130_fd_sc_hd__a22o_1
X_8101_ _8213_/A VGND VGND VPWR VPWR _8625_/A sky130_fd_sc_hd__clkinv_2
X_9081_ _9788_/CLK _9081_/D _9646_/SET_B VGND VGND VPWR VPWR _9081_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_88_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6293_ _6291_/Y _6027_/B _6292_/Y _4893_/X VGND VGND VPWR VPWR _6293_/X sky130_fd_sc_hd__o22a_1
XFILLER_114_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8032_ _8521_/A _8551_/A VGND VGND VPWR VPWR _8614_/B sky130_fd_sc_hd__nor2_1
X_5244_ _9552_/Q _5242_/A _8845_/X _5242_/Y VGND VGND VPWR VPWR _9552_/D sky130_fd_sc_hd__a22o_1
X_5175_ _9596_/Q _5169_/A _8841_/X _5169_/Y VGND VGND VPWR VPWR _9596_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8934_ _8933_/X _9678_/Q _9587_/Q VGND VGND VPWR VPWR _8934_/X sky130_fd_sc_hd__mux2_4
XFILLER_56_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8865_ _8864_/X _9171_/Q _9054_/Q VGND VGND VPWR VPWR _8865_/X sky130_fd_sc_hd__mux2_1
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7816_ _8202_/A _8097_/B VGND VGND VPWR VPWR _8094_/A sky130_fd_sc_hd__or2_1
XFILLER_24_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8796_ _8796_/A VGND VGND VPWR VPWR _8796_/X sky130_fd_sc_hd__clkbuf_1
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7747_ _9068_/Q _7747_/A2 _9067_/Q _7747_/B2 _7746_/X VGND VGND VPWR VPWR _7747_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_24_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4959_ _9048_/Q VGND VGND VPWR VPWR _6022_/B sky130_fd_sc_hd__clkinv_4
XFILLER_177_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7678_ _6528_/Y _7471_/X _7370_/A _7473_/X _7677_/X VGND VGND VPWR VPWR _7679_/D
+ sky130_fd_sc_hd__o221a_1
X_9417_ _9684_/CLK _9417_/D _9685_/SET_B VGND VGND VPWR VPWR _9417_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_177_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6629_ _6629_/A _6629_/B _6629_/C _6629_/D VGND VGND VPWR VPWR _6629_/Y sky130_fd_sc_hd__nand4_4
XFILLER_152_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9348_ _9352_/CLK _9348_/D _9646_/SET_B VGND VGND VPWR VPWR _9348_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9279_ _9279_/CLK _9279_/D _9633_/SET_B VGND VGND VPWR VPWR _9279_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6980_ _6475_/Y _6976_/A _9016_/Q _6976_/Y VGND VGND VPWR VPWR _9016_/D sky130_fd_sc_hd__o22a_2
X_5931_ _5931_/A _5931_/B input164/X input202/X VGND VGND VPWR VPWR _5935_/C sky130_fd_sc_hd__or4bb_1
XFILLER_80_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8650_ _8672_/C _8650_/B _8650_/C VGND VGND VPWR VPWR _8722_/B sky130_fd_sc_hd__or3_1
X_5862_ _8978_/X VGND VGND VPWR VPWR _5862_/Y sky130_fd_sc_hd__inv_2
X_8581_ _8005_/A _8279_/C _8280_/B VGND VGND VPWR VPWR _8582_/B sky130_fd_sc_hd__o21ai_1
X_7601_ _6098_/Y _7455_/X _6062_/Y _7457_/X VGND VGND VPWR VPWR _7601_/X sky130_fd_sc_hd__o22a_1
XFILLER_21_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4813_ _9761_/Q VGND VGND VPWR VPWR _4813_/Y sky130_fd_sc_hd__inv_2
X_5793_ _9215_/Q _5791_/A _5964_/B1 _5791_/Y VGND VGND VPWR VPWR _9215_/D sky130_fd_sc_hd__a22o_1
XFILLER_193_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4744_ _9390_/Q VGND VGND VPWR VPWR _4744_/Y sky130_fd_sc_hd__inv_2
X_7532_ _8747_/A _7461_/X _8787_/A _7463_/X _7531_/X VGND VGND VPWR VPWR _7535_/C
+ sky130_fd_sc_hd__o221a_1
X_4675_ _9364_/Q VGND VGND VPWR VPWR _4675_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_119_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9202_ _9440_/CLK _9202_/D _4628_/A VGND VGND VPWR VPWR _9202_/Q sky130_fd_sc_hd__dfrtp_1
X_7463_ _7463_/A VGND VGND VPWR VPWR _7463_/X sky130_fd_sc_hd__buf_8
X_6414_ _6409_/Y _5442_/B _6410_/Y _5583_/B _6413_/X VGND VGND VPWR VPWR _6433_/A
+ sky130_fd_sc_hd__o221a_1
X_7394_ _6429_/Y _7126_/X _6341_/Y _7128_/X VGND VGND VPWR VPWR _7394_/X sky130_fd_sc_hd__o22a_1
X_9133_ _9354_/CLK _9133_/D _9685_/SET_B VGND VGND VPWR VPWR _9133_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_127_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6345_ _6340_/Y _5259_/B _6341_/Y _5251_/B _6344_/X VGND VGND VPWR VPWR _6352_/C
+ sky130_fd_sc_hd__o221a_1
X_9064_ _4450_/A1 _9064_/D _6146_/A VGND VGND VPWR VPWR _9064_/Q sky130_fd_sc_hd__dfrtp_1
X_6276_ _9377_/Q VGND VGND VPWR VPWR _6276_/Y sky130_fd_sc_hd__inv_2
X_8015_ _7902_/B _8013_/B _8093_/A VGND VGND VPWR VPWR _8016_/D sky130_fd_sc_hd__a21oi_1
XFILLER_102_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5227_ _5259_/A _5227_/B VGND VGND VPWR VPWR _5230_/S sky130_fd_sc_hd__or2_1
Xinput108 sram_ro_data[23] VGND VGND VPWR VPWR _6100_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_102_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput119 sram_ro_data[4] VGND VGND VPWR VPWR _6451_/A sky130_fd_sc_hd__clkbuf_1
X_5158_ _5158_/A VGND VGND VPWR VPWR _5158_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5089_ _5545_/A _5089_/B VGND VGND VPWR VPWR _5090_/A sky130_fd_sc_hd__or2_1
X_8917_ _9609_/Q _8846_/X _8926_/S VGND VGND VPWR VPWR _8917_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8848_ _9602_/Q _8916_/A1 _8926_/S VGND VGND VPWR VPWR _8848_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8779_ _8779_/A VGND VGND VPWR VPWR _8780_/A sky130_fd_sc_hd__clkbuf_1
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_92 input77/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_70 _7482_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_81 _8822_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4460_ _8946_/X VGND VGND VPWR VPWR _4729_/A sky130_fd_sc_hd__clkinv_2
XFILLER_116_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6130_ _6128_/Y _5872_/B _6129_/Y _5045_/B VGND VGND VPWR VPWR _6130_/X sky130_fd_sc_hd__o22a_1
XFILLER_112_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ _9319_/Q VGND VGND VPWR VPWR _6061_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ _9048_/Q _8957_/S _4949_/A _9696_/Q _5011_/X VGND VGND VPWR VPWR _9696_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_38_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6963_ _6963_/A VGND VGND VPWR VPWR _6964_/A sky130_fd_sc_hd__clkbuf_4
X_9751_ _9755_/CLK _9751_/D _9757_/SET_B VGND VGND VPWR VPWR _9751_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_38_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8702_ _8732_/A _8735_/C VGND VGND VPWR VPWR _8702_/Y sky130_fd_sc_hd__nor2_1
X_6894_ _6889_/Y _5872_/B _6890_/Y _5776_/B _6893_/X VGND VGND VPWR VPWR _6901_/C
+ sky130_fd_sc_hd__o221a_1
X_5914_ _9126_/Q _5907_/A _8930_/A1 _5907_/Y VGND VGND VPWR VPWR _9126_/D sky130_fd_sc_hd__a22o_1
X_9682_ _9709_/CLK _9682_/D _5033_/X VGND VGND VPWR VPWR _9682_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5845_ _9179_/Q _5839_/A _8955_/A1 _5839_/Y VGND VGND VPWR VPWR _9179_/D sky130_fd_sc_hd__a22o_1
X_8633_ _8633_/A _8709_/C _8688_/C _8687_/C VGND VGND VPWR VPWR _8633_/Y sky130_fd_sc_hd__nor4_1
XFILLER_167_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8564_ _8636_/A _8636_/B _8636_/C _8563_/X VGND VGND VPWR VPWR _8564_/X sky130_fd_sc_hd__or4b_1
X_5776_ _6052_/A _5776_/B VGND VGND VPWR VPWR _5777_/A sky130_fd_sc_hd__or2_1
XFILLER_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8495_ _8341_/A _8498_/A _8189_/A _7885_/X VGND VGND VPWR VPWR _8496_/B sky130_fd_sc_hd__o22a_1
XFILLER_135_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7515_ _6650_/Y _7475_/X _6633_/Y _7477_/X VGND VGND VPWR VPWR _7515_/X sky130_fd_sc_hd__o22a_1
X_4727_ _4898_/A _4780_/B VGND VGND VPWR VPWR _5660_/B sky130_fd_sc_hd__or2_4
X_7446_ _7456_/A _7472_/A _7474_/D VGND VGND VPWR VPWR _7447_/A sky130_fd_sc_hd__or3_1
X_4658_ _9091_/Q _9090_/Q _9092_/Q VGND VGND VPWR VPWR _7003_/C sky130_fd_sc_hd__or3_2
Xinput90 spimemio_flash_io2_oeb VGND VGND VPWR VPWR input90/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7377_ _6362_/Y _7077_/C _6440_/Y _7077_/D _7376_/X VGND VGND VPWR VPWR _7377_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_1_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4589_ _6158_/A _4903_/B VGND VGND VPWR VPWR _4590_/B sky130_fd_sc_hd__or2_4
X_9116_ _9779_/CLK _9116_/D _9779_/SET_B VGND VGND VPWR VPWR _9116_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_107_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6328_ _9402_/Q VGND VGND VPWR VPWR _6328_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_130_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9047_ _9790_/CLK _9047_/D VGND VGND VPWR VPWR _9047_/Q sky130_fd_sc_hd__dfxtp_1
X_6259_ input8/X VGND VGND VPWR VPWR _6259_/Y sky130_fd_sc_hd__inv_2
XFILLER_190_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5630_ _9287_/Q _5623_/A _8840_/X _5623_/Y VGND VGND VPWR VPWR _9287_/D sky130_fd_sc_hd__a22o_1
X_5561_ _9335_/Q _5558_/A _8841_/X _5558_/Y VGND VGND VPWR VPWR _9335_/D sky130_fd_sc_hd__a22o_1
X_8280_ _8275_/X _8280_/B _8280_/C VGND VGND VPWR VPWR _8281_/B sky130_fd_sc_hd__nand3b_1
X_7300_ _4718_/Y _7112_/X _4699_/Y _7077_/B VGND VGND VPWR VPWR _7300_/X sky130_fd_sc_hd__o22a_1
XFILLER_117_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5492_ _9383_/Q _5490_/A _5964_/B1 _5490_/Y VGND VGND VPWR VPWR _9383_/D sky130_fd_sc_hd__a22o_1
X_4512_ _9772_/Q _4466_/A _5963_/B1 _4466_/Y VGND VGND VPWR VPWR _9772_/D sky130_fd_sc_hd__a22o_1
XFILLER_156_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7231_ _6301_/Y _7068_/A _6263_/Y _7105_/X VGND VGND VPWR VPWR _7231_/X sky130_fd_sc_hd__o22a_1
XFILLER_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4443_ _9588_/Q input80/X _8833_/S VGND VGND VPWR VPWR _9009_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7162_ _6736_/Y _7095_/X _6643_/Y _7068_/D _7161_/X VGND VGND VPWR VPWR _7167_/B
+ sky130_fd_sc_hd__o221a_1
X_6113_ _9457_/Q VGND VGND VPWR VPWR _6113_/Y sky130_fd_sc_hd__inv_2
X_7093_ _4740_/Y _7048_/B _4701_/Y _7077_/A _7092_/X VGND VGND VPWR VPWR _7108_/A
+ sky130_fd_sc_hd__o221a_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6044_ _6050_/A VGND VGND VPWR VPWR _6045_/A sky130_fd_sc_hd__clkbuf_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7995_ _8116_/B _7995_/B VGND VGND VPWR VPWR _7996_/A sky130_fd_sc_hd__or2_1
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9734_ _9774_/CLK _9734_/D _9757_/SET_B VGND VGND VPWR VPWR _9734_/Q sky130_fd_sc_hd__dfstp_1
X_6946_ _6946_/A _6946_/B _6946_/C VGND VGND VPWR VPWR _6946_/Y sky130_fd_sc_hd__nand3_4
XFILLER_54_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9665_ _4450_/A1 _9665_/D _6146_/A VGND VGND VPWR VPWR _9665_/Q sky130_fd_sc_hd__dfrtp_1
X_6877_ _6877_/A _6877_/B _6877_/C _6877_/D VGND VGND VPWR VPWR _6878_/D sky130_fd_sc_hd__and4_1
X_9596_ _9596_/CLK _9596_/D _9528_/SET_B VGND VGND VPWR VPWR _9596_/Q sky130_fd_sc_hd__dfrtp_1
X_5828_ _9190_/Q _5820_/A _8916_/A1 _5820_/Y VGND VGND VPWR VPWR _9190_/D sky130_fd_sc_hd__a22o_1
X_8616_ _8735_/A _8616_/B _8668_/D _8699_/C VGND VGND VPWR VPWR _8619_/A sky130_fd_sc_hd__or4_2
XFILLER_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5759_ _5759_/A VGND VGND VPWR VPWR _5759_/Y sky130_fd_sc_hd__inv_2
X_8547_ _8098_/A _8546_/Y _8398_/Y VGND VGND VPWR VPWR _8547_/X sky130_fd_sc_hd__o21a_1
XFILLER_108_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8478_ _8703_/D _8478_/B VGND VGND VPWR VPWR _8479_/B sky130_fd_sc_hd__or2_1
XFILLER_162_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7429_ _7476_/A _9251_/Q _7470_/B _9255_/Q VGND VGND VPWR VPWR _7430_/A sky130_fd_sc_hd__or4_1
XFILLER_78_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput209 _8752_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[10] sky130_fd_sc_hd__buf_2
XFILLER_141_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6800_ _9115_/Q VGND VGND VPWR VPWR _6800_/Y sky130_fd_sc_hd__inv_2
X_7780_ _8218_/B VGND VGND VPWR VPWR _7969_/A sky130_fd_sc_hd__inv_2
X_4992_ _8909_/X _9700_/Q _5001_/S VGND VGND VPWR VPWR _4993_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6731_ _9103_/Q VGND VGND VPWR VPWR _6731_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_51_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9450_ _9483_/CLK _9450_/D _9528_/SET_B VGND VGND VPWR VPWR _9450_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_149_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6662_ _9335_/Q VGND VGND VPWR VPWR _6662_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_31_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5613_ _9301_/Q _5612_/A _8846_/X _5612_/Y VGND VGND VPWR VPWR _9301_/D sky130_fd_sc_hd__a22o_1
X_8401_ _8401_/A _8401_/B VGND VGND VPWR VPWR _8401_/X sky130_fd_sc_hd__or2_1
X_9381_ _9771_/CLK _9381_/D _4628_/A VGND VGND VPWR VPWR _9381_/Q sky130_fd_sc_hd__dfrtp_1
X_6593_ _6593_/A VGND VGND VPWR VPWR _6593_/Y sky130_fd_sc_hd__clkinv_2
X_8332_ _8299_/A _8282_/C _8282_/B _8331_/X VGND VGND VPWR VPWR _8333_/C sky130_fd_sc_hd__a31o_1
XFILLER_129_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5544_ _9346_/Q _5536_/A _8916_/A1 _5536_/Y VGND VGND VPWR VPWR _9346_/D sky130_fd_sc_hd__a22o_1
X_5475_ _9394_/Q _5471_/A _8925_/A1 _5471_/Y VGND VGND VPWR VPWR _9394_/D sky130_fd_sc_hd__a22o_1
XFILLER_144_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8263_ _8263_/A _8369_/B VGND VGND VPWR VPWR _8265_/A sky130_fd_sc_hd__or2_1
X_8194_ _8204_/A VGND VGND VPWR VPWR _8346_/B sky130_fd_sc_hd__inv_2
XFILLER_105_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7214_ _6346_/Y _7118_/X _6436_/Y _7048_/C VGND VGND VPWR VPWR _7214_/X sky130_fd_sc_hd__o22a_1
XFILLER_132_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7145_ _7145_/A _7145_/B _7145_/C _7145_/D VGND VGND VPWR VPWR _7155_/B sky130_fd_sc_hd__and4_1
XFILLER_113_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7076_ _7076_/A VGND VGND VPWR VPWR _7077_/D sky130_fd_sc_hd__buf_8
X_6027_ _6052_/A _6027_/B VGND VGND VPWR VPWR _6028_/A sky130_fd_sc_hd__or2_1
XFILLER_100_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7978_ _8096_/A _8098_/A VGND VGND VPWR VPWR _7995_/B sky130_fd_sc_hd__or2_1
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_31_csclk clkbuf_opt_2_0_csclk/X VGND VGND VPWR VPWR _9379_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_81_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6929_ _9102_/Q VGND VGND VPWR VPWR _6929_/Y sky130_fd_sc_hd__inv_2
X_9717_ _9709_/CLK hold2/X _4639_/X VGND VGND VPWR VPWR _9717_/Q sky130_fd_sc_hd__dfrtn_1
X_9648_ _9652_/CLK _9648_/D _9646_/SET_B VGND VGND VPWR VPWR _9648_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_80_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9579_ _9674_/CLK _9579_/D _9633_/SET_B VGND VGND VPWR VPWR _9579_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_129_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_46_csclk _9329_/CLK VGND VGND VPWR VPWR _9775_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_170_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_1_0_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_89_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5260_ _5260_/A VGND VGND VPWR VPWR _5261_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_141_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5191_ _9052_/Q _5985_/B _9586_/Q VGND VGND VPWR VPWR _9586_/D sky130_fd_sc_hd__a21o_1
XFILLER_83_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8950_ _9714_/Q _6475_/Y _8957_/S VGND VGND VPWR VPWR _8950_/X sky130_fd_sc_hd__mux2_1
X_7901_ _8472_/A _8517_/A VGND VGND VPWR VPWR _7902_/B sky130_fd_sc_hd__or2_1
XFILLER_55_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8881_ _8880_/X _9141_/Q _9054_/Q VGND VGND VPWR VPWR _8881_/X sky130_fd_sc_hd__mux2_1
X_7832_ _7832_/A _7837_/B _7837_/C VGND VGND VPWR VPWR _7833_/A sky130_fd_sc_hd__or3_1
X_4975_ _4975_/A VGND VGND VPWR VPWR _4975_/X sky130_fd_sc_hd__clkbuf_1
X_7763_ _8394_/A _8379_/B _7838_/B VGND VGND VPWR VPWR _7764_/A sky130_fd_sc_hd__or3_1
X_9502_ _9527_/CLK _9502_/D _9528_/SET_B VGND VGND VPWR VPWR _9502_/Q sky130_fd_sc_hd__dfstp_1
X_6714_ _6712_/Y _5374_/B _6713_/Y _5382_/B VGND VGND VPWR VPWR _6714_/X sky130_fd_sc_hd__o22a_1
X_9433_ _9440_/CLK _9433_/D _4628_/A VGND VGND VPWR VPWR _9433_/Q sky130_fd_sc_hd__dfrtp_1
X_7694_ _6434_/Y _7461_/X _6340_/Y _7463_/X _7693_/X VGND VGND VPWR VPWR _7697_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_32_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6645_ _9242_/Q VGND VGND VPWR VPWR _6645_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9364_ _9508_/CLK _9364_/D _9647_/SET_B VGND VGND VPWR VPWR _9364_/Q sky130_fd_sc_hd__dfstp_1
X_6576_ _9531_/Q VGND VGND VPWR VPWR _8779_/A sky130_fd_sc_hd__clkinv_8
XFILLER_192_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9295_ _9371_/CLK _9295_/D _9295_/SET_B VGND VGND VPWR VPWR _9295_/Q sky130_fd_sc_hd__dfstp_1
X_5527_ _5527_/A VGND VGND VPWR VPWR _5528_/A sky130_fd_sc_hd__clkbuf_2
X_8315_ _8238_/A _8498_/B _8304_/Y _8313_/X _8314_/X VGND VGND VPWR VPWR _8318_/A
+ sky130_fd_sc_hd__o2111ai_1
X_8246_ _8341_/A _8246_/B VGND VGND VPWR VPWR _8490_/B sky130_fd_sc_hd__nor2_1
X_5458_ _5545_/A _5458_/B VGND VGND VPWR VPWR _5459_/A sky130_fd_sc_hd__or2_1
X_5389_ _9453_/Q _5384_/A _8842_/X _5384_/Y VGND VGND VPWR VPWR _9453_/D sky130_fd_sc_hd__a22o_1
X_8177_ _8720_/A _8560_/A _8177_/C VGND VGND VPWR VPWR _8178_/B sky130_fd_sc_hd__or3_1
XFILLER_115_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7128_ _7128_/A VGND VGND VPWR VPWR _7128_/X sky130_fd_sc_hd__buf_8
XFILLER_101_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7059_ _7059_/A _7059_/B _7059_/C _7059_/D VGND VGND VPWR VPWR _7078_/B sky130_fd_sc_hd__and4_1
XFILLER_27_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_160 _4450_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_171 _7021_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_182 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_193 _4629_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4760_ _4927_/A _4780_/B VGND VGND VPWR VPWR _5610_/B sky130_fd_sc_hd__or2_4
XFILLER_81_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4691_ _4919_/A _4843_/B VGND VGND VPWR VPWR _5024_/B sky130_fd_sc_hd__or2_4
X_6430_ _9074_/Q VGND VGND VPWR VPWR _6430_/Y sky130_fd_sc_hd__inv_4
XFILLER_174_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6361_ _9311_/Q VGND VGND VPWR VPWR _6361_/Y sky130_fd_sc_hd__clkinv_2
X_8100_ _8100_/A VGND VGND VPWR VPWR _8213_/A sky130_fd_sc_hd__buf_12
X_5312_ _9506_/Q _5308_/A _8925_/A1 _5308_/Y VGND VGND VPWR VPWR _9506_/D sky130_fd_sc_hd__a22o_1
X_9080_ _9709_/CLK _9080_/D _6021_/X VGND VGND VPWR VPWR _9080_/Q sky130_fd_sc_hd__dfrtp_4
X_6292_ _6292_/A VGND VGND VPWR VPWR _6292_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_142_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8031_ _8097_/B _8550_/A _8030_/X VGND VGND VPWR VPWR _8033_/A sky130_fd_sc_hd__o21ai_1
X_5243_ _9553_/Q _5242_/A _8846_/X _5242_/Y VGND VGND VPWR VPWR _9553_/D sky130_fd_sc_hd__a22o_1
X_5174_ _9597_/Q _5169_/A _8842_/X _5169_/Y VGND VGND VPWR VPWR _9597_/D sky130_fd_sc_hd__a22o_1
XFILLER_142_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8933_ _9085_/Q _9084_/Q _9051_/Q VGND VGND VPWR VPWR _8933_/X sky130_fd_sc_hd__mux2_1
X_8864_ _7626_/Y _9627_/Q _8978_/S VGND VGND VPWR VPWR _8864_/X sky130_fd_sc_hd__mux2_1
X_7815_ _7815_/A VGND VGND VPWR VPWR _8097_/B sky130_fd_sc_hd__buf_12
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8795_ _8795_/A VGND VGND VPWR VPWR _8796_/A sky130_fd_sc_hd__clkbuf_1
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7746_ _9066_/Q _7746_/B VGND VGND VPWR VPWR _7746_/X sky130_fd_sc_hd__and2_1
XFILLER_101_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4958_ _9091_/Q _6022_/C VGND VGND VPWR VPWR _4958_/Y sky130_fd_sc_hd__nor2_1
XFILLER_184_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7677_ _6549_/Y _7475_/X _6510_/Y _7477_/X VGND VGND VPWR VPWR _7677_/X sky130_fd_sc_hd__o22a_1
X_4889_ _4911_/A _4900_/B VGND VGND VPWR VPWR _5298_/B sky130_fd_sc_hd__or2_4
X_9416_ _9684_/CLK _9416_/D _9685_/SET_B VGND VGND VPWR VPWR _9416_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_137_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6628_ _6628_/A _6628_/B _6628_/C _6628_/D VGND VGND VPWR VPWR _6629_/D sky130_fd_sc_hd__and4_2
XFILLER_118_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9347_ _9352_/CLK _9347_/D _9646_/SET_B VGND VGND VPWR VPWR _9347_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_106_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6559_ _6557_/Y _5450_/B _6558_/Y _4841_/X VGND VGND VPWR VPWR _6559_/X sky130_fd_sc_hd__o22a_1
XFILLER_193_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9278_ _9279_/CLK _9278_/D _9633_/SET_B VGND VGND VPWR VPWR _9278_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_126_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8229_ _8510_/A _8232_/B VGND VGND VPWR VPWR _8658_/B sky130_fd_sc_hd__nor2_1
XFILLER_10_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5930_ _5930_/A _5930_/B input150/X input153/X VGND VGND VPWR VPWR _5935_/B sky130_fd_sc_hd__or4bb_1
XFILLER_25_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7600_ _6122_/Y _7441_/X _6114_/Y _7443_/X _7599_/X VGND VGND VPWR VPWR _7607_/A
+ sky130_fd_sc_hd__o221a_1
X_5861_ _5849_/X _8851_/X _8924_/X _9165_/Q VGND VGND VPWR VPWR _9165_/D sky130_fd_sc_hd__o22a_1
X_8580_ _8580_/A _8675_/C _8645_/D _8716_/A VGND VGND VPWR VPWR _8586_/A sky130_fd_sc_hd__or4_4
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5792_ _9216_/Q _5791_/A _5963_/B1 _5791_/Y VGND VGND VPWR VPWR _9216_/D sky130_fd_sc_hd__a22o_1
X_4812_ _4800_/Y _5290_/B _4804_/Y _5534_/B _4811_/X VGND VGND VPWR VPWR _4830_/B
+ sky130_fd_sc_hd__o221a_1
X_4743_ _4876_/B _4780_/B VGND VGND VPWR VPWR _5572_/B sky130_fd_sc_hd__or2_4
X_7531_ _8751_/A _7465_/X _8789_/A _7467_/X VGND VGND VPWR VPWR _7531_/X sky130_fd_sc_hd__o22a_1
X_7462_ _7462_/A _7476_/C _7474_/D VGND VGND VPWR VPWR _7463_/A sky130_fd_sc_hd__or3_1
XFILLER_162_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9201_ _9789_/CLK _9201_/D _4628_/A VGND VGND VPWR VPWR _9201_/Q sky130_fd_sc_hd__dfrtp_1
X_4674_ _4660_/Y _5556_/B _4664_/Y _5905_/B _4673_/X VGND VGND VPWR VPWR _4705_/A
+ sky130_fd_sc_hd__o221a_1
X_6413_ _6411_/Y _4822_/X _6412_/Y _5232_/B VGND VGND VPWR VPWR _6413_/X sky130_fd_sc_hd__o22a_2
X_7393_ _6391_/Y _5728_/X _6418_/Y _7040_/A _7392_/X VGND VGND VPWR VPWR _7396_/C
+ sky130_fd_sc_hd__o221a_1
X_9132_ _9379_/CLK _9132_/D _9779_/SET_B VGND VGND VPWR VPWR _9132_/Q sky130_fd_sc_hd__dfrtp_1
X_6344_ _6342_/Y _4613_/B _6343_/Y _5564_/B VGND VGND VPWR VPWR _6344_/X sky130_fd_sc_hd__o22a_1
X_9063_ _4450_/A1 _9063_/D _6146_/A VGND VGND VPWR VPWR _9063_/Q sky130_fd_sc_hd__dfrtp_1
X_6275_ _9533_/Q VGND VGND VPWR VPWR _6275_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5226_ _9561_/Q _5218_/Y _8848_/X _5218_/A VGND VGND VPWR VPWR _9561_/D sky130_fd_sc_hd__o22a_1
X_8014_ _8521_/A _8117_/A _8013_/X VGND VGND VPWR VPWR _8016_/C sky130_fd_sc_hd__o21ai_1
Xinput109 sram_ro_data[24] VGND VGND VPWR VPWR _4831_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_130_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5157_ _5157_/A VGND VGND VPWR VPWR _5158_/A sky130_fd_sc_hd__clkbuf_4
X_5088_ _5133_/A VGND VGND VPWR VPWR _5545_/A sky130_fd_sc_hd__buf_12
X_8916_ _9610_/Q _8916_/A1 _8930_/S VGND VGND VPWR VPWR _8916_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8847_ _7022_/Y _9640_/Q _9587_/Q VGND VGND VPWR VPWR _8847_/X sky130_fd_sc_hd__mux2_1
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8778_ _8778_/A VGND VGND VPWR VPWR _8778_/X sky130_fd_sc_hd__clkbuf_1
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7729_ _7727_/Y _7726_/Y _9700_/Q VGND VGND VPWR VPWR _7729_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_165_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_71 _8544_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_93 input77/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_82 _7019_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_60 _6819_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6060_ _6060_/A VGND VGND VPWR VPWR _8807_/B sky130_fd_sc_hd__inv_4
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5011_ _6022_/B _7003_/C VGND VGND VPWR VPWR _5011_/X sky130_fd_sc_hd__or2_1
XFILLER_81_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6962_ _6974_/B _6962_/B VGND VGND VPWR VPWR _6963_/A sky130_fd_sc_hd__or2_2
X_9750_ _9755_/CLK _9750_/D _9757_/SET_B VGND VGND VPWR VPWR _9750_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_53_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8701_ _8064_/C _8700_/Y _8016_/C _8527_/C _8613_/B VGND VGND VPWR VPWR _8735_/C
+ sky130_fd_sc_hd__a2111o_2
X_6893_ _6891_/Y _5679_/B _6892_/Y _5488_/B VGND VGND VPWR VPWR _6893_/X sky130_fd_sc_hd__o22a_1
X_5913_ _9127_/Q _5907_/A _8955_/A1 _5907_/Y VGND VGND VPWR VPWR _9127_/D sky130_fd_sc_hd__a22o_1
XFILLER_34_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9681_ _9681_/CLK _9681_/D _6146_/A VGND VGND VPWR VPWR _9681_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_179_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5844_ _9180_/Q _5839_/A _8929_/A1 _5839_/Y VGND VGND VPWR VPWR _9180_/D sky130_fd_sc_hd__a22o_1
X_8632_ _8632_/A _8632_/B VGND VGND VPWR VPWR _8687_/C sky130_fd_sc_hd__nor2_1
XFILLER_22_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8563_ _8563_/A _8713_/D _8713_/B _8636_/D VGND VGND VPWR VPWR _8563_/X sky130_fd_sc_hd__or4_1
XFILLER_166_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7514_ _6687_/Y _7461_/X _6735_/Y _7463_/X _7513_/X VGND VGND VPWR VPWR _7517_/C
+ sky130_fd_sc_hd__o221a_1
X_5775_ _9226_/Q _5770_/A _5967_/B1 _5770_/Y VGND VGND VPWR VPWR _9226_/D sky130_fd_sc_hd__a22o_1
XFILLER_159_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4726_ _9269_/Q VGND VGND VPWR VPWR _4726_/Y sky130_fd_sc_hd__clkinv_2
X_8494_ _8515_/B _8305_/A _8660_/A _8496_/A _8341_/B VGND VGND VPWR VPWR _8594_/A
+ sky130_fd_sc_hd__a311oi_2
XFILLER_162_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7445_ _7445_/A VGND VGND VPWR VPWR _7445_/X sky130_fd_sc_hd__buf_8
X_4657_ _4657_/A VGND VGND VPWR VPWR _4657_/X sky130_fd_sc_hd__clkbuf_1
Xinput91 spimemio_flash_io3_do VGND VGND VPWR VPWR input91/X sky130_fd_sc_hd__clkbuf_4
XFILLER_174_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput80 spi_sck VGND VGND VPWR VPWR input80/X sky130_fd_sc_hd__buf_6
X_7376_ _6348_/Y _7086_/X _6409_/Y _7088_/X VGND VGND VPWR VPWR _7376_/X sky130_fd_sc_hd__o22a_1
X_6327_ _6149_/A _6326_/Y _9041_/Q _6149_/Y VGND VGND VPWR VPWR _9041_/D sky130_fd_sc_hd__o22a_1
XFILLER_162_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9115_ _9129_/CLK _9115_/D _9779_/SET_B VGND VGND VPWR VPWR _9115_/Q sky130_fd_sc_hd__dfrtp_1
X_4588_ _4669_/A _4729_/D _8946_/X _4729_/B VGND VGND VPWR VPWR _4903_/B sky130_fd_sc_hd__or4_4
XFILLER_115_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9046_ _9790_/CLK _9046_/D VGND VGND VPWR VPWR _9046_/Q sky130_fd_sc_hd__dfxtp_1
X_6258_ _9737_/Q VGND VGND VPWR VPWR _6258_/Y sky130_fd_sc_hd__inv_2
XFILLER_191_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5209_ _9572_/Q _5203_/Y _8905_/X _5203_/A VGND VGND VPWR VPWR _9572_/D sky130_fd_sc_hd__o22a_1
XFILLER_29_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6189_ _9784_/Q VGND VGND VPWR VPWR _6189_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5560_ _9336_/Q _5558_/A _8842_/X _5558_/Y VGND VGND VPWR VPWR _9336_/D sky130_fd_sc_hd__a22o_1
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5491_ _9384_/Q _5490_/A _5963_/B1 _5490_/Y VGND VGND VPWR VPWR _9384_/D sky130_fd_sc_hd__a22o_1
X_4511_ _9773_/Q _4506_/A _5967_/B1 _4506_/Y VGND VGND VPWR VPWR _9773_/D sky130_fd_sc_hd__a22o_1
XFILLER_144_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7230_ _6296_/Y _7059_/B _6310_/Y _7068_/C _7229_/X VGND VGND VPWR VPWR _7233_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_117_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7161_ _6760_/Y _7097_/X _6735_/Y _7099_/X VGND VGND VPWR VPWR _7161_/X sky130_fd_sc_hd__o22a_1
XFILLER_98_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6112_ _6109_/Y _5267_/B _6110_/Y _5306_/B _6111_/X VGND VGND VPWR VPWR _6119_/C
+ sky130_fd_sc_hd__o221a_1
X_7092_ _4773_/Y _7040_/C _4664_/Y _7059_/C VGND VGND VPWR VPWR _7092_/X sky130_fd_sc_hd__o22a_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6043_ _6043_/A VGND VGND VPWR VPWR _6043_/X sky130_fd_sc_hd__clkbuf_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7994_ _7994_/A _7994_/B VGND VGND VPWR VPWR _8116_/B sky130_fd_sc_hd__nand2_4
XFILLER_39_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6945_ _6945_/A _6945_/B _6945_/C VGND VGND VPWR VPWR _6946_/C sky130_fd_sc_hd__and3_2
X_9733_ _9774_/CLK _9733_/D _9757_/SET_B VGND VGND VPWR VPWR _9733_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_54_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_2_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
X_9664_ _9664_/CLK _9664_/D _6146_/A VGND VGND VPWR VPWR _9664_/Q sky130_fd_sc_hd__dfrtp_1
X_6876_ _6871_/Y _5458_/B _6872_/Y _5480_/B _6875_/X VGND VGND VPWR VPWR _6877_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9595_ _9596_/CLK _9595_/D _9528_/SET_B VGND VGND VPWR VPWR _9595_/Q sky130_fd_sc_hd__dfrtp_1
X_5827_ _9191_/Q _5820_/A _8930_/A1 _5820_/Y VGND VGND VPWR VPWR _9191_/D sky130_fd_sc_hd__a22o_1
X_8615_ _8615_/A _8615_/B _8615_/C _8615_/D VGND VGND VPWR VPWR _8699_/C sky130_fd_sc_hd__or4_1
X_5758_ _5758_/A VGND VGND VPWR VPWR _5759_/A sky130_fd_sc_hd__clkbuf_4
X_8546_ _8546_/A _8566_/B VGND VGND VPWR VPWR _8546_/Y sky130_fd_sc_hd__nor2_1
XFILLER_163_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8477_ _8477_/A _8721_/C VGND VGND VPWR VPWR _8478_/B sky130_fd_sc_hd__or2_1
XFILLER_135_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4709_ _4929_/A _4780_/B VGND VGND VPWR VPWR _5776_/B sky130_fd_sc_hd__or2_4
X_5689_ _9256_/Q _5681_/A _8916_/A1 _5681_/Y VGND VGND VPWR VPWR _9256_/D sky130_fd_sc_hd__a22o_1
XFILLER_175_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7428_ _4816_/Y _7427_/X _4742_/Y _5699_/X VGND VGND VPWR VPWR _7428_/X sky130_fd_sc_hd__o22a_1
XFILLER_162_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7359_ _6604_/Y _7097_/X _6550_/Y _7099_/X VGND VGND VPWR VPWR _7359_/X sky130_fd_sc_hd__o22a_1
XFILLER_78_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9029_ _9039_/CLK _9029_/D VGND VGND VPWR VPWR _9029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6730_ _9512_/Q VGND VGND VPWR VPWR _6730_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_23_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4991_ _4991_/A _8957_/X VGND VGND VPWR VPWR _5001_/S sky130_fd_sc_hd__or2b_1
XFILLER_189_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6661_ _9322_/Q VGND VGND VPWR VPWR _6661_/Y sky130_fd_sc_hd__clkinv_2
X_5612_ _5612_/A VGND VGND VPWR VPWR _5612_/Y sky130_fd_sc_hd__clkinv_2
X_8400_ _8521_/A _8117_/A _8393_/Y _8401_/B _8399_/X VGND VGND VPWR VPWR _8400_/X
+ sky130_fd_sc_hd__o221a_1
X_9380_ _9380_/CLK _9380_/D _4628_/A VGND VGND VPWR VPWR _9380_/Q sky130_fd_sc_hd__dfrtp_1
X_6592_ input6/X VGND VGND VPWR VPWR _6592_/Y sky130_fd_sc_hd__inv_2
X_8331_ _8331_/A _8331_/B VGND VGND VPWR VPWR _8331_/X sky130_fd_sc_hd__or2_1
X_5543_ _9347_/Q _5536_/A _8930_/A1 _5536_/Y VGND VGND VPWR VPWR _9347_/D sky130_fd_sc_hd__a22o_1
XFILLER_129_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5474_ _9395_/Q _5471_/A _8844_/X _5471_/Y VGND VGND VPWR VPWR _9395_/D sky130_fd_sc_hd__a22o_1
XFILLER_144_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8262_ _8341_/A _8262_/B VGND VGND VPWR VPWR _8369_/B sky130_fd_sc_hd__nor2_1
X_8193_ _8193_/A _8193_/B _8195_/A VGND VGND VPWR VPWR _8204_/A sky130_fd_sc_hd__or3_2
XFILLER_160_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7213_ _6457_/Y _7040_/D _6398_/Y _7110_/X _7212_/X VGND VGND VPWR VPWR _7220_/A
+ sky130_fd_sc_hd__o221a_1
X_7144_ _6879_/Y _7048_/D _6908_/Y _7040_/B _7143_/X VGND VGND VPWR VPWR _7145_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_98_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7075_ _7075_/A _7123_/B VGND VGND VPWR VPWR _7076_/A sky130_fd_sc_hd__or2_1
XFILLER_58_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6026_ _9078_/Q _4466_/A _8955_/A1 _4466_/Y VGND VGND VPWR VPWR _9078_/D sky130_fd_sc_hd__a22o_1
XFILLER_39_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7977_ _8091_/B _7988_/A VGND VGND VPWR VPWR _8096_/A sky130_fd_sc_hd__nand2_4
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6928_ _9265_/Q VGND VGND VPWR VPWR _6928_/Y sky130_fd_sc_hd__clkinv_2
X_9716_ _9089_/CLK _9716_/D _4642_/X VGND VGND VPWR VPWR hold1/A sky130_fd_sc_hd__dfrtn_1
XFILLER_167_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9647_ _9652_/CLK _9647_/D _9647_/SET_B VGND VGND VPWR VPWR _9647_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6859_ _9373_/Q VGND VGND VPWR VPWR _6859_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9578_ _9674_/CLK _9578_/D _9633_/SET_B VGND VGND VPWR VPWR _9578_/Q sky130_fd_sc_hd__dfrtp_1
X_8529_ _8523_/Y _8528_/Y _8518_/X _8455_/B VGND VGND VPWR VPWR _8734_/D sky130_fd_sc_hd__a31o_1
XFILLER_182_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_3_0_mgmt_gpio_in[4] clkbuf_2_3_0_mgmt_gpio_in[4]/A VGND VGND VPWR VPWR _4446_/A1
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_173_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5190_ _5190_/A VGND VGND VPWR VPWR _5190_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_95_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7900_ _7900_/A _8528_/B VGND VGND VPWR VPWR _8517_/A sky130_fd_sc_hd__or2b_2
XFILLER_110_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8880_ _7221_/Y _9636_/Q _8959_/S VGND VGND VPWR VPWR _8880_/X sky130_fd_sc_hd__mux2_1
X_7831_ _8324_/A VGND VGND VPWR VPWR _7831_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4974_ _4994_/A VGND VGND VPWR VPWR _4975_/A sky130_fd_sc_hd__clkbuf_1
X_7762_ _8379_/D VGND VGND VPWR VPWR _8394_/A sky130_fd_sc_hd__clkinv_4
X_6713_ _9452_/Q VGND VGND VPWR VPWR _6713_/Y sky130_fd_sc_hd__inv_2
X_9501_ _9501_/CLK _9501_/D _9647_/SET_B VGND VGND VPWR VPWR _9501_/Q sky130_fd_sc_hd__dfrtp_1
X_7693_ _6369_/Y _7465_/X _6397_/Y _7467_/X VGND VGND VPWR VPWR _7693_/X sky130_fd_sc_hd__o22a_1
X_6644_ _9192_/Q VGND VGND VPWR VPWR _6644_/Y sky130_fd_sc_hd__inv_2
X_9432_ _9440_/CLK _9432_/D _4628_/A VGND VGND VPWR VPWR _9432_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_109_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6575_ _9375_/Q VGND VGND VPWR VPWR _8767_/A sky130_fd_sc_hd__clkinv_8
X_9363_ _9771_/CLK _9363_/D _4628_/A VGND VGND VPWR VPWR _9363_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9294_ _9371_/CLK _9294_/D _9295_/SET_B VGND VGND VPWR VPWR _9294_/Q sky130_fd_sc_hd__dfstp_1
X_5526_ _5671_/A _5526_/B VGND VGND VPWR VPWR _5527_/A sky130_fd_sc_hd__or2_1
X_8314_ _8316_/A _8264_/B _8454_/A VGND VGND VPWR VPWR _8314_/X sky130_fd_sc_hd__o21a_1
XFILLER_160_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8245_ _8245_/A _8362_/B _8575_/B VGND VGND VPWR VPWR _8248_/A sky130_fd_sc_hd__or3_1
X_5457_ _9406_/Q _5452_/A _5967_/B1 _5452_/Y VGND VGND VPWR VPWR _9406_/D sky130_fd_sc_hd__a22o_1
XFILLER_105_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5388_ _9454_/Q _5384_/A _8925_/A1 _5384_/Y VGND VGND VPWR VPWR _9454_/D sky130_fd_sc_hd__a22o_1
X_8176_ _8521_/A _8515_/A _8175_/Y VGND VGND VPWR VPWR _8177_/C sky130_fd_sc_hd__o21bai_1
XFILLER_120_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7127_ _7127_/A _7127_/B _7127_/C VGND VGND VPWR VPWR _7128_/A sky130_fd_sc_hd__or3_1
XFILLER_47_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7058_ _7058_/A VGND VGND VPWR VPWR _7059_/D sky130_fd_sc_hd__buf_8
XFILLER_101_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6009_ _6040_/A VGND VGND VPWR VPWR _6010_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_46_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_161 _9404_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_150 _6829_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_172 _7021_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_183 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_194 input82/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4690_ _9683_/Q VGND VGND VPWR VPWR _4692_/A sky130_fd_sc_hd__clkinv_4
XFILLER_174_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6360_ _9324_/Q VGND VGND VPWR VPWR _6360_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5311_ _9507_/Q _5308_/A _8844_/X _5308_/Y VGND VGND VPWR VPWR _9507_/D sky130_fd_sc_hd__a22o_1
XFILLER_127_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6291_ _9075_/Q VGND VGND VPWR VPWR _6291_/Y sky130_fd_sc_hd__inv_6
XFILLER_114_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8030_ _8389_/A _8550_/A _8027_/X _8410_/A _8029_/X VGND VGND VPWR VPWR _8030_/X
+ sky130_fd_sc_hd__o2111a_1
X_5242_ _5242_/A VGND VGND VPWR VPWR _5242_/Y sky130_fd_sc_hd__inv_2
X_5173_ _9598_/Q _5169_/A _8925_/A1 _5169_/Y VGND VGND VPWR VPWR _9598_/D sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_30_csclk clkbuf_2_1_0_csclk/X VGND VGND VPWR VPWR _9129_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_96_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput1 debug_mode VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_45_csclk _9329_/CLK VGND VGND VPWR VPWR _9777_/CLK sky130_fd_sc_hd__clkbuf_16
X_8932_ _8931_/X _9677_/Q _9587_/Q VGND VGND VPWR VPWR _8932_/X sky130_fd_sc_hd__mux2_4
XFILLER_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8863_ _8862_/X _9170_/Q _9054_/Q VGND VGND VPWR VPWR _8863_/X sky130_fd_sc_hd__mux2_1
X_7814_ _8379_/C _7839_/A _8394_/A _8394_/B VGND VGND VPWR VPWR _7815_/A sky130_fd_sc_hd__or4_1
XFILLER_24_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8794_ _8794_/A VGND VGND VPWR VPWR _8794_/X sky130_fd_sc_hd__clkbuf_1
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7745_ _9068_/Q _7745_/A2 _9067_/Q _7745_/B2 _7744_/X VGND VGND VPWR VPWR _7745_/X
+ sky130_fd_sc_hd__a221o_1
X_4957_ _4957_/A VGND VGND VPWR VPWR _4957_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_177_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7676_ _6486_/Y _7461_/X _6550_/Y _7463_/X _7675_/X VGND VGND VPWR VPWR _7679_/C
+ sky130_fd_sc_hd__o221a_1
X_4888_ _9510_/Q VGND VGND VPWR VPWR _4888_/Y sky130_fd_sc_hd__inv_2
XFILLER_192_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9415_ _9514_/CLK _9415_/D _4628_/A VGND VGND VPWR VPWR _9415_/Q sky130_fd_sc_hd__dfrtp_1
X_6627_ _6627_/A _6627_/B _6627_/C _6627_/D VGND VGND VPWR VPWR _6628_/D sky130_fd_sc_hd__and4_1
XFILLER_192_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9346_ _9352_/CLK _9346_/D _9646_/SET_B VGND VGND VPWR VPWR _9346_/Q sky130_fd_sc_hd__dfstp_1
X_6558_ _6558_/A VGND VGND VPWR VPWR _6558_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_106_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6489_ _9393_/Q VGND VGND VPWR VPWR _8797_/A sky130_fd_sc_hd__inv_4
X_5509_ _5509_/A VGND VGND VPWR VPWR _5509_/Y sky130_fd_sc_hd__inv_2
XFILLER_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9277_ _9280_/CLK _9277_/D _9757_/SET_B VGND VGND VPWR VPWR _9277_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_160_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8228_ _8230_/A _8264_/B VGND VGND VPWR VPWR _8676_/B sky130_fd_sc_hd__nor2_2
X_8159_ _8554_/A _8640_/B VGND VGND VPWR VPWR _8645_/A sky130_fd_sc_hd__nor2_1
XFILLER_86_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5860_ _5849_/X _8853_/X _8924_/X _9166_/Q VGND VGND VPWR VPWR _9166_/D sky130_fd_sc_hd__o22a_1
XFILLER_92_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4811_ _4931_/A _6158_/A _4808_/Y _4809_/Y _5251_/B VGND VGND VPWR VPWR _4811_/X
+ sky130_fd_sc_hd__o32a_1
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5791_ _5791_/A VGND VGND VPWR VPWR _5791_/Y sky130_fd_sc_hd__inv_2
XFILLER_178_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4742_ _9320_/Q VGND VGND VPWR VPWR _4742_/Y sky130_fd_sc_hd__inv_2
X_7530_ _8749_/A _7451_/X _8773_/A _7453_/X _7529_/X VGND VGND VPWR VPWR _7535_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_21_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4673_ _4668_/Y _5872_/B _4671_/Y _5526_/B VGND VGND VPWR VPWR _4673_/X sky130_fd_sc_hd__o22a_1
X_7461_ _7461_/A VGND VGND VPWR VPWR _7461_/X sky130_fd_sc_hd__buf_8
X_9200_ _9789_/CLK _9200_/D _4628_/A VGND VGND VPWR VPWR _9200_/Q sky130_fd_sc_hd__dfstp_1
X_6412_ _9558_/Q VGND VGND VPWR VPWR _6412_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_opt_5_0_csclk clkbuf_2_2_0_csclk/X VGND VGND VPWR VPWR clkbuf_leaf_6_csclk/A
+ sky130_fd_sc_hd__clkbuf_16
X_7392_ _7392_/A _7392_/B VGND VGND VPWR VPWR _7392_/X sky130_fd_sc_hd__or2_1
XFILLER_127_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9131_ _9379_/CLK _9131_/D _9779_/SET_B VGND VGND VPWR VPWR _9131_/Q sky130_fd_sc_hd__dfrtp_1
X_6343_ _9332_/Q VGND VGND VPWR VPWR _6343_/Y sky130_fd_sc_hd__inv_2
X_6274_ _9455_/Q VGND VGND VPWR VPWR _6274_/Y sky130_fd_sc_hd__clkinv_4
X_9062_ _4450_/A1 _9062_/D _6146_/A VGND VGND VPWR VPWR _9062_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_115_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5225_ _9562_/Q _5218_/Y _8919_/X _5218_/A VGND VGND VPWR VPWR _9562_/D sky130_fd_sc_hd__o22a_1
X_8013_ _8097_/B _8013_/B VGND VGND VPWR VPWR _8013_/X sky130_fd_sc_hd__or2_1
XFILLER_130_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5156_ _6135_/A _5156_/B VGND VGND VPWR VPWR _5157_/A sky130_fd_sc_hd__or2_1
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5087_ _9654_/Q _5082_/A _5967_/B1 _5082_/Y VGND VGND VPWR VPWR _9654_/D sky130_fd_sc_hd__a22o_1
X_8915_ _9623_/Q _8844_/X _8955_/S VGND VGND VPWR VPWR _8915_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8846_ _9707_/Q _9666_/Q _9587_/Q VGND VGND VPWR VPWR _8846_/X sky130_fd_sc_hd__mux2_8
XFILLER_52_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8777_ _8777_/A VGND VGND VPWR VPWR _8778_/A sky130_fd_sc_hd__clkbuf_1
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5989_ _6022_/C _5985_/B _5985_/Y VGND VGND VPWR VPWR _9090_/D sky130_fd_sc_hd__a21oi_1
XFILLER_24_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7728_ _7727_/Y _7726_/Y _9699_/Q _9698_/Q VGND VGND VPWR VPWR _7728_/X sky130_fd_sc_hd__a22o_1
XFILLER_177_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_50 _7216_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_72 _8375_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7659_ _6652_/Y _7475_/X _6634_/Y _7477_/X VGND VGND VPWR VPWR _7659_/X sky130_fd_sc_hd__o22a_1
XANTENNA_83 _7019_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_61 _6832_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_94 input77/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9329_ _9329_/CLK _9329_/D _4628_/A VGND VGND VPWR VPWR _9329_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_97_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_4_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A VGND VGND VPWR VPWR _9027_/CLK sky130_fd_sc_hd__clkbuf_2
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _5010_/A VGND VGND VPWR VPWR _5010_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_85_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6961_ _9062_/Q VGND VGND VPWR VPWR _6962_/B sky130_fd_sc_hd__inv_2
X_8700_ _8515_/B _8305_/A _8341_/B VGND VGND VPWR VPWR _8700_/Y sky130_fd_sc_hd__a21oi_1
X_5912_ _9128_/Q _5907_/A _8929_/A1 _5907_/Y VGND VGND VPWR VPWR _9128_/D sky130_fd_sc_hd__a22o_1
X_6892_ _9381_/Q VGND VGND VPWR VPWR _6892_/Y sky130_fd_sc_hd__clkinv_2
X_9680_ _9681_/CLK _9680_/D _6146_/A VGND VGND VPWR VPWR _9680_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_53_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5843_ _9181_/Q _5839_/A _8925_/A1 _5839_/Y VGND VGND VPWR VPWR _9181_/D sky130_fd_sc_hd__a22o_1
X_8631_ _8631_/A _8631_/B VGND VGND VPWR VPWR _8688_/C sky130_fd_sc_hd__or2_1
XFILLER_179_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8562_ _8562_/A _8672_/C _8673_/A VGND VGND VPWR VPWR _8636_/D sky130_fd_sc_hd__or3_1
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7513_ _6637_/Y _7465_/X _6717_/Y _7467_/X VGND VGND VPWR VPWR _7513_/X sky130_fd_sc_hd__o22a_1
X_5774_ _9227_/Q _5770_/A _5966_/B1 _5770_/Y VGND VGND VPWR VPWR _9227_/D sky130_fd_sc_hd__a22o_1
X_4725_ _4716_/Y _5837_/B _4718_/Y _5594_/B _4724_/X VGND VGND VPWR VPWR _4791_/B
+ sky130_fd_sc_hd__o221a_1
X_8493_ _8614_/A _8493_/B _8493_/C VGND VGND VPWR VPWR _8657_/C sky130_fd_sc_hd__or3_1
XFILLER_135_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7444_ _7462_/A _7470_/B _7474_/D VGND VGND VPWR VPWR _7445_/A sky130_fd_sc_hd__or3_1
X_4656_ _4994_/A VGND VGND VPWR VPWR _4657_/A sky130_fd_sc_hd__clkbuf_1
Xinput81 spi_sdo VGND VGND VPWR VPWR input81/X sky130_fd_sc_hd__buf_6
X_7375_ _7375_/A _7375_/B _7375_/C VGND VGND VPWR VPWR _7375_/Y sky130_fd_sc_hd__nand3_4
Xinput70 mgmt_gpio_in[7] VGND VGND VPWR VPWR _6060_/A sky130_fd_sc_hd__clkbuf_1
X_4587_ _9740_/Q _4579_/A _5967_/B1 _4579_/Y VGND VGND VPWR VPWR _9740_/D sky130_fd_sc_hd__a22o_1
Xinput92 spimemio_flash_io3_oeb VGND VGND VPWR VPWR input92/X sky130_fd_sc_hd__buf_2
XFILLER_162_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6326_ _6326_/A _6326_/B _6326_/C _6326_/D VGND VGND VPWR VPWR _6326_/Y sky130_fd_sc_hd__nand4_4
X_9114_ _9779_/CLK _9114_/D _9779_/SET_B VGND VGND VPWR VPWR _9114_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_130_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9045_ _9790_/CLK _9045_/D VGND VGND VPWR VPWR _9045_/Q sky130_fd_sc_hd__dfxtp_1
X_6257_ _6257_/A VGND VGND VPWR VPWR _6257_/Y sky130_fd_sc_hd__inv_2
XFILLER_190_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6188_ _9076_/Q VGND VGND VPWR VPWR _6188_/Y sky130_fd_sc_hd__clkinv_4
X_5208_ _9573_/Q _5203_/Y _8929_/X _5203_/A VGND VGND VPWR VPWR _9573_/D sky130_fd_sc_hd__o22a_1
XFILLER_130_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5139_ _9623_/Q _5136_/A _8844_/X _5136_/Y VGND VGND VPWR VPWR _9623_/D sky130_fd_sc_hd__a22o_1
XFILLER_29_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8829_ _9592_/Q input89/X _8835_/S VGND VGND VPWR VPWR _8829_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5490_ _5490_/A VGND VGND VPWR VPWR _5490_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4510_ _9774_/Q _4506_/A _5966_/B1 _4506_/Y VGND VGND VPWR VPWR _9774_/D sky130_fd_sc_hd__a22o_1
XFILLER_156_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7160_ _6644_/Y _7048_/B _6681_/Y _7077_/A _7159_/X VGND VGND VPWR VPWR _7167_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_171_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6111_ _6111_/A _6111_/B _9769_/Q VGND VGND VPWR VPWR _6111_/X sky130_fd_sc_hd__or3b_4
X_7091_ _4855_/Y _7082_/X _4850_/Y _7084_/X _7090_/X VGND VGND VPWR VPWR _7132_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_112_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6042_ _6050_/A VGND VGND VPWR VPWR _6043_/A sky130_fd_sc_hd__clkbuf_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7993_ _7993_/A VGND VGND VPWR VPWR _8137_/B sky130_fd_sc_hd__buf_4
X_6944_ _6944_/A _6944_/B _6944_/C VGND VGND VPWR VPWR _6945_/C sky130_fd_sc_hd__and3_1
XFILLER_81_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9732_ _9774_/CLK _9732_/D _9757_/SET_B VGND VGND VPWR VPWR _9732_/Q sky130_fd_sc_hd__dfstp_1
X_9663_ _9664_/CLK _9663_/D _6146_/A VGND VGND VPWR VPWR _9663_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8614_ _8614_/A _8614_/B _8614_/C _8614_/D VGND VGND VPWR VPWR _8668_/D sky130_fd_sc_hd__or4_1
X_6875_ _6873_/Y _5404_/B _6874_/Y _5290_/B VGND VGND VPWR VPWR _6875_/X sky130_fd_sc_hd__o22a_1
XFILLER_22_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9594_ _9596_/CLK _9594_/D _9528_/SET_B VGND VGND VPWR VPWR _9594_/Q sky130_fd_sc_hd__dfrtp_1
X_5826_ _9192_/Q _5820_/A _8955_/A1 _5820_/Y VGND VGND VPWR VPWR _9192_/D sky130_fd_sc_hd__a22o_1
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5757_ _6052_/A _5757_/B VGND VGND VPWR VPWR _5758_/A sky130_fd_sc_hd__or2_1
X_8545_ _8625_/B VGND VGND VPWR VPWR _8554_/B sky130_fd_sc_hd__clkinv_4
XFILLER_182_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8476_ _8476_/A _8476_/B VGND VGND VPWR VPWR _8721_/C sky130_fd_sc_hd__or2_2
X_4708_ _9218_/Q VGND VGND VPWR VPWR _4708_/Y sky130_fd_sc_hd__inv_2
X_5688_ _9257_/Q _5681_/A _8840_/X _5681_/Y VGND VGND VPWR VPWR _9257_/D sky130_fd_sc_hd__a22o_1
XFILLER_162_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7427_ _7427_/A VGND VGND VPWR VPWR _7427_/X sky130_fd_sc_hd__buf_8
X_4639_ _4639_/A VGND VGND VPWR VPWR _4639_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7358_ _6504_/Y _7048_/B _6539_/Y _7077_/A _7357_/X VGND VGND VPWR VPWR _7365_/A
+ sky130_fd_sc_hd__o221a_2
X_6309_ _9261_/Q VGND VGND VPWR VPWR _6309_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7289_ _4731_/A _7077_/C _4671_/Y _7077_/D _7288_/X VGND VGND VPWR VPWR _7289_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9028_ _9039_/CLK _9028_/D VGND VGND VPWR VPWR _9028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4990_ _7008_/A _5992_/B _4966_/A _6022_/B _4989_/X VGND VGND VPWR VPWR _4991_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_149_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6660_ _6656_/Y _4524_/B _6657_/Y _5412_/B _6659_/X VGND VGND VPWR VPWR _6691_/B
+ sky130_fd_sc_hd__o221a_1
X_5611_ _5611_/A VGND VGND VPWR VPWR _5612_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_149_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6591_ _9751_/Q VGND VGND VPWR VPWR _6591_/Y sky130_fd_sc_hd__inv_2
X_8330_ _8376_/A _8330_/B VGND VGND VPWR VPWR _8331_/B sky130_fd_sc_hd__or2_1
X_5542_ _9348_/Q _5536_/A _8955_/A1 _5536_/Y VGND VGND VPWR VPWR _9348_/D sky130_fd_sc_hd__a22o_1
XFILLER_129_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5473_ _9396_/Q _5471_/A _8845_/X _5471_/Y VGND VGND VPWR VPWR _9396_/D sky130_fd_sc_hd__a22o_1
X_8261_ _8261_/A _8578_/B VGND VGND VPWR VPWR _8263_/A sky130_fd_sc_hd__or2_1
X_8192_ _8195_/A _8193_/B _8193_/A VGND VGND VPWR VPWR _8346_/A sky130_fd_sc_hd__o21a_1
X_7212_ _6360_/Y _7112_/X _6468_/Y _7077_/B VGND VGND VPWR VPWR _7212_/X sky130_fd_sc_hd__o22a_1
XFILLER_125_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7143_ _6890_/Y _7068_/A _6860_/Y _7105_/X VGND VGND VPWR VPWR _7143_/X sky130_fd_sc_hd__o22a_1
XFILLER_140_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7074_ _7074_/A VGND VGND VPWR VPWR _7077_/C sky130_fd_sc_hd__buf_8
XFILLER_59_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6025_ _9079_/Q _4466_/A _8844_/X _4466_/Y VGND VGND VPWR VPWR _9079_/D sky130_fd_sc_hd__a22o_1
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7976_ _8583_/A _7966_/B _8195_/B VGND VGND VPWR VPWR _7988_/A sky130_fd_sc_hd__a21bo_1
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9715_ _9089_/CLK _9715_/D _4645_/X VGND VGND VPWR VPWR _9715_/Q sky130_fd_sc_hd__dfrtn_1
X_6927_ _9241_/Q VGND VGND VPWR VPWR _6927_/Y sky130_fd_sc_hd__inv_2
X_9646_ _9652_/CLK _9646_/D _9646_/SET_B VGND VGND VPWR VPWR _9646_/Q sky130_fd_sc_hd__dfstp_1
X_6858_ _6853_/Y _5382_/B _6854_/Y _5306_/B _6857_/X VGND VGND VPWR VPWR _6877_/A
+ sky130_fd_sc_hd__o221a_2
X_9577_ _9788_/CLK _9577_/D _9295_/SET_B VGND VGND VPWR VPWR _9577_/Q sky130_fd_sc_hd__dfrtp_1
X_5809_ _9053_/Q _9791_/Q _5643_/Y _5808_/X VGND VGND VPWR VPWR _9203_/D sky130_fd_sc_hd__a31o_1
XFILLER_182_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8528_ _8528_/A _8528_/B VGND VGND VPWR VPWR _8528_/Y sky130_fd_sc_hd__nor2_4
X_6789_ _9727_/Q VGND VGND VPWR VPWR _6789_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8459_ _8459_/A _8734_/C _8459_/C _8614_/C VGND VGND VPWR VPWR _8464_/A sky130_fd_sc_hd__or4_1
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7830_ _7903_/C _8528_/A _8583_/A _8189_/A VGND VGND VPWR VPWR _8324_/A sky130_fd_sc_hd__or4_4
X_4973_ _9705_/Q _4966_/A _9704_/Q _4966_/Y VGND VGND VPWR VPWR _9705_/D sky130_fd_sc_hd__a22o_1
X_7761_ _8299_/A _8282_/C _7836_/A VGND VGND VPWR VPWR _8636_/A sky130_fd_sc_hd__and3_2
XFILLER_91_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6712_ _9460_/Q VGND VGND VPWR VPWR _6712_/Y sky130_fd_sc_hd__inv_2
X_9500_ _9501_/CLK _9500_/D _9647_/SET_B VGND VGND VPWR VPWR _9500_/Q sky130_fd_sc_hd__dfrtp_1
X_7692_ _6467_/Y _7451_/X _6348_/Y _7453_/X _7691_/X VGND VGND VPWR VPWR _7697_/B
+ sky130_fd_sc_hd__o221a_1
X_9431_ _9508_/CLK _9431_/D _9295_/SET_B VGND VGND VPWR VPWR _9431_/Q sky130_fd_sc_hd__dfrtp_1
X_6643_ _9233_/Q VGND VGND VPWR VPWR _6643_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6574_ _9513_/Q VGND VGND VPWR VPWR _6574_/Y sky130_fd_sc_hd__inv_2
X_9362_ _9514_/CLK _9362_/D _4628_/A VGND VGND VPWR VPWR _9362_/Q sky130_fd_sc_hd__dfrtp_1
X_9293_ _9596_/CLK _9293_/D _9528_/SET_B VGND VGND VPWR VPWR _9293_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_145_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8313_ _8496_/A _8306_/X _8230_/A _8498_/B _8312_/X VGND VGND VPWR VPWR _8313_/X
+ sky130_fd_sc_hd__o221a_2
X_5525_ _9359_/Q _5520_/A _5967_/B1 _5520_/Y VGND VGND VPWR VPWR _9359_/D sky130_fd_sc_hd__a22o_1
XFILLER_160_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8244_ _8316_/A _8260_/B VGND VGND VPWR VPWR _8575_/B sky130_fd_sc_hd__nor2_1
X_5456_ _9407_/Q _5452_/A _5966_/B1 _5452_/Y VGND VGND VPWR VPWR _9407_/D sky130_fd_sc_hd__a22o_1
XFILLER_145_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5387_ _9455_/Q _5384_/A _8844_/X _5384_/Y VGND VGND VPWR VPWR _9455_/D sky130_fd_sc_hd__a22o_1
XFILLER_160_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8175_ _8175_/A _8175_/B VGND VGND VPWR VPWR _8175_/Y sky130_fd_sc_hd__nand2_1
XFILLER_113_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7126_ _7126_/A VGND VGND VPWR VPWR _7126_/X sky130_fd_sc_hd__buf_8
XFILLER_140_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7057_ _7073_/C _7087_/B VGND VGND VPWR VPWR _7058_/A sky130_fd_sc_hd__or2_1
XFILLER_101_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6008_ _9085_/Q _5995_/A _8910_/X _5995_/Y VGND VGND VPWR VPWR _9085_/D sky130_fd_sc_hd__a22o_1
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7959_ _7959_/A _8583_/A _7966_/B VGND VGND VPWR VPWR _8193_/B sky130_fd_sc_hd__or3_2
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9629_ _9757_/CLK _9629_/D _9757_/SET_B VGND VGND VPWR VPWR _9629_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_24_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_151 _6902_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_140 _5013_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_173 _7021_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_184 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_162 _6629_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_195 _6271_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6290_ _9481_/Q VGND VGND VPWR VPWR _6290_/Y sky130_fd_sc_hd__inv_6
X_5310_ _9508_/Q _5308_/A _8845_/X _5308_/Y VGND VGND VPWR VPWR _9508_/D sky130_fd_sc_hd__a22o_1
XFILLER_115_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5241_ _5241_/A VGND VGND VPWR VPWR _5242_/A sky130_fd_sc_hd__clkbuf_4
X_5172_ _9599_/Q _5169_/A _8844_/X _5169_/Y VGND VGND VPWR VPWR _9599_/D sky130_fd_sc_hd__a22o_1
XFILLER_122_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput2 debug_oeb VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__clkbuf_4
X_8931_ _9084_/Q _9083_/Q _9051_/Q VGND VGND VPWR VPWR _8931_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_opt_1_0_csclk _9329_/CLK VGND VGND VPWR VPWR clkbuf_leaf_2_csclk/A sky130_fd_sc_hd__clkbuf_16
XFILLER_49_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8862_ _7608_/Y _9639_/Q _8978_/S VGND VGND VPWR VPWR _8862_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8793_ _8793_/A VGND VGND VPWR VPWR _8794_/A sky130_fd_sc_hd__clkbuf_1
X_7813_ _7813_/A VGND VGND VPWR VPWR _8341_/A sky130_fd_sc_hd__clkbuf_16
X_7744_ _9066_/Q _7744_/B VGND VGND VPWR VPWR _7744_/X sky130_fd_sc_hd__and2_1
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4956_ _4994_/A VGND VGND VPWR VPWR _4957_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_165_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7675_ _6498_/Y _7465_/X _6574_/Y _7467_/X VGND VGND VPWR VPWR _7675_/X sky130_fd_sc_hd__o22a_1
X_4887_ _9732_/Q VGND VGND VPWR VPWR _4887_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9414_ _9514_/CLK _9414_/D _9685_/SET_B VGND VGND VPWR VPWR _9414_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6626_ _6621_/Y _4524_/B _8787_/A _5278_/B _6625_/X VGND VGND VPWR VPWR _6627_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_192_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9345_ _9371_/CLK _9345_/D _9295_/SET_B VGND VGND VPWR VPWR _9345_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6557_ _9409_/Q VGND VGND VPWR VPWR _6557_/Y sky130_fd_sc_hd__inv_2
XFILLER_192_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5508_ _5508_/A VGND VGND VPWR VPWR _5509_/A sky130_fd_sc_hd__clkbuf_4
X_9276_ _9596_/CLK _9276_/D _9528_/SET_B VGND VGND VPWR VPWR _9276_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_105_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6488_ _8761_/A _5610_/B _6484_/Y _5594_/B _6487_/X VGND VGND VPWR VPWR _6501_/B
+ sky130_fd_sc_hd__o221a_1
X_5439_ _9418_/Q _5433_/A _8841_/X _5433_/Y VGND VGND VPWR VPWR _9418_/D sky130_fd_sc_hd__a22o_1
XFILLER_160_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput350 _9022_/Q VGND VGND VPWR VPWR wb_dat_o[2] sky130_fd_sc_hd__buf_2
X_8227_ _8595_/B _8227_/B _8571_/B _8499_/B VGND VGND VPWR VPWR _8231_/A sky130_fd_sc_hd__or4_1
XFILLER_126_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8158_ _8158_/A _8630_/B VGND VGND VPWR VPWR _8160_/A sky130_fd_sc_hd__or2_1
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7109_ _7127_/C _7109_/B VGND VGND VPWR VPWR _7110_/A sky130_fd_sc_hd__or2_1
XFILLER_59_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8089_ _8218_/B _7837_/A _8102_/B VGND VGND VPWR VPWR _8120_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4810_ _4891_/A _4931_/B VGND VGND VPWR VPWR _5251_/B sky130_fd_sc_hd__or2_4
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5790_ _5790_/A VGND VGND VPWR VPWR _5791_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_147_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4741_ _4805_/A _4780_/B VGND VGND VPWR VPWR _5818_/B sky130_fd_sc_hd__or2_4
XFILLER_174_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4672_ _4919_/A _4787_/A VGND VGND VPWR VPWR _5526_/B sky130_fd_sc_hd__or2_4
X_7460_ _7462_/A _7474_/C _9255_/Q VGND VGND VPWR VPWR _7461_/A sky130_fd_sc_hd__or3_1
X_6411_ _6411_/A VGND VGND VPWR VPWR _6411_/Y sky130_fd_sc_hd__clkinv_2
X_9130_ _9379_/CLK _9130_/D _9779_/SET_B VGND VGND VPWR VPWR _9130_/Q sky130_fd_sc_hd__dfrtp_1
X_7391_ _6458_/Y _7059_/D _6424_/Y _7116_/X _7390_/X VGND VGND VPWR VPWR _7396_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_155_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6342_ _9725_/Q VGND VGND VPWR VPWR _6342_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_170_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9061_ _4450_/A1 _9061_/D _6146_/A VGND VGND VPWR VPWR _9061_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_103_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6273_ _6268_/Y _4524_/B _6269_/Y _5458_/B _6272_/X VGND VGND VPWR VPWR _6280_/C
+ sky130_fd_sc_hd__o221a_1
X_5224_ _9563_/Q _5218_/Y _8922_/X _5218_/A VGND VGND VPWR VPWR _9563_/D sky130_fd_sc_hd__o22a_1
X_8012_ _8523_/A _8517_/A VGND VGND VPWR VPWR _8013_/B sky130_fd_sc_hd__or2_1
XFILLER_102_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5155_ _9610_/Q _5147_/A _8916_/A1 _5147_/Y VGND VGND VPWR VPWR _9610_/D sky130_fd_sc_hd__a22o_1
XFILLER_69_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5086_ _9655_/Q _5082_/A _8930_/A1 _5082_/Y VGND VGND VPWR VPWR _9655_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8914_ _9625_/Q _8846_/X _8955_/S VGND VGND VPWR VPWR _8914_/X sky130_fd_sc_hd__mux2_1
X_8845_ _9706_/Q _9665_/Q _9587_/Q VGND VGND VPWR VPWR _8845_/X sky130_fd_sc_hd__mux2_8
XFILLER_71_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8776_ _8776_/A VGND VGND VPWR VPWR _8776_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_188_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5988_ _5988_/A VGND VGND VPWR VPWR _5988_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7727_ _9699_/Q VGND VGND VPWR VPWR _7727_/Y sky130_fd_sc_hd__inv_2
X_4939_ _4939_/A VGND VGND VPWR VPWR _4939_/X sky130_fd_sc_hd__clkbuf_1
X_7658_ _6674_/Y _7461_/X _6711_/Y _7463_/X _7657_/X VGND VGND VPWR VPWR _7661_/C
+ sky130_fd_sc_hd__o221a_1
XANTENNA_40 _6111_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_73 _8586_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_51 _6595_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_84 _7019_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_62 _6847_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6609_ _9544_/Q VGND VGND VPWR VPWR _6609_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_192_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7589_ _7589_/A _7589_/B _7589_/C _7589_/D VGND VGND VPWR VPWR _7590_/D sky130_fd_sc_hd__and4_1
XANTENNA_95 input77/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9328_ _9380_/CLK _9328_/D _4628_/A VGND VGND VPWR VPWR _9328_/Q sky130_fd_sc_hd__dfrtp_1
X_9259_ _9601_/CLK _9259_/D _9295_/SET_B VGND VGND VPWR VPWR _9259_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_97_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_44_csclk _9329_/CLK VGND VGND VPWR VPWR _9755_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_97_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6960_ _4936_/Y _6952_/A _9028_/Q _6952_/Y VGND VGND VPWR VPWR _9028_/D sky130_fd_sc_hd__o22a_1
XFILLER_26_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5911_ _9129_/Q _5907_/A _8925_/A1 _5907_/Y VGND VGND VPWR VPWR _9129_/D sky130_fd_sc_hd__a22o_1
X_6891_ _9257_/Q VGND VGND VPWR VPWR _6891_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_81_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5842_ _9182_/Q _5839_/A _8844_/X _5839_/Y VGND VGND VPWR VPWR _9182_/D sky130_fd_sc_hd__a22o_1
X_8630_ _8630_/A _8630_/B _8630_/C _8630_/D VGND VGND VPWR VPWR _8709_/C sky130_fd_sc_hd__or4_2
XFILLER_61_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8561_ _8624_/B _8632_/B VGND VGND VPWR VPWR _8713_/B sky130_fd_sc_hd__nor2_1
X_5773_ _9228_/Q _5770_/A _5965_/B1 _5770_/Y VGND VGND VPWR VPWR _9228_/D sky130_fd_sc_hd__a22o_1
X_7512_ _6644_/Y _7451_/X _6713_/Y _7453_/X _7511_/X VGND VGND VPWR VPWR _7517_/B
+ sky130_fd_sc_hd__o221a_1
X_4724_ _4720_/Y _5679_/B _4722_/Y _5768_/B VGND VGND VPWR VPWR _4724_/X sky130_fd_sc_hd__o22a_1
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8492_ _8492_/A VGND VGND VPWR VPWR _8614_/A sky130_fd_sc_hd__inv_2
XFILLER_190_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7443_ _7443_/A VGND VGND VPWR VPWR _7443_/X sky130_fd_sc_hd__buf_8
X_4655_ _9712_/Q _4636_/A _8952_/X _4636_/Y VGND VGND VPWR VPWR _9712_/D sky130_fd_sc_hd__a22o_1
Xinput60 mgmt_gpio_in[31] VGND VGND VPWR VPWR _6132_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_128_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput82 spi_sdoenb VGND VGND VPWR VPWR input82/X sky130_fd_sc_hd__buf_4
X_7374_ _7374_/A _7374_/B _7374_/C _7374_/D VGND VGND VPWR VPWR _7375_/C sky130_fd_sc_hd__and4_1
Xinput71 mgmt_gpio_in[8] VGND VGND VPWR VPWR _4737_/A sky130_fd_sc_hd__clkbuf_2
X_4586_ _9741_/Q _4579_/A _5966_/B1 _4579_/Y VGND VGND VPWR VPWR _9741_/D sky130_fd_sc_hd__a22o_1
X_6325_ _6325_/A _6325_/B _6325_/C VGND VGND VPWR VPWR _6326_/D sky130_fd_sc_hd__and3_2
X_9113_ _9378_/CLK _9113_/D _9646_/SET_B VGND VGND VPWR VPWR _9113_/Q sky130_fd_sc_hd__dfrtp_1
Xinput93 sram_ro_data[0] VGND VGND VPWR VPWR _4860_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_143_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9044_ _9790_/CLK _9044_/D VGND VGND VPWR VPWR _9044_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6256_ _9473_/Q VGND VGND VPWR VPWR _6256_/Y sky130_fd_sc_hd__inv_4
XFILLER_130_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5207_ _9574_/Q _5203_/Y _8906_/X _5203_/A VGND VGND VPWR VPWR _9574_/D sky130_fd_sc_hd__o22a_1
XFILLER_130_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6187_ _6187_/A _6187_/B _6187_/C VGND VGND VPWR VPWR _6237_/B sky130_fd_sc_hd__and3_1
XFILLER_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5138_ _9624_/Q _5136_/A _8845_/X _5136_/Y VGND VGND VPWR VPWR _9624_/D sky130_fd_sc_hd__a22o_1
XFILLER_123_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5069_ _5069_/A VGND VGND VPWR VPWR _9664_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8828_ _9591_/Q input81/X _8833_/S VGND VGND VPWR VPWR _8828_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8759_ _8759_/A VGND VGND VPWR VPWR _8760_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_12_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6110_ _9509_/Q VGND VGND VPWR VPWR _6110_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7090_ _4720_/Y _7077_/C _4751_/Y _7077_/D _7089_/X VGND VGND VPWR VPWR _7090_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6041_ _6041_/A VGND VGND VPWR VPWR _6041_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7992_ _8116_/A _7992_/B VGND VGND VPWR VPWR _7993_/A sky130_fd_sc_hd__or2_1
XFILLER_93_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6943_ _6938_/Y _5594_/B _6939_/Y _5757_/B _6942_/X VGND VGND VPWR VPWR _6944_/C
+ sky130_fd_sc_hd__o221a_1
X_9731_ _9774_/CLK _9731_/D _7011_/B VGND VGND VPWR VPWR _9731_/Q sky130_fd_sc_hd__dfrtp_1
X_9662_ _9664_/CLK _9662_/D _6146_/A VGND VGND VPWR VPWR _9662_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_81_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6874_ _9516_/Q VGND VGND VPWR VPWR _6874_/Y sky130_fd_sc_hd__inv_2
X_8613_ _8666_/C _8613_/B _8666_/D VGND VGND VPWR VPWR _8616_/B sky130_fd_sc_hd__or3_1
X_5825_ _9193_/Q _5820_/A _8929_/A1 _5820_/Y VGND VGND VPWR VPWR _9193_/D sky130_fd_sc_hd__a22o_1
XFILLER_22_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9593_ _9601_/CLK _9593_/D _9295_/SET_B VGND VGND VPWR VPWR _9593_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8544_ _8544_/A _8544_/B _8544_/C VGND VGND VPWR VPWR _8625_/B sky130_fd_sc_hd__or3_2
X_5756_ _5713_/Y _5750_/Y _5755_/Y _9239_/Q _5755_/A VGND VGND VPWR VPWR _9239_/D
+ sky130_fd_sc_hd__a32o_1
X_5687_ _9258_/Q _5681_/A _8955_/A1 _5681_/Y VGND VGND VPWR VPWR _9258_/D sky130_fd_sc_hd__a22o_1
X_8475_ _8703_/C _8617_/A _8475_/C VGND VGND VPWR VPWR _8477_/A sky130_fd_sc_hd__or3_1
X_4707_ _4925_/A _4780_/B VGND VGND VPWR VPWR _5671_/B sky130_fd_sc_hd__or2_4
X_7426_ _7472_/A _7476_/C _7474_/D VGND VGND VPWR VPWR _7427_/A sky130_fd_sc_hd__or3_1
X_4638_ _4994_/A VGND VGND VPWR VPWR _4639_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_162_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4569_ _9753_/Q _4566_/A _8844_/X _4566_/Y VGND VGND VPWR VPWR _9753_/D sky130_fd_sc_hd__a22o_1
X_7357_ _6533_/Y _7040_/C _6479_/Y _7059_/C VGND VGND VPWR VPWR _7357_/X sky130_fd_sc_hd__o22a_1
X_6308_ _9236_/Q VGND VGND VPWR VPWR _6308_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_143_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7288_ _4899_/Y _7086_/X _4848_/Y _7088_/X VGND VGND VPWR VPWR _7288_/X sky130_fd_sc_hd__o22a_1
X_6239_ _9429_/Q VGND VGND VPWR VPWR _6239_/Y sky130_fd_sc_hd__inv_2
X_9027_ _9027_/CLK _9027_/D VGND VGND VPWR VPWR _9027_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5610_ _6052_/A _5610_/B VGND VGND VPWR VPWR _5611_/A sky130_fd_sc_hd__or2_1
X_6590_ _8777_/A _5306_/B _6589_/Y _5366_/B VGND VGND VPWR VPWR _6590_/X sky130_fd_sc_hd__o22a_2
XFILLER_157_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5541_ _9349_/Q _5536_/A _8929_/A1 _5536_/Y VGND VGND VPWR VPWR _9349_/D sky130_fd_sc_hd__a22o_1
XFILLER_145_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8260_ _8260_/A _8260_/B VGND VGND VPWR VPWR _8578_/B sky130_fd_sc_hd__nor2_1
X_5472_ _9397_/Q _5471_/A _8846_/X _5471_/Y VGND VGND VPWR VPWR _9397_/D sky130_fd_sc_hd__a22o_1
X_7211_ _7211_/A _7211_/B _7211_/C _7211_/D VGND VGND VPWR VPWR _7221_/B sky130_fd_sc_hd__and4_1
X_8191_ _8345_/A VGND VGND VPWR VPWR _8583_/B sky130_fd_sc_hd__inv_2
XFILLER_172_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7142_ _6914_/Y _7059_/B _6905_/Y _7068_/C _7141_/X VGND VGND VPWR VPWR _7145_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_113_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7073_ _7098_/C _7127_/A _7073_/C VGND VGND VPWR VPWR _7074_/A sky130_fd_sc_hd__or3_1
XFILLER_98_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6024_ _9709_/Q _6023_/Y _9080_/Q _6023_/A VGND VGND VPWR VPWR _9080_/D sky130_fd_sc_hd__a22o_1
XFILLER_39_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7975_ _7975_/A VGND VGND VPWR VPWR _8389_/A sky130_fd_sc_hd__buf_8
X_6926_ _9270_/Q VGND VGND VPWR VPWR _6926_/Y sky130_fd_sc_hd__inv_2
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9714_ _9089_/CLK _9714_/D _4648_/X VGND VGND VPWR VPWR _9714_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_14_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6857_ _6855_/Y _5420_/B _6856_/Y _5374_/B VGND VGND VPWR VPWR _6857_/X sky130_fd_sc_hd__o22a_1
XFILLER_120_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9645_ _9774_/CLK _9645_/D _7011_/B VGND VGND VPWR VPWR _9645_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_167_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9576_ _9788_/CLK _9576_/D _9646_/SET_B VGND VGND VPWR VPWR _9576_/Q sky130_fd_sc_hd__dfrtp_1
X_6788_ _9529_/Q VGND VGND VPWR VPWR _6788_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5808_ _9056_/Q _5691_/A _5643_/Y _5753_/B _9203_/Q VGND VGND VPWR VPWR _5808_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_136_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8527_ _8612_/B _8527_/B _8527_/C _8666_/A VGND VGND VPWR VPWR _8531_/B sky130_fd_sc_hd__or4_1
X_5739_ _9055_/Q _7125_/A _7127_/A _5737_/A _5713_/Y VGND VGND VPWR VPWR _5740_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_135_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8458_ _7864_/X _8319_/A _8097_/B _8550_/A VGND VGND VPWR VPWR _8614_/C sky130_fd_sc_hd__o22ai_1
XFILLER_151_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8389_ _8389_/A VGND VGND VPWR VPWR _8518_/B sky130_fd_sc_hd__inv_2
X_7409_ _7456_/A _7472_/A _9255_/Q VGND VGND VPWR VPWR _7410_/A sky130_fd_sc_hd__or3_1
XFILLER_104_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4972_ _4972_/A VGND VGND VPWR VPWR _4972_/X sky130_fd_sc_hd__clkbuf_1
X_7760_ _8394_/D VGND VGND VPWR VPWR _7836_/A sky130_fd_sc_hd__inv_2
XFILLER_91_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7691_ _6363_/Y _7455_/X _6445_/Y _7457_/X VGND VGND VPWR VPWR _7691_/X sky130_fd_sc_hd__o22a_1
X_6711_ _9538_/Q VGND VGND VPWR VPWR _6711_/Y sky130_fd_sc_hd__clkinv_4
X_9430_ _9508_/CLK _9430_/D _9295_/SET_B VGND VGND VPWR VPWR _9430_/Q sky130_fd_sc_hd__dfrtp_1
X_6642_ _6637_/Y _5797_/B _6638_/Y _5768_/B _6641_/X VGND VGND VPWR VPWR _6649_/B
+ sky130_fd_sc_hd__o221a_1
X_9361_ _9545_/CLK _9361_/D _4628_/A VGND VGND VPWR VPWR _9361_/Q sky130_fd_sc_hd__dfstp_1
X_8312_ _8310_/X _8676_/B _8592_/A _8312_/D VGND VGND VPWR VPWR _8312_/X sky130_fd_sc_hd__and4bb_1
XFILLER_118_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6573_ _8789_/A _5317_/B _6569_/Y _4590_/B _6572_/X VGND VGND VPWR VPWR _6586_/A
+ sky130_fd_sc_hd__o221a_1
X_9292_ _9596_/CLK _9292_/D _9528_/SET_B VGND VGND VPWR VPWR _9292_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_1_1_0_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR clkbuf_1_1_1_mgmt_gpio_in[4]/A
+ sky130_fd_sc_hd__clkbuf_2
X_5524_ _9360_/Q _5520_/A _5966_/B1 _5520_/Y VGND VGND VPWR VPWR _9360_/D sky130_fd_sc_hd__a22o_1
XFILLER_133_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5455_ _9408_/Q _5452_/A _5965_/B1 _5452_/Y VGND VGND VPWR VPWR _9408_/D sky130_fd_sc_hd__a22o_1
X_8243_ _8243_/A VGND VGND VPWR VPWR _8362_/B sky130_fd_sc_hd__inv_2
X_8174_ _8376_/A _8174_/B VGND VGND VPWR VPWR _8175_/B sky130_fd_sc_hd__nor2_1
XFILLER_132_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5386_ _9456_/Q _5384_/A _8845_/X _5384_/Y VGND VGND VPWR VPWR _9456_/D sky130_fd_sc_hd__a22o_1
XFILLER_132_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7125_ _7125_/A _7127_/B _7127_/C VGND VGND VPWR VPWR _7126_/A sky130_fd_sc_hd__or3_1
XFILLER_113_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7056_ _9248_/Q _7056_/B _9246_/Q _9245_/Q VGND VGND VPWR VPWR _7087_/B sky130_fd_sc_hd__or4_1
X_6007_ _6007_/A VGND VGND VPWR VPWR _6007_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_55_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7958_ _8189_/A _8099_/B VGND VGND VPWR VPWR _7966_/B sky130_fd_sc_hd__or2_1
XFILLER_131_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6909_ _9160_/Q VGND VGND VPWR VPWR _6909_/Y sky130_fd_sc_hd__clkinv_4
X_7889_ _8525_/A _8189_/A _7903_/C _8193_/A VGND VGND VPWR VPWR _7890_/A sky130_fd_sc_hd__or4_1
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9628_ _9639_/CLK _9628_/D _9757_/SET_B VGND VGND VPWR VPWR _9628_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9559_ _9776_/CLK _9559_/D _4628_/A VGND VGND VPWR VPWR _9559_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_183_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_152 _7879_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_130 _7331_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_141 _5045_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_185 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_174 _8803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_163 _9080_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_196 _6586_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5240_ _5545_/A _5240_/B VGND VGND VPWR VPWR _5241_/A sky130_fd_sc_hd__or2_1
XFILLER_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5171_ _9600_/Q _5169_/A _8845_/X _5169_/Y VGND VGND VPWR VPWR _9600_/D sky130_fd_sc_hd__a22o_1
XFILLER_96_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8930_ _9611_/Q _8930_/A1 _8930_/S VGND VGND VPWR VPWR _8930_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput3 debug_out VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__buf_4
X_8861_ _8860_/X _9169_/Q _9054_/Q VGND VGND VPWR VPWR _8861_/X sky130_fd_sc_hd__mux2_1
X_8792_ _8792_/A VGND VGND VPWR VPWR _8792_/X sky130_fd_sc_hd__clkbuf_1
X_7812_ _8379_/D _8379_/B _7838_/B VGND VGND VPWR VPWR _7813_/A sky130_fd_sc_hd__or3_1
XFILLER_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7743_ _9068_/Q _7743_/A2 _9067_/Q _7743_/B2 _7742_/X VGND VGND VPWR VPWR _7743_/X
+ sky130_fd_sc_hd__a221o_1
X_4955_ _4949_/Y _4951_/Y _4952_/Y _4954_/X VGND VGND VPWR VPWR _9709_/D sky130_fd_sc_hd__o22ai_1
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7674_ _6504_/Y _7451_/X _6556_/Y _7453_/X _7673_/X VGND VGND VPWR VPWR _7679_/B
+ sky130_fd_sc_hd__o221a_1
X_4886_ _4882_/Y _4504_/B _4883_/Y _5259_/B _4885_/X VGND VGND VPWR VPWR _4896_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_192_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9413_ _9514_/CLK _9413_/D _9685_/SET_B VGND VGND VPWR VPWR _9413_/Q sky130_fd_sc_hd__dfstp_1
X_6625_ _8781_/A _4491_/B _6624_/Y _4822_/X VGND VGND VPWR VPWR _6625_/X sky130_fd_sc_hd__o22a_1
XFILLER_165_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9344_ _9344_/CLK _9344_/D _9295_/SET_B VGND VGND VPWR VPWR _9344_/Q sky130_fd_sc_hd__dfrtp_1
X_6556_ _9440_/Q VGND VGND VPWR VPWR _6556_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_20_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9275_ _9371_/CLK _9275_/D _9295_/SET_B VGND VGND VPWR VPWR _9275_/Q sky130_fd_sc_hd__dfrtp_1
X_5507_ _5545_/A _5507_/B VGND VGND VPWR VPWR _5508_/A sky130_fd_sc_hd__or2_1
X_6487_ _6485_/Y _5583_/B _6486_/Y _5864_/B VGND VGND VPWR VPWR _6487_/X sky130_fd_sc_hd__o22a_1
X_8226_ _8341_/A _8305_/B _8226_/C VGND VGND VPWR VPWR _8499_/B sky130_fd_sc_hd__nor3_1
X_5438_ _9419_/Q _5433_/A _8842_/X _5433_/Y VGND VGND VPWR VPWR _9419_/D sky130_fd_sc_hd__a22o_1
Xoutput351 _9042_/Q VGND VGND VPWR VPWR wb_dat_o[30] sky130_fd_sc_hd__buf_2
XFILLER_160_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput340 _9032_/Q VGND VGND VPWR VPWR wb_dat_o[20] sky130_fd_sc_hd__buf_2
XFILLER_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8157_ _8164_/A _8554_/A VGND VGND VPWR VPWR _8630_/B sky130_fd_sc_hd__nor2_1
X_5369_ _9467_/Q _5368_/A _5963_/B1 _5368_/Y VGND VGND VPWR VPWR _9467_/D sky130_fd_sc_hd__a22o_1
X_8088_ _8188_/B _8389_/A VGND VGND VPWR VPWR _8433_/B sky130_fd_sc_hd__nor2_1
X_7108_ _7108_/A _7108_/B _7108_/C _7108_/D VGND VGND VPWR VPWR _7132_/B sky130_fd_sc_hd__and4_1
XFILLER_101_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7039_ _7039_/A VGND VGND VPWR VPWR _7040_/D sky130_fd_sc_hd__clkbuf_16
XFILLER_59_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4740_ _9190_/Q VGND VGND VPWR VPWR _4740_/Y sky130_fd_sc_hd__clkinv_2
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4671_ _9354_/Q VGND VGND VPWR VPWR _4671_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6410_ _9316_/Q VGND VGND VPWR VPWR _6410_/Y sky130_fd_sc_hd__clkinv_2
X_7390_ _6330_/Y _7118_/X _6335_/Y _7048_/C VGND VGND VPWR VPWR _7390_/X sky130_fd_sc_hd__o22a_1
XFILLER_174_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6341_ _9545_/Q VGND VGND VPWR VPWR _6341_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_155_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9060_ _4450_/A1 _9060_/D _6146_/A VGND VGND VPWR VPWR _9065_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_142_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6272_ _6270_/Y _4861_/X _6271_/Y _5278_/B VGND VGND VPWR VPWR _6272_/X sky130_fd_sc_hd__o22a_1
X_5223_ _9564_/Q _5218_/Y _8926_/X _5218_/A VGND VGND VPWR VPWR _9564_/D sky130_fd_sc_hd__o22a_1
XFILLER_170_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8011_ _8583_/A _8538_/B _8525_/C VGND VGND VPWR VPWR _8523_/A sky130_fd_sc_hd__or3_2
XFILLER_130_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5154_ _9611_/Q _5147_/A _8930_/A1 _5147_/Y VGND VGND VPWR VPWR _9611_/D sky130_fd_sc_hd__a22o_1
XFILLER_69_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5085_ _9656_/Q _5082_/A _5965_/B1 _5082_/Y VGND VGND VPWR VPWR _9656_/D sky130_fd_sc_hd__a22o_1
XFILLER_112_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8913_ _7723_/X _9087_/Q _9051_/Q VGND VGND VPWR VPWR _8913_/X sky130_fd_sc_hd__mux2_1
X_8844_ _9705_/Q _9664_/Q _9587_/Q VGND VGND VPWR VPWR _8844_/X sky130_fd_sc_hd__mux2_8
XFILLER_64_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8775_ _8775_/A VGND VGND VPWR VPWR _8776_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_169_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5987_ _6040_/A VGND VGND VPWR VPWR _5988_/A sky130_fd_sc_hd__clkbuf_1
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7726_ _9698_/Q VGND VGND VPWR VPWR _7726_/Y sky130_fd_sc_hd__clkinv_4
X_4938_ _4994_/A VGND VGND VPWR VPWR _4939_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_138_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_41 _6117_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7657_ _6646_/Y _7465_/X _6730_/Y _7467_/X VGND VGND VPWR VPWR _7657_/X sky130_fd_sc_hd__o22a_1
X_4869_ input4/X VGND VGND VPWR VPWR _4869_/Y sky130_fd_sc_hd__inv_2
XANTENNA_30 _4858_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_74 _8586_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_52 _6651_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_63 _6877_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6608_ _8775_/A _5344_/B _6604_/Y _5328_/B _6607_/X VGND VGND VPWR VPWR _6627_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_20_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_85 _7019_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_96 input78/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7588_ _6212_/Y _7471_/X _7260_/A _7473_/X _7587_/X VGND VGND VPWR VPWR _7589_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_192_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9327_ _9352_/CLK _9327_/D _9646_/SET_B VGND VGND VPWR VPWR _9327_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6539_ _9117_/Q VGND VGND VPWR VPWR _6539_/Y sky130_fd_sc_hd__inv_2
X_9258_ _9601_/CLK _9258_/D _9295_/SET_B VGND VGND VPWR VPWR _9258_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8209_ _8660_/A _8226_/C VGND VGND VPWR VPWR _8210_/A sky130_fd_sc_hd__or2_1
X_9189_ _9655_/CLK _9189_/D _9633_/SET_B VGND VGND VPWR VPWR _9189_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_153_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5910_ _9130_/Q _5907_/A _8844_/X _5907_/Y VGND VGND VPWR VPWR _9130_/D sky130_fd_sc_hd__a22o_1
XFILLER_19_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6890_ _9219_/Q VGND VGND VPWR VPWR _6890_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5841_ _9183_/Q _5839_/A _8845_/X _5839_/Y VGND VGND VPWR VPWR _9183_/D sky130_fd_sc_hd__a22o_1
XFILLER_34_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8560_ _8560_/A _8560_/B VGND VGND VPWR VPWR _8713_/D sky130_fd_sc_hd__or2_2
X_5772_ _9229_/Q _5770_/A _5964_/B1 _5770_/Y VGND VGND VPWR VPWR _9229_/D sky130_fd_sc_hd__a22o_1
XFILLER_61_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7511_ _6737_/Y _7455_/X _6773_/Y _7457_/X VGND VGND VPWR VPWR _7511_/X sky130_fd_sc_hd__o22a_1
X_4723_ _6111_/B _4780_/B VGND VGND VPWR VPWR _5768_/B sky130_fd_sc_hd__or2_4
X_8491_ _7862_/Y _8302_/Y _8667_/A _8369_/B VGND VGND VPWR VPWR _8599_/D sky130_fd_sc_hd__a211o_1
XFILLER_187_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7442_ _7476_/A _9251_/Q _7476_/C _7474_/D VGND VGND VPWR VPWR _7443_/A sky130_fd_sc_hd__or4_1
X_4654_ _4654_/A VGND VGND VPWR VPWR _4654_/X sky130_fd_sc_hd__clkbuf_1
Xinput61 mgmt_gpio_in[32] VGND VGND VPWR VPWR input61/X sky130_fd_sc_hd__clkbuf_4
Xinput50 mgmt_gpio_in[22] VGND VGND VPWR VPWR input50/X sky130_fd_sc_hd__clkbuf_4
XFILLER_174_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput72 mgmt_gpio_in[9] VGND VGND VPWR VPWR _6941_/A sky130_fd_sc_hd__clkbuf_1
X_4585_ _9742_/Q _4579_/A _5965_/B1 _4579_/Y VGND VGND VPWR VPWR _9742_/D sky130_fd_sc_hd__a22o_1
X_7373_ _6587_/Y _7124_/X _6480_/Y _7068_/B _7372_/X VGND VGND VPWR VPWR _7374_/D
+ sky130_fd_sc_hd__o221a_1
Xinput83 spimemio_flash_clk VGND VGND VPWR VPWR input83/X sky130_fd_sc_hd__buf_6
X_6324_ _6320_/Y _5572_/B _6321_/Y _5507_/B _6323_/Y VGND VGND VPWR VPWR _6325_/C
+ sky130_fd_sc_hd__o221a_1
X_9112_ _9379_/CLK _9112_/D _9779_/SET_B VGND VGND VPWR VPWR _9112_/Q sky130_fd_sc_hd__dfrtp_1
Xinput94 sram_ro_data[10] VGND VGND VPWR VPWR _6778_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_9043_ _9664_/CLK _9043_/D VGND VGND VPWR VPWR _9043_/Q sky130_fd_sc_hd__dfxtp_1
X_6255_ _6239_/Y _5420_/B _6242_/X _6248_/X _6254_/X VGND VGND VPWR VPWR _6326_/A
+ sky130_fd_sc_hd__o2111a_1
X_5206_ _9575_/Q _5203_/Y _8928_/X _5203_/A VGND VGND VPWR VPWR _9575_/D sky130_fd_sc_hd__o22a_1
XFILLER_115_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6186_ _7260_/A _5610_/B _6182_/Y _5776_/B _6185_/X VGND VGND VPWR VPWR _6187_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_130_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5137_ _9625_/Q _5136_/A _8846_/X _5136_/Y VGND VGND VPWR VPWR _9625_/D sky130_fd_sc_hd__a22o_1
X_5068_ _8966_/X _9664_/Q _5078_/S VGND VGND VPWR VPWR _5069_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8827_ _8826_/X _7020_/B _9586_/Q VGND VGND VPWR VPWR _8827_/X sky130_fd_sc_hd__mux2_4
X_8758_ _8758_/A VGND VGND VPWR VPWR _8758_/X sky130_fd_sc_hd__clkbuf_1
X_7709_ _9083_/Q _9082_/Q VGND VGND VPWR VPWR _7711_/A sky130_fd_sc_hd__nand2_1
X_8689_ _8689_/A _8709_/D _8713_/C _8714_/D VGND VGND VPWR VPWR _8689_/X sky130_fd_sc_hd__or4_1
XFILLER_193_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ _6040_/A VGND VGND VPWR VPWR _6041_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_66_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7991_ _7991_/A VGND VGND VPWR VPWR _8550_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_93_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6942_ _6940_/Y _5080_/B _6941_/Y _6134_/A VGND VGND VPWR VPWR _6942_/X sky130_fd_sc_hd__o22a_1
X_9730_ _9774_/CLK _9730_/D _7011_/B VGND VGND VPWR VPWR _9730_/Q sky130_fd_sc_hd__dfstp_2
X_9661_ _9664_/CLK _9661_/D _6146_/A VGND VGND VPWR VPWR _9661_/Q sky130_fd_sc_hd__dfrtp_1
X_6873_ _9438_/Q VGND VGND VPWR VPWR _6873_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_179_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8612_ _8612_/A _8612_/B VGND VGND VPWR VPWR _8666_/D sky130_fd_sc_hd__or2_1
X_5824_ _9194_/Q _5820_/A _8925_/A1 _5820_/Y VGND VGND VPWR VPWR _9194_/D sky130_fd_sc_hd__a22o_1
X_9592_ _9617_/CLK _9592_/D _9295_/SET_B VGND VGND VPWR VPWR _9592_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8543_ _8543_/A VGND VGND VPWR VPWR _8543_/Y sky130_fd_sc_hd__inv_2
X_5755_ _5755_/A VGND VGND VPWR VPWR _5755_/Y sky130_fd_sc_hd__inv_2
X_5686_ _9259_/Q _5681_/A _8842_/X _5681_/Y VGND VGND VPWR VPWR _9259_/D sky130_fd_sc_hd__a22o_1
XFILLER_147_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4706_ _9264_/Q VGND VGND VPWR VPWR _4706_/Y sky130_fd_sc_hd__clkinv_2
X_8474_ _8474_/A _8474_/B VGND VGND VPWR VPWR _8475_/C sky130_fd_sc_hd__or2_1
XFILLER_190_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4637_ _9718_/Q _4636_/A _8953_/X _4636_/Y VGND VGND VPWR VPWR _9718_/D sky130_fd_sc_hd__a22o_1
X_7425_ _7425_/A VGND VGND VPWR VPWR _7425_/X sky130_fd_sc_hd__buf_8
XFILLER_162_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7356_ _6574_/Y _7082_/X _6615_/Y _7084_/X _7355_/X VGND VGND VPWR VPWR _7375_/A
+ sky130_fd_sc_hd__o221a_1
X_4568_ _9754_/Q _4566_/A _8845_/X _4566_/Y VGND VGND VPWR VPWR _9754_/D sky130_fd_sc_hd__a22o_1
X_7287_ _7287_/A _7287_/B _7287_/C VGND VGND VPWR VPWR _7287_/Y sky130_fd_sc_hd__nand3_4
XFILLER_116_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6307_ _6307_/A _6307_/B _6307_/C _6307_/D VGND VGND VPWR VPWR _6326_/C sky130_fd_sc_hd__and4_1
XFILLER_89_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4499_ _9780_/Q _4493_/A _5965_/B1 _4493_/Y VGND VGND VPWR VPWR _9780_/D sky130_fd_sc_hd__a22o_1
X_6238_ _6149_/A _6237_/Y _9042_/Q _6149_/Y VGND VGND VPWR VPWR _9042_/D sky130_fd_sc_hd__o22a_1
XFILLER_134_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9026_ _9027_/CLK _9026_/D VGND VGND VPWR VPWR _9026_/Q sky130_fd_sc_hd__dfxtp_1
X_6169_ _9508_/Q VGND VGND VPWR VPWR _6169_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_43_csclk _9329_/CLK VGND VGND VPWR VPWR _9758_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_13_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5540_ _9350_/Q _5536_/A _8925_/A1 _5536_/Y VGND VGND VPWR VPWR _9350_/D sky130_fd_sc_hd__a22o_1
X_5471_ _5471_/A VGND VGND VPWR VPWR _5471_/Y sky130_fd_sc_hd__inv_2
XFILLER_157_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7210_ _6367_/Y _7048_/D _6439_/Y _7040_/B _7209_/X VGND VGND VPWR VPWR _7211_/D
+ sky130_fd_sc_hd__o221a_1
X_8190_ _8189_/A _8213_/A _8189_/Y VGND VGND VPWR VPWR _8345_/A sky130_fd_sc_hd__a21oi_1
X_7141_ _6819_/Y _7079_/B _6926_/Y _7059_/A VGND VGND VPWR VPWR _7141_/X sky130_fd_sc_hd__o22a_1
XFILLER_125_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7072_ _7072_/A VGND VGND VPWR VPWR _7077_/B sky130_fd_sc_hd__buf_8
XFILLER_98_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6023_ _6023_/A VGND VGND VPWR VPWR _6023_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7974_ _8379_/B _8093_/A VGND VGND VPWR VPWR _7975_/A sky130_fd_sc_hd__or2_1
XFILLER_27_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6925_ _6925_/A _6925_/B _6925_/C _6925_/D VGND VGND VPWR VPWR _6945_/B sky130_fd_sc_hd__and4_1
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9713_ _9089_/CLK _9713_/D _4651_/X VGND VGND VPWR VPWR _9713_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_120_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6856_ _9459_/Q VGND VGND VPWR VPWR _6856_/Y sky130_fd_sc_hd__clkinv_2
X_9644_ _9776_/CLK _9644_/D _4628_/A VGND VGND VPWR VPWR _9644_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_50_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6787_ _9469_/Q VGND VGND VPWR VPWR _6787_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_167_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5807_ _9204_/Q _5799_/A _8916_/A1 _5799_/Y VGND VGND VPWR VPWR _9204_/D sky130_fd_sc_hd__a22o_1
X_9575_ _9613_/CLK _9575_/D _9646_/SET_B VGND VGND VPWR VPWR _9575_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8526_ _8525_/Y _8517_/Y _8518_/X _8449_/A VGND VGND VPWR VPWR _8666_/A sky130_fd_sc_hd__a31o_1
X_5738_ _9246_/Q _5738_/B VGND VGND VPWR VPWR _7127_/A sky130_fd_sc_hd__or2_2
XFILLER_182_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5669_ _9270_/Q _5662_/A _8840_/X _5662_/Y VGND VGND VPWR VPWR _9270_/D sky130_fd_sc_hd__a22o_1
XFILLER_163_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8457_ _8521_/B _8246_/B _8029_/X VGND VGND VPWR VPWR _8459_/C sky130_fd_sc_hd__o21ai_2
XFILLER_190_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8388_ _8098_/B _8397_/B _8171_/X VGND VGND VPWR VPWR _8631_/A sky130_fd_sc_hd__o21ai_1
X_7408_ _7408_/A VGND VGND VPWR VPWR _7408_/X sky130_fd_sc_hd__buf_6
XFILLER_2_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7339_ _6657_/Y _7079_/B _6634_/Y _7059_/A VGND VGND VPWR VPWR _7339_/X sky130_fd_sc_hd__o22a_1
XFILLER_89_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9009_ _9009_/A _8795_/A VGND VGND VPWR VPWR mgmt_gpio_out[32] sky130_fd_sc_hd__ebufn_8
XFILLER_131_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_1_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_110_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4971_ _4994_/A VGND VGND VPWR VPWR _4972_/A sky130_fd_sc_hd__clkbuf_1
X_6710_ _9426_/Q VGND VGND VPWR VPWR _6710_/Y sky130_fd_sc_hd__inv_2
X_7690_ _6374_/Y _7441_/X _6387_/Y _7443_/X _7689_/X VGND VGND VPWR VPWR _7697_/A
+ sky130_fd_sc_hd__o221a_1
X_6641_ _6639_/Y _5776_/B _6640_/Y _5789_/B VGND VGND VPWR VPWR _6641_/X sky130_fd_sc_hd__o22a_1
XFILLER_32_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9360_ _9771_/CLK _9360_/D _4628_/A VGND VGND VPWR VPWR _9360_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8311_ _8640_/A _8311_/B VGND VGND VPWR VPWR _8592_/A sky130_fd_sc_hd__or2_2
XFILLER_157_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6572_ _6570_/Y _4907_/X _8773_/A _5382_/B VGND VGND VPWR VPWR _6572_/X sky130_fd_sc_hd__o22a_1
X_9291_ _9596_/CLK _9291_/D _9528_/SET_B VGND VGND VPWR VPWR _9291_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_157_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5523_ _9361_/Q _5520_/A _5965_/B1 _5520_/Y VGND VGND VPWR VPWR _9361_/D sky130_fd_sc_hd__a22o_1
XFILLER_172_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5454_ _9409_/Q _5452_/A _5964_/B1 _5452_/Y VGND VGND VPWR VPWR _9409_/D sky130_fd_sc_hd__a22o_1
X_8242_ _8510_/A _8246_/B VGND VGND VPWR VPWR _8243_/A sky130_fd_sc_hd__or2_1
X_5385_ _9457_/Q _5384_/A _8846_/X _5384_/Y VGND VGND VPWR VPWR _9457_/D sky130_fd_sc_hd__a22o_1
XFILLER_132_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8173_ _8688_/A _8173_/B VGND VGND VPWR VPWR _8174_/B sky130_fd_sc_hd__or2_1
XFILLER_105_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7124_ _7124_/A VGND VGND VPWR VPWR _7124_/X sky130_fd_sc_hd__buf_8
XFILLER_59_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7055_ _7055_/A VGND VGND VPWR VPWR _7059_/C sky130_fd_sc_hd__buf_6
X_6006_ _6040_/A VGND VGND VPWR VPWR _6007_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7957_ _8583_/A _8189_/A _8099_/B VGND VGND VPWR VPWR _8195_/B sky130_fd_sc_hd__or3_1
XFILLER_82_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6908_ _9647_/Q VGND VGND VPWR VPWR _6908_/Y sky130_fd_sc_hd__inv_2
X_7888_ _8496_/A _8521_/B VGND VGND VPWR VPWR _7896_/A sky130_fd_sc_hd__or2_1
XFILLER_168_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6839_ _9757_/Q VGND VGND VPWR VPWR _6839_/Y sky130_fd_sc_hd__inv_2
X_9627_ _9757_/CLK _9627_/D _9757_/SET_B VGND VGND VPWR VPWR _9627_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9558_ _9758_/CLK _9558_/D _9633_/SET_B VGND VGND VPWR VPWR _9558_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_136_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8509_ _8509_/A _8693_/A _8600_/B _8662_/B VGND VGND VPWR VPWR _8512_/B sky130_fd_sc_hd__or4_1
X_9489_ _9493_/CLK _9489_/D _4628_/A VGND VGND VPWR VPWR _9489_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_6_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_120 _8816_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_142 _4814_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_131 _7375_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_153 _7992_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_175 _4629_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_164 _9571_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_186 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_197 _8801_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5170_ _9601_/Q _5169_/A _8846_/X _5169_/Y VGND VGND VPWR VPWR _9601_/D sky130_fd_sc_hd__a22o_1
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput4 mask_rev_in[0] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8860_ _7590_/Y _9638_/Q _8978_/S VGND VGND VPWR VPWR _8860_/X sky130_fd_sc_hd__mux2_1
X_8791_ _8791_/A VGND VGND VPWR VPWR _8792_/A sky130_fd_sc_hd__clkbuf_1
X_7811_ _7811_/A VGND VGND VPWR VPWR _8202_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_51_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7742_ _9066_/Q _7742_/B VGND VGND VPWR VPWR _7742_/X sky130_fd_sc_hd__and2_1
X_4954_ _4953_/Y _7008_/A _9092_/Q _9048_/Q _9091_/Q VGND VGND VPWR VPWR _4954_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7673_ _6508_/Y _7455_/X _6551_/Y _7457_/X VGND VGND VPWR VPWR _7673_/X sky130_fd_sc_hd__o22a_1
X_9412_ _9493_/CLK _9412_/D _4628_/A VGND VGND VPWR VPWR _9412_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4885_ _6158_/A _6086_/B input34/X VGND VGND VPWR VPWR _4885_/X sky130_fd_sc_hd__or3b_1
XFILLER_165_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6624_ _6624_/A VGND VGND VPWR VPWR _6624_/Y sky130_fd_sc_hd__clkinv_2
X_9343_ _9344_/CLK _9343_/D _9295_/SET_B VGND VGND VPWR VPWR _9343_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6555_ _9362_/Q VGND VGND VPWR VPWR _6555_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_180_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9274_ _9371_/CLK _9274_/D _9295_/SET_B VGND VGND VPWR VPWR _9274_/Q sky130_fd_sc_hd__dfrtp_1
X_5506_ _9372_/Q _5498_/A _8916_/A1 _5498_/Y VGND VGND VPWR VPWR _9372_/D sky130_fd_sc_hd__a22o_1
X_6486_ _9162_/Q VGND VGND VPWR VPWR _6486_/Y sky130_fd_sc_hd__inv_2
X_8225_ _8305_/B _8260_/B VGND VGND VPWR VPWR _8571_/B sky130_fd_sc_hd__nor2_2
XFILLER_10_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5437_ _9420_/Q _5433_/A _8925_/A1 _5433_/Y VGND VGND VPWR VPWR _9420_/D sky130_fd_sc_hd__a22o_1
Xoutput352 _9043_/Q VGND VGND VPWR VPWR wb_dat_o[31] sky130_fd_sc_hd__buf_2
Xoutput341 _9033_/Q VGND VGND VPWR VPWR wb_dat_o[21] sky130_fd_sc_hd__buf_2
Xoutput330 _9015_/Q VGND VGND VPWR VPWR wb_dat_o[11] sky130_fd_sc_hd__buf_2
XFILLER_105_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5368_ _5368_/A VGND VGND VPWR VPWR _5368_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8156_ _8156_/A _8578_/A VGND VGND VPWR VPWR _8158_/A sky130_fd_sc_hd__or2_1
X_8087_ _8514_/B _8086_/Y VGND VGND VPWR VPWR _8296_/A sky130_fd_sc_hd__or2b_1
X_7107_ _4734_/Y _7048_/D _4769_/Y _7040_/B _7106_/X VGND VGND VPWR VPWR _7108_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_113_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5299_ _5299_/A VGND VGND VPWR VPWR _5300_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7038_ _9246_/Q _9245_/Q _7127_/B _7073_/C VGND VGND VPWR VPWR _7039_/A sky130_fd_sc_hd__or4_1
X_8989_ _9574_/Q _8755_/A VGND VGND VPWR VPWR mgmt_gpio_out[12] sky130_fd_sc_hd__ebufn_8
XFILLER_35_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4670_ _4927_/A _4843_/B VGND VGND VPWR VPWR _5872_/B sky130_fd_sc_hd__or2_4
XFILLER_147_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6340_ _9540_/Q VGND VGND VPWR VPWR _6340_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_127_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6271_ _9525_/Q VGND VGND VPWR VPWR _6271_/Y sky130_fd_sc_hd__inv_6
XFILLER_170_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5222_ _9565_/Q _5218_/Y _8925_/X _5218_/A VGND VGND VPWR VPWR _9565_/D sky130_fd_sc_hd__o22a_1
XFILLER_170_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8010_ _7864_/X _8085_/A _8009_/X VGND VGND VPWR VPWR _8016_/B sky130_fd_sc_hd__o21ai_1
XFILLER_130_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5153_ _9612_/Q _5147_/A _8955_/A1 _5147_/Y VGND VGND VPWR VPWR _9612_/D sky130_fd_sc_hd__a22o_1
XFILLER_130_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5084_ _9657_/Q _5082_/A _5964_/B1 _5082_/Y VGND VGND VPWR VPWR _9657_/D sky130_fd_sc_hd__a22o_1
X_8912_ _7720_/X _9086_/Q _9051_/Q VGND VGND VPWR VPWR _8912_/X sky130_fd_sc_hd__mux2_1
X_8843_ _9704_/Q _9663_/Q _9587_/Q VGND VGND VPWR VPWR _8843_/X sky130_fd_sc_hd__mux2_8
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8774_ _8774_/A VGND VGND VPWR VPWR _8774_/X sky130_fd_sc_hd__clkbuf_1
X_5986_ _9091_/Q _5985_/Y _5981_/X VGND VGND VPWR VPWR _9091_/D sky130_fd_sc_hd__o21ba_1
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4937_ _4636_/Y _8957_/S _4936_/Y _9711_/Q _4636_/A VGND VGND VPWR VPWR _9711_/D
+ sky130_fd_sc_hd__a32o_1
X_7725_ _9088_/Q _7722_/B _7724_/Y _9089_/Q _7722_/Y VGND VGND VPWR VPWR _7725_/X
+ sky130_fd_sc_hd__a32o_1
X_7656_ _6682_/Y _7451_/X _6723_/Y _7453_/X _7655_/X VGND VGND VPWR VPWR _7661_/B
+ sky130_fd_sc_hd__o221a_1
XANTENNA_20 _7662_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_31 _4867_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4868_ _6111_/A _4898_/A VGND VGND VPWR VPWR _4868_/X sky130_fd_sc_hd__or2_4
XANTENNA_53 _6658_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_64 _6863_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6607_ _8769_/A _5458_/B _6606_/Y _5290_/B VGND VGND VPWR VPWR _6607_/X sky130_fd_sc_hd__o22a_1
XANTENNA_42 _6252_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_75 _8783_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_86 _7019_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_97 input80/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7587_ _6188_/Y _7475_/X _6179_/Y _7477_/X VGND VGND VPWR VPWR _7587_/X sky130_fd_sc_hd__o22a_1
X_9326_ _9352_/CLK _9326_/D _9646_/SET_B VGND VGND VPWR VPWR _9326_/Q sky130_fd_sc_hd__dfrtp_1
X_4799_ _4792_/Y _4564_/B _4793_/Y _5240_/B _4798_/X VGND VGND VPWR VPWR _4830_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_4_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6538_ _6538_/A VGND VGND VPWR VPWR _6538_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_137_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9257_ _9601_/CLK _9257_/D _9295_/SET_B VGND VGND VPWR VPWR _9257_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_106_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6469_ _9766_/Q VGND VGND VPWR VPWR _6469_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8208_ _8305_/B _8264_/B VGND VGND VPWR VPWR _8595_/C sky130_fd_sc_hd__nor2_1
XFILLER_79_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9188_ _9758_/CLK _9188_/D _9633_/SET_B VGND VGND VPWR VPWR _9188_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_121_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8139_ _8550_/A _8640_/B VGND VGND VPWR VPWR _8730_/A sky130_fd_sc_hd__nor2_1
XFILLER_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5840_ _9184_/Q _5839_/A _8846_/X _5839_/Y VGND VGND VPWR VPWR _9184_/D sky130_fd_sc_hd__a22o_1
XFILLER_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5771_ _9230_/Q _5770_/A _5963_/B1 _5770_/Y VGND VGND VPWR VPWR _9230_/D sky130_fd_sc_hd__a22o_1
XFILLER_34_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7510_ _6643_/Y _7441_/X _6704_/Y _7443_/X _7509_/X VGND VGND VPWR VPWR _7517_/A
+ sky130_fd_sc_hd__o221a_1
X_4722_ _9226_/Q VGND VGND VPWR VPWR _4722_/Y sky130_fd_sc_hd__inv_2
X_8490_ _8734_/A _8490_/B _8490_/C VGND VGND VPWR VPWR _8597_/D sky130_fd_sc_hd__or3_1
XFILLER_187_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7441_ _7441_/A VGND VGND VPWR VPWR _7441_/X sky130_fd_sc_hd__buf_8
Xinput40 mgmt_gpio_in[13] VGND VGND VPWR VPWR _6317_/A sky130_fd_sc_hd__clkbuf_1
X_4653_ _4994_/A VGND VGND VPWR VPWR _4654_/A sky130_fd_sc_hd__clkbuf_1
Xinput62 mgmt_gpio_in[33] VGND VGND VPWR VPWR input62/X sky130_fd_sc_hd__clkbuf_4
Xinput51 mgmt_gpio_in[23] VGND VGND VPWR VPWR input51/X sky130_fd_sc_hd__clkbuf_2
X_4584_ _9743_/Q _4579_/A _5964_/B1 _4579_/Y VGND VGND VPWR VPWR _9743_/D sky130_fd_sc_hd__a22o_1
Xinput73 pad_flash_io0_di VGND VGND VPWR VPWR _7018_/B sky130_fd_sc_hd__clkbuf_1
X_7372_ _6549_/Y _7126_/X _6609_/Y _7128_/X VGND VGND VPWR VPWR _7372_/X sky130_fd_sc_hd__o22a_1
X_6323_ _8818_/A _4680_/Y input57/X _6322_/Y VGND VGND VPWR VPWR _6323_/Y sky130_fd_sc_hd__a22oi_4
Xinput84 spimemio_flash_csb VGND VGND VPWR VPWR input84/X sky130_fd_sc_hd__buf_4
XFILLER_143_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9111_ _9379_/CLK _9111_/D _9646_/SET_B VGND VGND VPWR VPWR _9111_/Q sky130_fd_sc_hd__dfrtp_1
Xinput95 sram_ro_data[11] VGND VGND VPWR VPWR _6552_/A sky130_fd_sc_hd__clkbuf_1
X_9042_ _9664_/CLK _9042_/D VGND VGND VPWR VPWR _9042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6254_ _6249_/Y _4832_/X _6250_/Y _5110_/B _6253_/X VGND VGND VPWR VPWR _6254_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_170_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5205_ _9576_/Q _5203_/Y _8927_/X _5203_/A VGND VGND VPWR VPWR _9576_/D sky130_fd_sc_hd__o22a_1
XFILLER_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6185_ _6183_/Y _5757_/B _6184_/Y _5797_/B VGND VGND VPWR VPWR _6185_/X sky130_fd_sc_hd__o22a_1
XFILLER_69_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5136_ _5136_/A VGND VGND VPWR VPWR _5136_/Y sky130_fd_sc_hd__inv_2
X_5067_ _5067_/A VGND VGND VPWR VPWR _9665_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8826_ _8825_/X _6505_/A _9682_/Q VGND VGND VPWR VPWR _8826_/X sky130_fd_sc_hd__mux2_1
X_5969_ _5969_/A VGND VGND VPWR VPWR _5970_/A sky130_fd_sc_hd__clkbuf_4
X_8757_ _8757_/A VGND VGND VPWR VPWR _8758_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_25_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7708_ _9082_/Q VGND VGND VPWR VPWR _7708_/Y sky130_fd_sc_hd__clkinv_2
X_8688_ _8688_/A _8688_/B _8688_/C VGND VGND VPWR VPWR _8714_/D sky130_fd_sc_hd__or3_1
X_7639_ _6897_/Y _7465_/X _6848_/Y _7467_/X VGND VGND VPWR VPWR _7639_/X sky130_fd_sc_hd__o22a_1
XFILLER_180_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9309_ _9789_/CLK _9309_/D _9647_/SET_B VGND VGND VPWR VPWR _9309_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_180_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7990_ _8050_/B _7992_/B VGND VGND VPWR VPWR _7991_/A sky130_fd_sc_hd__or2_1
XFILLER_66_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6941_ _6941_/A VGND VGND VPWR VPWR _6941_/Y sky130_fd_sc_hd__inv_2
X_9660_ _9664_/CLK _9660_/D _6146_/A VGND VGND VPWR VPWR _9660_/Q sky130_fd_sc_hd__dfrtp_1
X_6872_ _9386_/Q VGND VGND VPWR VPWR _6872_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_34_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9591_ _9601_/CLK _9591_/D _9295_/SET_B VGND VGND VPWR VPWR _9591_/Q sky130_fd_sc_hd__dfrtp_1
X_8611_ _8064_/C _8610_/Y _8016_/A _8527_/B VGND VGND VPWR VPWR _8613_/B sky130_fd_sc_hd__a211o_1
X_5823_ _9195_/Q _5820_/A _8844_/X _5820_/Y VGND VGND VPWR VPWR _9195_/D sky130_fd_sc_hd__a22o_1
XFILLER_179_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8542_ _8703_/B _8605_/A _8705_/A _8541_/Y VGND VGND VPWR VPWR _8543_/A sky130_fd_sc_hd__or4b_1
XFILLER_147_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5754_ _6997_/A _5643_/Y _5713_/Y _5753_/X VGND VGND VPWR VPWR _5755_/A sky130_fd_sc_hd__a31o_1
X_5685_ _9260_/Q _5681_/A _8925_/A1 _5681_/Y VGND VGND VPWR VPWR _9260_/D sky130_fd_sc_hd__a22o_1
XFILLER_175_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8473_ _8471_/Y _8472_/Y _8061_/A _8708_/C VGND VGND VPWR VPWR _8474_/B sky130_fd_sc_hd__a31o_1
X_4705_ _4705_/A _4705_/B _4705_/C _4705_/D VGND VGND VPWR VPWR _4936_/A sky130_fd_sc_hd__and4_1
XFILLER_147_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4636_ _4636_/A VGND VGND VPWR VPWR _4636_/Y sky130_fd_sc_hd__inv_2
X_7424_ _7462_/A _7470_/B _9255_/Q VGND VGND VPWR VPWR _7425_/A sky130_fd_sc_hd__or3_1
XFILLER_162_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7355_ _6497_/Y _7077_/C _6583_/Y _7077_/D _7354_/X VGND VGND VPWR VPWR _7355_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_190_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6306_ _6301_/Y _5776_/B _6302_/Y _5872_/B _6305_/X VGND VGND VPWR VPWR _6307_/D
+ sky130_fd_sc_hd__o221a_1
X_4567_ _9755_/Q _4566_/A _8846_/X _4566_/Y VGND VGND VPWR VPWR _9755_/D sky130_fd_sc_hd__a22o_1
XFILLER_143_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7286_ _7286_/A _7286_/B _7286_/C _7286_/D VGND VGND VPWR VPWR _7287_/C sky130_fd_sc_hd__and4_1
X_4498_ _9781_/Q _4493_/A _5964_/B1 _4493_/Y VGND VGND VPWR VPWR _9781_/D sky130_fd_sc_hd__a22o_1
X_9025_ _9027_/CLK _9025_/D VGND VGND VPWR VPWR _9025_/Q sky130_fd_sc_hd__dfxtp_1
X_6237_ _6237_/A _6237_/B _6237_/C _6237_/D VGND VGND VPWR VPWR _6237_/Y sky130_fd_sc_hd__nand4_4
X_6168_ _9526_/Q VGND VGND VPWR VPWR _6168_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5119_ _9633_/Q _5112_/A _5966_/B1 _5112_/Y VGND VGND VPWR VPWR _9633_/D sky130_fd_sc_hd__a22o_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6099_ _6099_/A VGND VGND VPWR VPWR _6099_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_27_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_3_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A VGND VGND VPWR VPWR _9279_/CLK sky130_fd_sc_hd__clkbuf_2
X_8809_ _8809_/A VGND VGND VPWR VPWR _8813_/B sky130_fd_sc_hd__inv_2
XFILLER_53_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9789_ _9789_/CLK _9789_/D _9685_/SET_B VGND VGND VPWR VPWR _9789_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5470_ _5470_/A VGND VGND VPWR VPWR _5471_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_157_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7140_ _6865_/Y _7095_/X _6939_/Y _7068_/D _7139_/X VGND VGND VPWR VPWR _7145_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_113_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7071_ _7096_/B _7073_/C VGND VGND VPWR VPWR _7072_/A sky130_fd_sc_hd__or2_1
XFILLER_98_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6022_ _6022_/A _6022_/B _6022_/C _6022_/D VGND VGND VPWR VPWR _6023_/A sky130_fd_sc_hd__or4_1
XFILLER_39_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7973_ _7973_/A VGND VGND VPWR VPWR _8554_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_27_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6924_ _6919_/Y _5949_/B _6920_/Y _5837_/B _6923_/X VGND VGND VPWR VPWR _6925_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_81_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9712_ _9089_/CLK _9712_/D _4654_/X VGND VGND VPWR VPWR _9712_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_81_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9643_ _9776_/CLK _9643_/D _7011_/B VGND VGND VPWR VPWR _9643_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6855_ _9425_/Q VGND VGND VPWR VPWR _6855_/Y sky130_fd_sc_hd__clkinv_2
X_6786_ _6149_/A _6785_/Y _9038_/Q _6149_/Y VGND VGND VPWR VPWR _9038_/D sky130_fd_sc_hd__o22a_1
X_9574_ _9788_/CLK _9574_/D _9646_/SET_B VGND VGND VPWR VPWR _9574_/Q sky130_fd_sc_hd__dfrtp_1
X_5806_ _9205_/Q _5799_/A _8930_/A1 _5799_/Y VGND VGND VPWR VPWR _9205_/D sky130_fd_sc_hd__a22o_1
XFILLER_22_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8525_ _8525_/A _8538_/B _8525_/C VGND VGND VPWR VPWR _8525_/Y sky130_fd_sc_hd__nor3_4
X_5737_ _5737_/A _9245_/Q VGND VGND VPWR VPWR _7125_/A sky130_fd_sc_hd__or2_2
XFILLER_135_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8456_ _7864_/X _8316_/A _8097_/B _8137_/B VGND VGND VPWR VPWR _8734_/C sky130_fd_sc_hd__o22ai_1
X_5668_ _9271_/Q _5662_/A _8841_/X _5662_/Y VGND VGND VPWR VPWR _9271_/D sky130_fd_sc_hd__a22o_1
XFILLER_135_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7407_ _7476_/A _9251_/Q _7470_/B _7474_/D VGND VGND VPWR VPWR _7408_/A sky130_fd_sc_hd__or4_1
XFILLER_151_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5599_ _9309_/Q _5596_/A _8841_/X _5596_/Y VGND VGND VPWR VPWR _9309_/D sky130_fd_sc_hd__a22o_1
X_8387_ _8389_/A _8632_/B VGND VGND VPWR VPWR _8687_/B sky130_fd_sc_hd__nor2_1
X_4619_ _9722_/Q _4615_/A _5966_/B1 _4615_/Y VGND VGND VPWR VPWR _9722_/D sky130_fd_sc_hd__a22o_1
XFILLER_150_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7338_ _6729_/Y _7095_/X _6638_/Y _7068_/D _7337_/X VGND VGND VPWR VPWR _7343_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_89_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7269_ _6129_/Y _7040_/C _6123_/Y _7059_/C VGND VGND VPWR VPWR _7269_/X sky130_fd_sc_hd__o22a_1
X_9008_ _9601_/Q _8793_/A VGND VGND VPWR VPWR mgmt_gpio_out[31] sky130_fd_sc_hd__ebufn_8
XFILLER_18_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4970_ _9706_/Q _4966_/A _9705_/Q _4966_/Y VGND VGND VPWR VPWR _9706_/D sky130_fd_sc_hd__a22o_1
XFILLER_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6640_ _9214_/Q VGND VGND VPWR VPWR _6640_/Y sky130_fd_sc_hd__clkinv_2
X_6571_ _9453_/Q VGND VGND VPWR VPWR _8773_/A sky130_fd_sc_hd__inv_6
XFILLER_145_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8310_ _8571_/B _8310_/B _8497_/A _8309_/X VGND VGND VPWR VPWR _8310_/X sky130_fd_sc_hd__or4b_1
X_5522_ _9362_/Q _5520_/A _5964_/B1 _5520_/Y VGND VGND VPWR VPWR _9362_/D sky130_fd_sc_hd__a22o_1
X_9290_ _9483_/CLK _9290_/D _9528_/SET_B VGND VGND VPWR VPWR _9290_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_117_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5453_ _9410_/Q _5452_/A _5963_/B1 _5452_/Y VGND VGND VPWR VPWR _9410_/D sky130_fd_sc_hd__a22o_1
X_8241_ _8241_/A _8574_/B _8361_/B _8730_/B VGND VGND VPWR VPWR _8245_/A sky130_fd_sc_hd__or4_1
X_5384_ _5384_/A VGND VGND VPWR VPWR _5384_/Y sky130_fd_sc_hd__inv_2
X_8172_ _8172_/A _8373_/A _8171_/X VGND VGND VPWR VPWR _8173_/B sky130_fd_sc_hd__or3b_1
XFILLER_5_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7123_ _7127_/C _7123_/B VGND VGND VPWR VPWR _7124_/A sky130_fd_sc_hd__or2_1
XFILLER_59_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7054_ _7094_/B _7073_/C VGND VGND VPWR VPWR _7055_/A sky130_fd_sc_hd__or2_1
XFILLER_67_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6005_ _9086_/Q _5995_/A _8911_/X _5995_/Y VGND VGND VPWR VPWR _9086_/D sky130_fd_sc_hd__a22o_1
XFILLER_67_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7956_ _8379_/C _8394_/A _8394_/B VGND VGND VPWR VPWR _8099_/B sky130_fd_sc_hd__or3_1
XFILLER_82_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6907_ _6902_/Y _5024_/B _6903_/Y _6135_/A _6906_/X VGND VGND VPWR VPWR _6925_/A
+ sky130_fd_sc_hd__o221a_1
X_7887_ _7836_/B _7879_/Y _7886_/X VGND VGND VPWR VPWR _7887_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_145_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9626_ _8837_/A1 _9626_/D _5130_/X VGND VGND VPWR VPWR _9626_/Q sky130_fd_sc_hd__dfrtp_4
X_6838_ _9633_/Q VGND VGND VPWR VPWR _6838_/Y sky130_fd_sc_hd__inv_2
X_9557_ _9755_/CLK _9557_/D _9633_/SET_B VGND VGND VPWR VPWR _9557_/Q sky130_fd_sc_hd__dfrtp_1
X_8508_ _8282_/C _7831_/Y _8394_/A _7767_/C _8331_/B VGND VGND VPWR VPWR _8662_/B
+ sky130_fd_sc_hd__a41o_1
X_6769_ input5/X VGND VGND VPWR VPWR _6769_/Y sky130_fd_sc_hd__inv_2
X_9488_ _9777_/CLK _9488_/D _9757_/SET_B VGND VGND VPWR VPWR _9488_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_40_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8439_ _8518_/A _8064_/B _8061_/C _8062_/B VGND VGND VPWR VPWR _8617_/A sky130_fd_sc_hd__a31o_1
XFILLER_108_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_110 input86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_132 _7375_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_121 _7015_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_143 _4814_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_154 _8544_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_165 _4901_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_176 _8801_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_187 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput5 mask_rev_in[10] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7810_ _8660_/C _7878_/A VGND VGND VPWR VPWR _7811_/A sky130_fd_sc_hd__or2_1
X_8790_ _8790_/A VGND VGND VPWR VPWR _8790_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_91_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7741_ _9068_/Q _7741_/A2 _9067_/Q _7741_/B2 _7740_/X VGND VGND VPWR VPWR _7741_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4953_ _9708_/Q VGND VGND VPWR VPWR _4953_/Y sky130_fd_sc_hd__inv_2
X_7672_ _6477_/Y _7441_/X _6615_/Y _7443_/X _7671_/X VGND VGND VPWR VPWR _7679_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9411_ _9514_/CLK _9411_/D _9685_/SET_B VGND VGND VPWR VPWR _9411_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6623_ _9781_/Q VGND VGND VPWR VPWR _8781_/A sky130_fd_sc_hd__inv_6
X_4884_ _4911_/A _6111_/B VGND VGND VPWR VPWR _5259_/B sky130_fd_sc_hd__or2_4
XFILLER_165_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9342_ _9508_/CLK _9342_/D _9647_/SET_B VGND VGND VPWR VPWR _9342_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6554_ _6549_/Y _4504_/B _6550_/Y _5259_/B _6553_/X VGND VGND VPWR VPWR _6567_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_173_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9273_ _9535_/CLK _9273_/D _9528_/SET_B VGND VGND VPWR VPWR _9273_/Q sky130_fd_sc_hd__dfrtp_1
X_6485_ _9315_/Q VGND VGND VPWR VPWR _6485_/Y sky130_fd_sc_hd__inv_4
XFILLER_145_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5505_ _9373_/Q _5498_/A _8930_/A1 _5498_/Y VGND VGND VPWR VPWR _9373_/D sky130_fd_sc_hd__a22o_1
X_5436_ _9421_/Q _5433_/A _8844_/X _5433_/Y VGND VGND VPWR VPWR _9421_/D sky130_fd_sc_hd__a22o_1
XFILLER_118_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8224_ _8595_/C _8224_/B _8224_/C _8223_/X VGND VGND VPWR VPWR _8227_/B sky130_fd_sc_hd__or4b_2
Xoutput342 _9034_/Q VGND VGND VPWR VPWR wb_dat_o[22] sky130_fd_sc_hd__buf_2
Xoutput331 _9016_/Q VGND VGND VPWR VPWR wb_dat_o[12] sky130_fd_sc_hd__buf_2
XFILLER_126_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput353 _9023_/Q VGND VGND VPWR VPWR wb_dat_o[3] sky130_fd_sc_hd__buf_2
Xoutput320 _9765_/Q VGND VGND VPWR VPWR sram_ro_addr[3] sky130_fd_sc_hd__buf_2
XFILLER_99_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5367_ _5367_/A VGND VGND VPWR VPWR _5368_/A sky130_fd_sc_hd__clkbuf_2
X_8155_ _8213_/A _8552_/A VGND VGND VPWR VPWR _8578_/A sky130_fd_sc_hd__nor2_1
X_8086_ _8086_/A _8086_/B VGND VGND VPWR VPWR _8086_/Y sky130_fd_sc_hd__nand2_1
XFILLER_141_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7106_ _4708_/Y _7068_/A _4793_/Y _7105_/X VGND VGND VPWR VPWR _7106_/X sky130_fd_sc_hd__o22a_1
X_5298_ _5671_/A _5298_/B VGND VGND VPWR VPWR _5299_/A sky130_fd_sc_hd__or2_1
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7037_ _7037_/A _9247_/Q VGND VGND VPWR VPWR _7127_/B sky130_fd_sc_hd__or2_2
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8988_ _9573_/Q _8753_/A VGND VGND VPWR VPWR mgmt_gpio_out[11] sky130_fd_sc_hd__ebufn_8
XFILLER_15_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7939_ _8202_/A _8510_/A _7938_/Y VGND VGND VPWR VPWR _7939_/X sky130_fd_sc_hd__o21ba_1
XFILLER_70_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9609_ _9617_/CLK _9609_/D _9295_/SET_B VGND VGND VPWR VPWR _9609_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6270_ _6270_/A VGND VGND VPWR VPWR _6270_/Y sky130_fd_sc_hd__clkinv_2
X_5221_ _9566_/Q _5218_/Y _8921_/X _5218_/A VGND VGND VPWR VPWR _9566_/D sky130_fd_sc_hd__o22a_1
XFILLER_88_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5152_ _9613_/Q _5147_/A _8929_/A1 _5147_/Y VGND VGND VPWR VPWR _9613_/D sky130_fd_sc_hd__a22o_1
XFILLER_110_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5083_ _9658_/Q _5082_/A _5963_/B1 _5082_/Y VGND VGND VPWR VPWR _9658_/D sky130_fd_sc_hd__a22o_1
XFILLER_110_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8911_ _7717_/X _9085_/Q _9051_/Q VGND VGND VPWR VPWR _8911_/X sky130_fd_sc_hd__mux2_1
X_8842_ _9703_/Q _9662_/Q _9587_/Q VGND VGND VPWR VPWR _8842_/X sky130_fd_sc_hd__mux2_8
XFILLER_25_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8773_ _8773_/A VGND VGND VPWR VPWR _8774_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_64_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5985_ _6022_/C _5985_/B VGND VGND VPWR VPWR _5985_/Y sky130_fd_sc_hd__nor2_1
X_7724_ _9089_/Q VGND VGND VPWR VPWR _7724_/Y sky130_fd_sc_hd__inv_2
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4936_ _4936_/A _4936_/B _4936_/C VGND VGND VPWR VPWR _4936_/Y sky130_fd_sc_hd__nand3_4
XFILLER_52_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4867_ _4867_/A VGND VGND VPWR VPWR _4867_/Y sky130_fd_sc_hd__inv_4
X_7655_ _6662_/Y _7455_/X _6745_/Y _7457_/X VGND VGND VPWR VPWR _7655_/X sky130_fd_sc_hd__o22a_1
XANTENNA_10 _7287_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_32 _4910_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_21 _5259_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7586_ _6194_/Y _7461_/X _6168_/Y _7463_/X _7585_/X VGND VGND VPWR VPWR _7589_/C
+ sky130_fd_sc_hd__o221a_1
XANTENNA_43 _6254_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_65 _7133_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_54 _6676_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6606_ _9518_/Q VGND VGND VPWR VPWR _6606_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_87 _7019_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_98 input81/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_76 _4450_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_9325_ _9613_/CLK _9325_/D _9646_/SET_B VGND VGND VPWR VPWR _9325_/Q sky130_fd_sc_hd__dfrtp_1
X_6537_ _9109_/Q VGND VGND VPWR VPWR _7703_/A sky130_fd_sc_hd__clkinv_4
X_4798_ _4795_/Y _5121_/B _4797_/Y _4613_/B VGND VGND VPWR VPWR _4798_/X sky130_fd_sc_hd__o22a_1
XFILLER_192_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9256_ _9601_/CLK _9256_/D _9528_/SET_B VGND VGND VPWR VPWR _9256_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_97_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6468_ _9155_/Q VGND VGND VPWR VPWR _6468_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8207_ _8207_/A VGND VGND VPWR VPWR _8264_/B sky130_fd_sc_hd__buf_6
XFILLER_106_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5419_ _9432_/Q _5414_/A _5967_/B1 _5414_/Y VGND VGND VPWR VPWR _9432_/D sky130_fd_sc_hd__a22o_1
X_6399_ _9467_/Q VGND VGND VPWR VPWR _6399_/Y sky130_fd_sc_hd__inv_2
X_9187_ _9757_/CLK _9187_/D _9633_/SET_B VGND VGND VPWR VPWR _9187_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_153_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8138_ _8164_/A _8550_/A VGND VGND VPWR VPWR _8361_/A sky130_fd_sc_hd__nor2_1
XFILLER_87_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8069_ _8069_/A _8203_/A VGND VGND VPWR VPWR _8069_/Y sky130_fd_sc_hd__nand2_1
XFILLER_153_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5770_ _5770_/A VGND VGND VPWR VPWR _5770_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4721_ _4917_/A _4780_/B VGND VGND VPWR VPWR _5679_/B sky130_fd_sc_hd__or2_4
XFILLER_61_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7440_ _7462_/A _7476_/C _9255_/Q VGND VGND VPWR VPWR _7441_/A sky130_fd_sc_hd__or3_1
X_4652_ _9713_/Q _4636_/A _8951_/X _4636_/Y VGND VGND VPWR VPWR _9713_/D sky130_fd_sc_hd__a22o_1
XFILLER_147_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput30 mask_rev_in[4] VGND VGND VPWR VPWR _6470_/A sky130_fd_sc_hd__clkbuf_1
Xinput63 mgmt_gpio_in[34] VGND VGND VPWR VPWR _8803_/A sky130_fd_sc_hd__buf_6
Xinput52 mgmt_gpio_in[24] VGND VGND VPWR VPWR _4781_/A sky130_fd_sc_hd__clkbuf_1
Xinput41 mgmt_gpio_in[14] VGND VGND VPWR VPWR input41/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7371_ _6543_/Y _5728_/X _6529_/Y _7040_/A _7370_/X VGND VGND VPWR VPWR _7374_/C
+ sky130_fd_sc_hd__o221a_1
X_9110_ _9695_/CLK _9110_/D _9779_/SET_B VGND VGND VPWR VPWR _9110_/Q sky130_fd_sc_hd__dfrtp_1
X_4583_ _9744_/Q _4579_/A _5963_/B1 _4579_/Y VGND VGND VPWR VPWR _9744_/D sky130_fd_sc_hd__a22o_1
Xinput85 spimemio_flash_io0_do VGND VGND VPWR VPWR input85/X sky130_fd_sc_hd__buf_4
X_6322_ _6322_/A VGND VGND VPWR VPWR _6322_/Y sky130_fd_sc_hd__inv_6
XFILLER_155_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput74 pad_flash_io1_di VGND VGND VPWR VPWR _7020_/B sky130_fd_sc_hd__buf_2
Xinput96 sram_ro_data[12] VGND VGND VPWR VPWR _6336_/A sky130_fd_sc_hd__clkbuf_1
X_9041_ _9664_/CLK _9041_/D VGND VGND VPWR VPWR _9041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6253_ _8822_/X _6251_/Y _6252_/Y _4841_/X VGND VGND VPWR VPWR _6253_/X sky130_fd_sc_hd__o2bb2a_1
X_5204_ _9577_/Q _5203_/Y _8898_/X _5203_/A VGND VGND VPWR VPWR _9577_/D sky130_fd_sc_hd__o22a_1
XFILLER_103_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6184_ _9210_/Q VGND VGND VPWR VPWR _6184_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_111_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5135_ _5135_/A VGND VGND VPWR VPWR _5136_/A sky130_fd_sc_hd__clkbuf_4
X_5066_ _8967_/X _9665_/Q _5078_/S VGND VGND VPWR VPWR _5067_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8825_ _9579_/Q _9718_/Q _8977_/S VGND VGND VPWR VPWR _8825_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5968_ _6052_/A _5968_/B VGND VGND VPWR VPWR _5969_/A sky130_fd_sc_hd__or2_1
X_8756_ _8756_/A VGND VGND VPWR VPWR _8756_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_166_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7707_ _9049_/Q _9052_/Q VGND VGND VPWR VPWR _7707_/Y sky130_fd_sc_hd__nor2_1
X_4919_ _4919_/A _4931_/B VGND VGND VPWR VPWR _5480_/B sky130_fd_sc_hd__or2_4
XFILLER_178_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5899_ _5899_/A VGND VGND VPWR VPWR _5899_/Y sky130_fd_sc_hd__inv_2
X_8687_ _8720_/A _8687_/B _8687_/C VGND VGND VPWR VPWR _8713_/C sky130_fd_sc_hd__or3_1
XFILLER_32_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7638_ _6883_/Y _7451_/X _6873_/Y _7453_/X _7637_/X VGND VGND VPWR VPWR _7643_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_20_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7569_ _6291_/Y _7475_/X _6316_/Y _7477_/X VGND VGND VPWR VPWR _7569_/X sky130_fd_sc_hd__o22a_1
XFILLER_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9308_ _9789_/CLK _9308_/D _9647_/SET_B VGND VGND VPWR VPWR _9308_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9239_ _9279_/CLK _9239_/D _9757_/SET_B VGND VGND VPWR VPWR _9239_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_164_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6940_ _9655_/Q VGND VGND VPWR VPWR _6940_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_66_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6871_ _9399_/Q VGND VGND VPWR VPWR _6871_/Y sky130_fd_sc_hd__clkinv_4
X_9590_ _9601_/CLK _9590_/D _9295_/SET_B VGND VGND VPWR VPWR _9590_/Q sky130_fd_sc_hd__dfrtp_1
X_8610_ _8189_/A _7885_/X _7881_/A VGND VGND VPWR VPWR _8610_/Y sky130_fd_sc_hd__o21ai_1
X_5822_ _9196_/Q _5820_/A _8845_/X _5820_/Y VGND VGND VPWR VPWR _9196_/D sky130_fd_sc_hd__a22o_1
XFILLER_148_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8541_ _8541_/A _8617_/B _8705_/D _8619_/D VGND VGND VPWR VPWR _8541_/Y sky130_fd_sc_hd__nor4_1
X_5753_ _9056_/Q _5753_/B _5787_/A VGND VGND VPWR VPWR _5753_/X sky130_fd_sc_hd__and3_1
X_4704_ _4694_/Y _5864_/B _4696_/Y _6165_/A _4703_/X VGND VGND VPWR VPWR _4705_/D
+ sky130_fd_sc_hd__o221a_1
X_5684_ _9261_/Q _5681_/A _8844_/X _5681_/Y VGND VGND VPWR VPWR _9261_/D sky130_fd_sc_hd__a22o_1
X_8472_ _8472_/A VGND VGND VPWR VPWR _8472_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_30_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7423_ _4708_/Y _7415_/X _4701_/Y _7417_/X _7422_/X VGND VGND VPWR VPWR _7481_/B
+ sky130_fd_sc_hd__o221a_1
X_4635_ _4635_/A VGND VGND VPWR VPWR _4636_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_147_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7354_ _6556_/Y _7086_/X _6612_/Y _7088_/X VGND VGND VPWR VPWR _7354_/X sky130_fd_sc_hd__o22a_1
X_4566_ _4566_/A VGND VGND VPWR VPWR _4566_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_150_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6305_ _6303_/Y _5968_/B _6304_/Y _5905_/B VGND VGND VPWR VPWR _6305_/X sky130_fd_sc_hd__o22a_1
X_9024_ _9027_/CLK _9024_/D VGND VGND VPWR VPWR _9024_/Q sky130_fd_sc_hd__dfxtp_1
X_7285_ _6090_/Y _7124_/X _6061_/Y _7068_/B _7284_/X VGND VGND VPWR VPWR _7286_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_103_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4497_ _9782_/Q _4493_/A _5963_/B1 _4493_/Y VGND VGND VPWR VPWR _9782_/D sky130_fd_sc_hd__a22o_1
XFILLER_103_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6236_ _6236_/A _6236_/B _6236_/C _6236_/D VGND VGND VPWR VPWR _6237_/D sky130_fd_sc_hd__and4_2
X_6167_ _6163_/Y _5583_/B _6164_/Y _5458_/B _6166_/Y VGND VGND VPWR VPWR _6174_/C
+ sky130_fd_sc_hd__o221a_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5118_ _9634_/Q _5112_/A _5965_/B1 _5112_/Y VGND VGND VPWR VPWR _9634_/D sky130_fd_sc_hd__a22o_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6098_ _9353_/Q VGND VGND VPWR VPWR _6098_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5049_ _9673_/Q _5047_/A _8845_/X _5047_/Y VGND VGND VPWR VPWR _9673_/D sky130_fd_sc_hd__a22o_1
XFILLER_57_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8808_ _8808_/A _8808_/B VGND VGND VPWR VPWR _8808_/Y sky130_fd_sc_hd__nor2_2
X_9788_ _9788_/CLK _9788_/D _9646_/SET_B VGND VGND VPWR VPWR _9788_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_80_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8739_ _8739_/A VGND VGND VPWR VPWR _8739_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7070_ _7070_/A VGND VGND VPWR VPWR _7077_/A sky130_fd_sc_hd__buf_8
XFILLER_113_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6021_ _6021_/A VGND VGND VPWR VPWR _6021_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_58_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_1_csclk clkbuf_1_1_1_csclk/A VGND VGND VPWR VPWR clkbuf_2_3_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_39_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7972_ _8096_/B _8116_/A VGND VGND VPWR VPWR _7973_/A sky130_fd_sc_hd__or2_1
XFILLER_94_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6923_ _6921_/Y _5013_/B _6922_/Y _5916_/B VGND VGND VPWR VPWR _6923_/X sky130_fd_sc_hd__o22a_1
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9711_ _9709_/CLK _9711_/D _4657_/X VGND VGND VPWR VPWR _9711_/Q sky130_fd_sc_hd__dfrtn_1
X_9642_ _9776_/CLK _9642_/D _4628_/A VGND VGND VPWR VPWR _9642_/Q sky130_fd_sc_hd__dfrtp_1
X_6854_ _9503_/Q VGND VGND VPWR VPWR _6854_/Y sky130_fd_sc_hd__inv_2
XFILLER_167_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5805_ _9206_/Q _5799_/A _8955_/A1 _5799_/Y VGND VGND VPWR VPWR _9206_/D sky130_fd_sc_hd__a22o_1
X_9573_ _9613_/CLK _9573_/D _9646_/SET_B VGND VGND VPWR VPWR _9573_/Q sky130_fd_sc_hd__dfrtp_1
X_6785_ _6785_/A _6785_/B _6785_/C VGND VGND VPWR VPWR _6785_/Y sky130_fd_sc_hd__nand3_4
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8524_ _8523_/Y _8517_/Y _8518_/X _8444_/A VGND VGND VPWR VPWR _8527_/C sky130_fd_sc_hd__a31o_1
XFILLER_22_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5736_ _5724_/B _7104_/A _7056_/B _5692_/A _5735_/X VGND VGND VPWR VPWR _9247_/D
+ sky130_fd_sc_hd__o311a_1
X_5667_ _9272_/Q _5662_/A _8929_/A1 _5662_/Y VGND VGND VPWR VPWR _9272_/D sky130_fd_sc_hd__a22o_1
XFILLER_148_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8455_ _8455_/A _8455_/B VGND VGND VPWR VPWR _8459_/A sky130_fd_sc_hd__or2_1
XFILLER_175_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4618_ _9723_/Q _4615_/A _5965_/B1 _4615_/Y VGND VGND VPWR VPWR _9723_/D sky130_fd_sc_hd__a22o_1
X_7406_ _9254_/Q _7406_/B VGND VGND VPWR VPWR _7470_/B sky130_fd_sc_hd__or2_4
XFILLER_190_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8386_ _8386_/A _8386_/B VGND VGND VPWR VPWR _8632_/B sky130_fd_sc_hd__or2_1
XFILLER_135_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5598_ _9310_/Q _5596_/A _8842_/X _5596_/Y VGND VGND VPWR VPWR _9310_/D sky130_fd_sc_hd__a22o_1
XFILLER_190_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4549_ _8811_/A _8975_/S VGND VGND VPWR VPWR _4551_/B sky130_fd_sc_hd__nand2_8
XFILLER_150_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7337_ _6780_/Y _7097_/X _6711_/Y _7099_/X VGND VGND VPWR VPWR _7337_/X sky130_fd_sc_hd__o22a_1
XFILLER_145_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7268_ _6073_/Y _7082_/X _6114_/Y _7084_/X _7267_/X VGND VGND VPWR VPWR _7287_/A
+ sky130_fd_sc_hd__o221a_1
X_9007_ _9600_/Q _8791_/A VGND VGND VPWR VPWR mgmt_gpio_out[30] sky130_fd_sc_hd__ebufn_8
XFILLER_131_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6219_ _6219_/A VGND VGND VPWR VPWR _6219_/Y sky130_fd_sc_hd__clkinv_2
X_7199_ _7199_/A _7199_/B _7199_/C VGND VGND VPWR VPWR _7199_/Y sky130_fd_sc_hd__nand3_4
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6570_ _6570_/A VGND VGND VPWR VPWR _6570_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5521_ _9363_/Q _5520_/A _5963_/B1 _5520_/Y VGND VGND VPWR VPWR _9363_/D sky130_fd_sc_hd__a22o_1
XFILLER_117_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8240_ _8316_/A _8264_/B VGND VGND VPWR VPWR _8730_/B sky130_fd_sc_hd__nor2_1
XFILLER_172_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5452_ _5452_/A VGND VGND VPWR VPWR _5452_/Y sky130_fd_sc_hd__clkinv_2
X_5383_ _5383_/A VGND VGND VPWR VPWR _5384_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_145_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8171_ _8396_/A _8397_/B VGND VGND VPWR VPWR _8171_/X sky130_fd_sc_hd__or2_1
XFILLER_117_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7122_ _4816_/Y _5728_/X _4842_/Y _7040_/A _7121_/X VGND VGND VPWR VPWR _7131_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_140_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7053_ _7053_/A VGND VGND VPWR VPWR _7059_/B sky130_fd_sc_hd__buf_8
XFILLER_115_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6004_ _6004_/A VGND VGND VPWR VPWR _6004_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_101_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7955_ _8437_/B _8164_/A VGND VGND VPWR VPWR _8585_/B sky130_fd_sc_hd__nor2_2
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7886_ _8566_/A _7886_/B _7879_/B _7885_/X VGND VGND VPWR VPWR _7886_/X sky130_fd_sc_hd__or4bb_1
X_6906_ _6904_/Y _5526_/B _6905_/Y _6081_/B VGND VGND VPWR VPWR _6906_/X sky130_fd_sc_hd__o22a_1
X_6837_ _9628_/Q VGND VGND VPWR VPWR _6837_/Y sky130_fd_sc_hd__inv_2
X_9625_ _9674_/CLK _9625_/D _9633_/SET_B VGND VGND VPWR VPWR _9625_/Q sky130_fd_sc_hd__dfrtp_1
X_9556_ _9777_/CLK _9556_/D _9633_/SET_B VGND VGND VPWR VPWR _9556_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_24_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8507_ _7879_/A _7881_/A _7848_/A _8300_/B _7931_/A VGND VGND VPWR VPWR _8600_/B
+ sky130_fd_sc_hd__o221ai_2
X_6768_ _9750_/Q VGND VGND VPWR VPWR _6768_/Y sky130_fd_sc_hd__inv_2
X_6699_ _9742_/Q VGND VGND VPWR VPWR _6699_/Y sky130_fd_sc_hd__inv_2
X_9487_ _9777_/CLK _9487_/D _7011_/B VGND VGND VPWR VPWR _9487_/Q sky130_fd_sc_hd__dfrtp_1
X_5719_ _5737_/A _5738_/B VGND VGND VPWR VPWR _7104_/A sky130_fd_sc_hd__or2_2
XFILLER_163_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8438_ _8515_/A _8521_/B VGND VGND VPWR VPWR _8703_/D sky130_fd_sc_hd__nor2_1
XFILLER_156_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8369_ _8630_/B _8369_/B VGND VGND VPWR VPWR _8645_/C sky130_fd_sc_hd__or2_1
XFILLER_151_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_100 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_111 input86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_122 _7015_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_133 _7554_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_155 _8544_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_144 _4850_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_166 _8801_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_177 _8801_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_188 _6135_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput6 mask_rev_in[11] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7740_ _9066_/Q _7740_/B VGND VGND VPWR VPWR _7740_/X sky130_fd_sc_hd__and2_1
XFILLER_101_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4952_ _9709_/Q VGND VGND VPWR VPWR _4952_/Y sky130_fd_sc_hd__inv_2
XFILLER_177_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7671_ _6612_/Y _7445_/X _6587_/Y _7447_/X VGND VGND VPWR VPWR _7671_/X sky130_fd_sc_hd__o22a_1
X_4883_ _9536_/Q VGND VGND VPWR VPWR _4883_/Y sky130_fd_sc_hd__inv_2
X_6622_ _9523_/Q VGND VGND VPWR VPWR _8787_/A sky130_fd_sc_hd__inv_8
X_9410_ _9514_/CLK _9410_/D _4628_/A VGND VGND VPWR VPWR _9410_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9341_ _9344_/CLK _9341_/D _9295_/SET_B VGND VGND VPWR VPWR _9341_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6553_ _6551_/Y _5100_/B _6552_/Y _4893_/X VGND VGND VPWR VPWR _6553_/X sky130_fd_sc_hd__o22a_1
X_9272_ _9344_/CLK _9272_/D _9295_/SET_B VGND VGND VPWR VPWR _9272_/Q sky130_fd_sc_hd__dfrtp_1
X_6484_ _9310_/Q VGND VGND VPWR VPWR _6484_/Y sky130_fd_sc_hd__inv_2
X_5504_ _9374_/Q _5498_/A _8955_/A1 _5498_/Y VGND VGND VPWR VPWR _9374_/D sky130_fd_sc_hd__a22o_1
X_5435_ _9422_/Q _5433_/A _8845_/X _5433_/Y VGND VGND VPWR VPWR _9422_/D sky130_fd_sc_hd__a22o_1
XFILLER_173_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8223_ _8223_/A _8223_/B VGND VGND VPWR VPWR _8223_/X sky130_fd_sc_hd__and2_1
XFILLER_118_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput310 _8820_/X VGND VGND VPWR VPWR serial_load sky130_fd_sc_hd__buf_2
Xoutput343 _9035_/Q VGND VGND VPWR VPWR wb_dat_o[23] sky130_fd_sc_hd__buf_2
Xoutput332 _9017_/Q VGND VGND VPWR VPWR wb_dat_o[13] sky130_fd_sc_hd__buf_2
Xoutput321 _9766_/Q VGND VGND VPWR VPWR sram_ro_addr[4] sky130_fd_sc_hd__buf_2
Xoutput354 _9024_/Q VGND VGND VPWR VPWR wb_dat_o[4] sky130_fd_sc_hd__buf_2
X_5366_ _5671_/A _5366_/B VGND VGND VPWR VPWR _5367_/A sky130_fd_sc_hd__or2_1
X_8154_ _8154_/A _8367_/A VGND VGND VPWR VPWR _8156_/A sky130_fd_sc_hd__or2_1
X_8085_ _8085_/A _8538_/D VGND VGND VPWR VPWR _8086_/B sky130_fd_sc_hd__or2_1
XFILLER_99_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5297_ _9515_/Q _5292_/A _5967_/B1 _5292_/Y VGND VGND VPWR VPWR _9515_/D sky130_fd_sc_hd__a22o_1
X_7105_ _7105_/A VGND VGND VPWR VPWR _7105_/X sky130_fd_sc_hd__buf_8
XFILLER_142_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7036_ _7036_/A VGND VGND VPWR VPWR _7040_/C sky130_fd_sc_hd__buf_6
XFILLER_142_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8987_ _8987_/A _8751_/A VGND VGND VPWR VPWR mgmt_gpio_out[10] sky130_fd_sc_hd__ebufn_8
XFILLER_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7938_ _8094_/A _7938_/B VGND VGND VPWR VPWR _7938_/Y sky130_fd_sc_hd__nand2_1
XFILLER_27_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9608_ _9617_/CLK _9608_/D _9295_/SET_B VGND VGND VPWR VPWR _9608_/Q sky130_fd_sc_hd__dfrtp_1
X_7869_ _8226_/C _8316_/A VGND VGND VPWR VPWR _7870_/A sky130_fd_sc_hd__or2_1
XFILLER_11_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9539_ _9768_/CLK _9539_/D _4628_/A VGND VGND VPWR VPWR _9539_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_136_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_41_csclk clkbuf_2_1_0_csclk/X VGND VGND VPWR VPWR _9779_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_159_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5220_ _9567_/Q _5218_/Y _8918_/X _5218_/A VGND VGND VPWR VPWR _9567_/D sky130_fd_sc_hd__o22a_1
XFILLER_155_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5151_ _9614_/Q _5147_/A _8925_/A1 _5147_/Y VGND VGND VPWR VPWR _9614_/D sky130_fd_sc_hd__a22o_1
XFILLER_142_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5082_ _5082_/A VGND VGND VPWR VPWR _5082_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8910_ _7715_/Y _9084_/Q _9051_/Q VGND VGND VPWR VPWR _8910_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8841_ _9702_/Q _9661_/Q _9587_/Q VGND VGND VPWR VPWR _8841_/X sky130_fd_sc_hd__mux2_8
XFILLER_112_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8772_ _8772_/A VGND VGND VPWR VPWR _8772_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_92_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5984_ _5984_/A VGND VGND VPWR VPWR _5984_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7723_ _9088_/Q _7722_/B _7722_/Y VGND VGND VPWR VPWR _7723_/X sky130_fd_sc_hd__o21a_1
X_4935_ _4935_/A _4935_/B _4935_/C _4935_/D VGND VGND VPWR VPWR _4936_/C sky130_fd_sc_hd__and4_2
XFILLER_177_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_22 _4481_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7654_ _6638_/Y _7441_/X _6705_/Y _7443_/X _7653_/X VGND VGND VPWR VPWR _7661_/A
+ sky130_fd_sc_hd__o221a_1
XANTENNA_11 _7309_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4866_ _4911_/A _4925_/A VGND VGND VPWR VPWR _5336_/B sky130_fd_sc_hd__or2_4
XFILLER_165_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7585_ _6184_/Y _7465_/X _6160_/Y _7467_/X VGND VGND VPWR VPWR _7585_/X sky130_fd_sc_hd__o22a_1
XANTENNA_33 _5278_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_66 _7308_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_55 _6716_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4797_ _9721_/Q VGND VGND VPWR VPWR _4797_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6605_ _9401_/Q VGND VGND VPWR VPWR _8769_/A sky130_fd_sc_hd__inv_8
XANTENNA_44 _6256_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9324_ _9352_/CLK _9324_/D _9646_/SET_B VGND VGND VPWR VPWR _9324_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_88 input37/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6536_ _6531_/Y _6322_/A _7699_/A _5872_/B _6535_/X VGND VGND VPWR VPWR _6536_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_20_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_99 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_77 _6326_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6467_ _9189_/Q VGND VGND VPWR VPWR _6467_/Y sky130_fd_sc_hd__inv_2
X_9255_ _9279_/CLK _9255_/D _9779_/SET_B VGND VGND VPWR VPWR _9255_/Q sky130_fd_sc_hd__dfstp_4
X_8206_ _8272_/A _8226_/C VGND VGND VPWR VPWR _8207_/A sky130_fd_sc_hd__or2_1
X_5418_ _9433_/Q _5414_/A _5966_/B1 _5414_/Y VGND VGND VPWR VPWR _9433_/D sky130_fd_sc_hd__a22o_1
X_6398_ _9350_/Q VGND VGND VPWR VPWR _6398_/Y sky130_fd_sc_hd__inv_2
X_9186_ _9758_/CLK _9186_/D _9633_/SET_B VGND VGND VPWR VPWR _9186_/Q sky130_fd_sc_hd__dfrtp_1
X_5349_ _9481_/Q _5346_/A _8844_/X _5346_/Y VGND VGND VPWR VPWR _9481_/D sky130_fd_sc_hd__a22o_1
XFILLER_133_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8137_ _8213_/A _8137_/B VGND VGND VPWR VPWR _8574_/A sky130_fd_sc_hd__nor2_1
X_8068_ _8515_/A _8164_/A VGND VGND VPWR VPWR _8203_/A sky130_fd_sc_hd__or2_1
XFILLER_153_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7019_ _7019_/A VGND VGND VPWR VPWR _7019_/X sky130_fd_sc_hd__buf_6
XFILLER_28_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4720_ _9256_/Q VGND VGND VPWR VPWR _4720_/Y sky130_fd_sc_hd__clkinv_4
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4651_ _4651_/A VGND VGND VPWR VPWR _4651_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_147_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput31 mask_rev_in[5] VGND VGND VPWR VPWR _6257_/A sky130_fd_sc_hd__clkbuf_1
Xinput20 mask_rev_in[24] VGND VGND VPWR VPWR _4821_/A sky130_fd_sc_hd__clkbuf_1
Xinput64 mgmt_gpio_in[35] VGND VGND VPWR VPWR _6538_/A sky130_fd_sc_hd__clkbuf_1
Xinput53 mgmt_gpio_in[25] VGND VGND VPWR VPWR input53/X sky130_fd_sc_hd__clkbuf_4
XFILLER_162_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput42 mgmt_gpio_in[15] VGND VGND VPWR VPWR input42/X sky130_fd_sc_hd__clkbuf_1
X_7370_ _7370_/A _7392_/B VGND VGND VPWR VPWR _7370_/X sky130_fd_sc_hd__or2_1
X_4582_ _9745_/Q _4579_/A _8844_/X _4579_/Y VGND VGND VPWR VPWR _9745_/D sky130_fd_sc_hd__a22o_1
Xinput86 spimemio_flash_io0_oeb VGND VGND VPWR VPWR input86/X sky130_fd_sc_hd__buf_6
X_6321_ _9369_/Q VGND VGND VPWR VPWR _6321_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_115_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput75 porb VGND VGND VPWR VPWR _7011_/B sky130_fd_sc_hd__buf_12
Xinput97 sram_ro_data[13] VGND VGND VPWR VPWR _6292_/A sky130_fd_sc_hd__clkbuf_1
X_9040_ _9664_/CLK _9040_/D VGND VGND VPWR VPWR _9040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6252_ _6252_/A VGND VGND VPWR VPWR _6252_/Y sky130_fd_sc_hd__clkinv_2
X_6183_ _9237_/Q VGND VGND VPWR VPWR _6183_/Y sky130_fd_sc_hd__clkinv_2
X_5203_ _5203_/A VGND VGND VPWR VPWR _5203_/Y sky130_fd_sc_hd__inv_2
X_5134_ _6165_/A _5156_/B VGND VGND VPWR VPWR _5135_/A sky130_fd_sc_hd__or2_1
XFILLER_111_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5065_ _5065_/A VGND VGND VPWR VPWR _9666_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8824_ _9578_/Q input3/X input1/X VGND VGND VPWR VPWR _8824_/X sky130_fd_sc_hd__mux2_2
XFILLER_16_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8755_ _8755_/A VGND VGND VPWR VPWR _8756_/A sky130_fd_sc_hd__clkbuf_1
X_5967_ _9101_/Q _5962_/A _5967_/B1 _5962_/Y VGND VGND VPWR VPWR _9101_/D sky130_fd_sc_hd__a22o_1
XFILLER_40_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8686_ _8686_/A _8686_/B _8686_/C _8686_/D VGND VGND VPWR VPWR _8709_/D sky130_fd_sc_hd__or4_2
X_4918_ _9385_/Q VGND VGND VPWR VPWR _4918_/Y sky130_fd_sc_hd__clkinv_2
X_7706_ _7706_/A VGND VGND VPWR VPWR _7706_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_166_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5898_ _5898_/A VGND VGND VPWR VPWR _5899_/A sky130_fd_sc_hd__clkbuf_2
X_7637_ _6898_/Y _7455_/X _6833_/Y _7457_/X VGND VGND VPWR VPWR _7637_/X sky130_fd_sc_hd__o22a_1
XFILLER_32_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4849_ _6111_/B _4931_/B VGND VGND VPWR VPWR _5442_/B sky130_fd_sc_hd__or2_4
X_7568_ _6284_/Y _7461_/X _6271_/Y _7463_/X _7567_/X VGND VGND VPWR VPWR _7571_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_180_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9307_ _9789_/CLK _9307_/D _9685_/SET_B VGND VGND VPWR VPWR _9307_/Q sky130_fd_sc_hd__dfrtp_1
X_7499_ _7499_/A _7499_/B _7499_/C _7499_/D VGND VGND VPWR VPWR _7500_/D sky130_fd_sc_hd__and4_1
X_6519_ _8749_/A _5818_/B _8759_/A _5660_/B _6518_/X VGND VGND VPWR VPWR _6526_/C
+ sky130_fd_sc_hd__o221a_1
X_9238_ _9371_/CLK _9238_/D _9295_/SET_B VGND VGND VPWR VPWR _9238_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_134_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9169_ _9203_/CLK _9169_/D _9633_/SET_B VGND VGND VPWR VPWR _9169_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6870_ _6865_/Y _5344_/B _6866_/Y _5366_/B _6869_/X VGND VGND VPWR VPWR _6877_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_179_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5821_ _9197_/Q _5820_/A _8846_/X _5820_/Y VGND VGND VPWR VPWR _9197_/D sky130_fd_sc_hd__a22o_1
X_8540_ _8540_/A _8704_/B VGND VGND VPWR VPWR _8619_/D sky130_fd_sc_hd__or2_1
XFILLER_15_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5752_ _9280_/Q _9279_/Q _9278_/Q VGND VGND VPWR VPWR _5787_/A sky130_fd_sc_hd__or3_1
XFILLER_148_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4703_ _4699_/Y _5897_/B _4701_/Y _5013_/B VGND VGND VPWR VPWR _4703_/X sky130_fd_sc_hd__o22a_1
X_5683_ _9262_/Q _5681_/A _8845_/X _5681_/Y VGND VGND VPWR VPWR _9262_/D sky130_fd_sc_hd__a22o_1
X_8471_ _8538_/C VGND VGND VPWR VPWR _8471_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_30_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7422_ _4773_/Y _7419_/X _4857_/Y _7421_/X VGND VGND VPWR VPWR _7422_/X sky130_fd_sc_hd__o22a_1
X_4634_ _5214_/A _4964_/B VGND VGND VPWR VPWR _4635_/A sky130_fd_sc_hd__or2_1
XFILLER_175_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7353_ _7353_/A _7353_/B _7353_/C VGND VGND VPWR VPWR _7353_/Y sky130_fd_sc_hd__nand3_4
X_4565_ _4565_/A VGND VGND VPWR VPWR _4566_/A sky130_fd_sc_hd__buf_2
X_6304_ _9130_/Q VGND VGND VPWR VPWR _6304_/Y sky130_fd_sc_hd__inv_2
X_9023_ _9027_/CLK _9023_/D VGND VGND VPWR VPWR _9023_/Q sky130_fd_sc_hd__dfxtp_1
X_7284_ _6104_/Y _7126_/X _6116_/Y _7128_/X VGND VGND VPWR VPWR _7284_/X sky130_fd_sc_hd__o22a_1
X_4496_ _9783_/Q _4493_/A _8844_/X _4493_/Y VGND VGND VPWR VPWR _9783_/D sky130_fd_sc_hd__a22o_1
XFILLER_103_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6235_ _6230_/Y _5968_/B _6231_/Y _5110_/B _6234_/X VGND VGND VPWR VPWR _6236_/D
+ sky130_fd_sc_hd__o221a_1
X_6166_ input69/X _8955_/S input50/X _8926_/S VGND VGND VPWR VPWR _6166_/Y sky130_fd_sc_hd__a22oi_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6097_ _6097_/A VGND VGND VPWR VPWR _6097_/Y sky130_fd_sc_hd__clkinv_2
X_5117_ _9635_/Q _5112_/A _5964_/B1 _5112_/Y VGND VGND VPWR VPWR _9635_/D sky130_fd_sc_hd__a22o_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5048_ _9674_/Q _5047_/A _8846_/X _5047_/Y VGND VGND VPWR VPWR _9674_/D sky130_fd_sc_hd__a22o_1
XFILLER_150_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8807_ _8807_/A _8807_/B VGND VGND VPWR VPWR _8807_/Y sky130_fd_sc_hd__nor2_2
X_9787_ _9790_/CLK _9787_/D _9757_/SET_B VGND VGND VPWR VPWR _9787_/Q sky130_fd_sc_hd__dfrtp_4
X_8738_ _8738_/A VGND VGND VPWR VPWR _8738_/Y sky130_fd_sc_hd__inv_2
X_6999_ _6999_/A VGND VGND VPWR VPWR _6999_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8669_ _8713_/A _8703_/D _8706_/B VGND VGND VPWR VPWR _8670_/C sky130_fd_sc_hd__or3_1
XFILLER_193_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6020_ _6040_/A VGND VGND VPWR VPWR _6021_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_100_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7971_ _7971_/A _8098_/A VGND VGND VPWR VPWR _8116_/A sky130_fd_sc_hd__or2_1
XFILLER_94_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6922_ _9121_/Q VGND VGND VPWR VPWR _6922_/Y sky130_fd_sc_hd__clkinv_2
X_9710_ _9709_/CLK _9710_/D _4939_/X VGND VGND VPWR VPWR _9710_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_47_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6853_ _9451_/Q VGND VGND VPWR VPWR _6853_/Y sky130_fd_sc_hd__inv_2
X_9641_ _9774_/CLK _9641_/D _7011_/B VGND VGND VPWR VPWR _9641_/Q sky130_fd_sc_hd__dfrtp_1
X_5804_ _9207_/Q _5799_/A _8842_/X _5799_/Y VGND VGND VPWR VPWR _9207_/D sky130_fd_sc_hd__a22o_1
XFILLER_62_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9572_ _9788_/CLK _9572_/D _9646_/SET_B VGND VGND VPWR VPWR _9572_/Q sky130_fd_sc_hd__dfrtp_2
X_6784_ _6784_/A _6784_/B _6784_/C _6784_/D VGND VGND VPWR VPWR _6785_/C sky130_fd_sc_hd__and4_1
XFILLER_22_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8523_ _8523_/A VGND VGND VPWR VPWR _8523_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5735_ _9246_/Q _9245_/Q _9055_/Q _9247_/Q VGND VGND VPWR VPWR _5735_/X sky130_fd_sc_hd__a31o_1
X_5666_ _9273_/Q _5662_/A _8925_/A1 _5662_/Y VGND VGND VPWR VPWR _9273_/D sky130_fd_sc_hd__a22o_1
XFILLER_129_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8454_ _8454_/A _8454_/B VGND VGND VPWR VPWR _8455_/B sky130_fd_sc_hd__nand2_1
XFILLER_163_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7405_ _7405_/A VGND VGND VPWR VPWR _7405_/X sky130_fd_sc_hd__buf_6
X_4617_ _9724_/Q _4615_/A _5964_/B1 _4615_/Y VGND VGND VPWR VPWR _9724_/D sky130_fd_sc_hd__a22o_1
X_8385_ _8650_/C _8385_/B VGND VGND VPWR VPWR _8436_/A sky130_fd_sc_hd__or2_1
X_5597_ _9311_/Q _5596_/A _8843_/X _5596_/Y VGND VGND VPWR VPWR _9311_/D sky130_fd_sc_hd__a22o_1
XFILLER_190_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4548_ _4548_/A VGND VGND VPWR VPWR _8975_/S sky130_fd_sc_hd__buf_12
XFILLER_150_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7336_ _6682_/Y _7048_/B _6772_/Y _7077_/A _7335_/X VGND VGND VPWR VPWR _7343_/A
+ sky130_fd_sc_hd__o221a_2
X_7267_ _6139_/Y _7077_/C _6133_/Y _7077_/D _7266_/X VGND VGND VPWR VPWR _7267_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_104_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4479_ _4729_/A _4729_/B _4669_/A _8932_/X VGND VGND VPWR VPWR _4931_/A sky130_fd_sc_hd__or4_4
X_9006_ _9599_/Q _8789_/A VGND VGND VPWR VPWR mgmt_gpio_out[29] sky130_fd_sc_hd__ebufn_8
XFILLER_89_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6218_ _9112_/Q VGND VGND VPWR VPWR _6218_/Y sky130_fd_sc_hd__clkinv_4
X_7198_ _7198_/A _7198_/B _7198_/C _7198_/D VGND VGND VPWR VPWR _7199_/C sky130_fd_sc_hd__and4_1
X_6149_ _6149_/A VGND VGND VPWR VPWR _6149_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_97_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5520_ _5520_/A VGND VGND VPWR VPWR _5520_/Y sky130_fd_sc_hd__inv_2
XFILLER_157_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5451_ _5451_/A VGND VGND VPWR VPWR _5452_/A sky130_fd_sc_hd__buf_2
XFILLER_172_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5382_ _5545_/A _5382_/B VGND VGND VPWR VPWR _5383_/A sky130_fd_sc_hd__or2_1
X_8170_ _8170_/A _8389_/A VGND VGND VPWR VPWR _8396_/A sky130_fd_sc_hd__or2_1
XFILLER_160_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7121_ _7121_/A _7392_/B VGND VGND VPWR VPWR _7121_/X sky130_fd_sc_hd__or2_1
XFILLER_99_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7052_ _7075_/A _7085_/B VGND VGND VPWR VPWR _7053_/A sky130_fd_sc_hd__or2_1
XFILLER_140_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6003_ _6040_/A VGND VGND VPWR VPWR _6004_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_67_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7954_ _7954_/A VGND VGND VPWR VPWR _8164_/A sky130_fd_sc_hd__buf_12
XFILLER_82_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6905_ _9391_/Q VGND VGND VPWR VPWR _6905_/Y sky130_fd_sc_hd__clkinv_2
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7885_ _8515_/B _7885_/B VGND VGND VPWR VPWR _7885_/X sky130_fd_sc_hd__or2_1
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6836_ _6831_/Y _4822_/X _6832_/Y _5278_/B _6835_/X VGND VGND VPWR VPWR _6878_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9624_ _9674_/CLK _9624_/D _9633_/SET_B VGND VGND VPWR VPWR _9624_/Q sky130_fd_sc_hd__dfrtp_1
X_9555_ _9758_/CLK _9555_/D _7011_/B VGND VGND VPWR VPWR _9555_/Q sky130_fd_sc_hd__dfrtp_1
X_6767_ _9400_/Q VGND VGND VPWR VPWR _6767_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8506_ _8615_/A _8506_/B _8506_/C VGND VGND VPWR VPWR _8693_/A sky130_fd_sc_hd__or3_2
X_5718_ _9245_/Q VGND VGND VPWR VPWR _5738_/B sky130_fd_sc_hd__inv_2
X_6698_ _9078_/Q VGND VGND VPWR VPWR _6698_/Y sky130_fd_sc_hd__clkinv_2
X_9486_ _9777_/CLK _9486_/D _7011_/B VGND VGND VPWR VPWR _9486_/Q sky130_fd_sc_hd__dfstp_1
X_8437_ _8632_/A _8437_/B VGND VGND VPWR VPWR _8704_/B sky130_fd_sc_hd__nor2_1
X_5649_ _5649_/A _5649_/B _9278_/Q _9277_/Q VGND VGND VPWR VPWR _6997_/C sky130_fd_sc_hd__or4_1
XFILLER_156_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8368_ _8368_/A _8577_/C _8675_/A _8578_/C VGND VGND VPWR VPWR _8372_/A sky130_fd_sc_hd__or4_2
XFILLER_163_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7319_ _6932_/Y _7068_/A _6805_/Y _7105_/X VGND VGND VPWR VPWR _7319_/X sky130_fd_sc_hd__o22a_1
XFILLER_49_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8299_ _8299_/A _8299_/B VGND VGND VPWR VPWR _8300_/B sky130_fd_sc_hd__nor2_1
XFILLER_104_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_123 _7015_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_112 input86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_101 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_134 _7626_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_156 _8544_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_145 _5355_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_167 _8822_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_189 _6158_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_178 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_1_1_1_csclk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_127_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput7 mask_rev_in[12] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4951_ _9048_/Q _4951_/B VGND VGND VPWR VPWR _4951_/Y sky130_fd_sc_hd__nand2_1
XFILLER_24_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7670_ _6516_/Y _7425_/X _7667_/X _7669_/X VGND VGND VPWR VPWR _7680_/C sky130_fd_sc_hd__o211a_1
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4882_ _9773_/Q VGND VGND VPWR VPWR _4882_/Y sky130_fd_sc_hd__inv_2
X_6621_ _9765_/Q VGND VGND VPWR VPWR _6621_/Y sky130_fd_sc_hd__clkinv_2
X_9340_ _9535_/CLK _9340_/D _9528_/SET_B VGND VGND VPWR VPWR _9340_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6552_ _6552_/A VGND VGND VPWR VPWR _6552_/Y sky130_fd_sc_hd__inv_2
XFILLER_173_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6483_ _9297_/Q VGND VGND VPWR VPWR _8761_/A sky130_fd_sc_hd__inv_6
X_9271_ _9535_/CLK _9271_/D _9528_/SET_B VGND VGND VPWR VPWR _9271_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_145_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5503_ _9375_/Q _5498_/A _8929_/A1 _5498_/Y VGND VGND VPWR VPWR _9375_/D sky130_fd_sc_hd__a22o_1
XFILLER_9_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5434_ _9423_/Q _5433_/A _8846_/X _5433_/Y VGND VGND VPWR VPWR _9423_/D sky130_fd_sc_hd__a22o_1
XFILLER_145_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8222_ _8341_/A _8498_/A _8640_/A VGND VGND VPWR VPWR _8223_/B sky130_fd_sc_hd__or3_1
XFILLER_118_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput300 _9741_/Q VGND VGND VPWR VPWR pll_trim[9] sky130_fd_sc_hd__buf_2
Xoutput344 _9036_/Q VGND VGND VPWR VPWR wb_dat_o[24] sky130_fd_sc_hd__buf_2
Xoutput333 _9018_/Q VGND VGND VPWR VPWR wb_dat_o[14] sky130_fd_sc_hd__buf_2
XFILLER_133_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8153_ _8552_/A _8378_/B VGND VGND VPWR VPWR _8367_/A sky130_fd_sc_hd__nor2_1
Xoutput322 _9767_/Q VGND VGND VPWR VPWR sram_ro_addr[5] sky130_fd_sc_hd__buf_2
Xoutput311 _8821_/X VGND VGND VPWR VPWR serial_resetn sky130_fd_sc_hd__buf_2
XFILLER_160_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5365_ _9468_/Q _5357_/A _8839_/X _5357_/Y VGND VGND VPWR VPWR _9468_/D sky130_fd_sc_hd__a22o_1
Xoutput355 _9025_/Q VGND VGND VPWR VPWR wb_dat_o[5] sky130_fd_sc_hd__buf_2
X_7104_ _7104_/A _7127_/B _7127_/C VGND VGND VPWR VPWR _7105_/A sky130_fd_sc_hd__or3_1
X_8084_ _8084_/A _8521_/B VGND VGND VPWR VPWR _8538_/D sky130_fd_sc_hd__or2_1
XFILLER_113_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5296_ _9516_/Q _5292_/A _5966_/B1 _5292_/Y VGND VGND VPWR VPWR _9516_/D sky130_fd_sc_hd__a22o_1
XFILLER_87_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7035_ _7115_/B _7073_/C VGND VGND VPWR VPWR _7036_/A sky130_fd_sc_hd__or2_1
XFILLER_142_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8986_ _8986_/A _8749_/A VGND VGND VPWR VPWR mgmt_gpio_out[9] sky130_fd_sc_hd__ebufn_2
XFILLER_70_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7937_ _8282_/C _7836_/C _8282_/B _8703_/A _7936_/X VGND VGND VPWR VPWR _7938_/B
+ sky130_fd_sc_hd__a311oi_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7868_ _7868_/A VGND VGND VPWR VPWR _8316_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_42_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_0_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_3_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9607_ _9617_/CLK _9607_/D _9295_/SET_B VGND VGND VPWR VPWR _9607_/Q sky130_fd_sc_hd__dfrtp_1
X_6819_ _9417_/Q VGND VGND VPWR VPWR _6819_/Y sky130_fd_sc_hd__inv_4
XFILLER_11_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7799_ _8394_/C VGND VGND VPWR VPWR _8379_/C sky130_fd_sc_hd__inv_6
XFILLER_11_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9538_ _9768_/CLK _9538_/D _4628_/A VGND VGND VPWR VPWR _9538_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9469_ _9684_/CLK _9469_/D _9685_/SET_B VGND VGND VPWR VPWR _9469_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_167_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5150_ _9615_/Q _5147_/A _8844_/X _5147_/Y VGND VGND VPWR VPWR _9615_/D sky130_fd_sc_hd__a22o_1
XFILLER_69_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5081_ _5081_/A VGND VGND VPWR VPWR _5082_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_96_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8840_ _9701_/Q _9660_/Q _9587_/Q VGND VGND VPWR VPWR _8840_/X sky130_fd_sc_hd__mux2_8
XFILLER_64_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8771_ _8771_/A VGND VGND VPWR VPWR _8772_/A sky130_fd_sc_hd__clkbuf_1
X_5983_ _6040_/A VGND VGND VPWR VPWR _5984_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_25_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4934_ _4934_/A _4934_/B _4934_/C _4934_/D VGND VGND VPWR VPWR _4935_/D sky130_fd_sc_hd__and4_1
XFILLER_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7722_ _9088_/Q _7722_/B VGND VGND VPWR VPWR _7722_/Y sky130_fd_sc_hd__nand2_1
XFILLER_177_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7653_ _6695_/Y _7445_/X _6700_/Y _7447_/X VGND VGND VPWR VPWR _7653_/X sky130_fd_sc_hd__o22a_1
XANTENNA_23 _4481_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4865_ _9484_/Q VGND VGND VPWR VPWR _4865_/Y sky130_fd_sc_hd__clkinv_4
XANTENNA_12 _7353_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_34 _5278_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7584_ _6175_/Y _7451_/X _6159_/Y _7453_/X _7583_/X VGND VGND VPWR VPWR _7589_/B
+ sky130_fd_sc_hd__o221a_1
XANTENNA_56 _6716_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_45 _6271_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4796_ _6111_/A _4903_/B VGND VGND VPWR VPWR _5121_/B sky130_fd_sc_hd__or2_4
X_6604_ _9492_/Q VGND VGND VPWR VPWR _6604_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_192_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9323_ _9613_/CLK _9323_/D _9646_/SET_B VGND VGND VPWR VPWR _9323_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_118_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_78 _9571_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_67 _7330_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_89 _6505_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6535_ _6533_/Y _5080_/B _6534_/Y _6052_/C VGND VGND VPWR VPWR _6535_/X sky130_fd_sc_hd__o22a_1
XFILLER_137_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9254_ _9681_/CLK _9254_/D _9633_/SET_B VGND VGND VPWR VPWR _9254_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_173_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8205_ _8510_/A _8305_/B _8226_/C VGND VGND VPWR VPWR _8595_/B sky130_fd_sc_hd__nor3_2
X_6466_ _6461_/Y _5545_/B _6462_/Y _5013_/B _6465_/X VGND VGND VPWR VPWR _6473_/C
+ sky130_fd_sc_hd__o221a_1
X_5417_ _9434_/Q _5414_/A _5965_/B1 _5414_/Y VGND VGND VPWR VPWR _9434_/D sky130_fd_sc_hd__a22o_1
X_6397_ _9514_/Q VGND VGND VPWR VPWR _6397_/Y sky130_fd_sc_hd__inv_2
X_9185_ _9655_/CLK _9185_/D _9633_/SET_B VGND VGND VPWR VPWR _9185_/Q sky130_fd_sc_hd__dfrtp_1
X_5348_ _9482_/Q _5346_/A _8845_/X _5346_/Y VGND VGND VPWR VPWR _9482_/D sky130_fd_sc_hd__a22o_1
XFILLER_121_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8136_ _8136_/A _8358_/A _8642_/A _8359_/A VGND VGND VPWR VPWR _8140_/A sky130_fd_sc_hd__or4_1
X_8067_ _8067_/A _8539_/A VGND VGND VPWR VPWR _8069_/A sky130_fd_sc_hd__nor2_1
X_5279_ _5279_/A VGND VGND VPWR VPWR _5280_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_101_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7018_ _9626_/Q _7018_/B VGND VGND VPWR VPWR _7019_/A sky130_fd_sc_hd__and2b_1
XFILLER_46_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8969_ _8296_/Y _7944_/X _8975_/S VGND VGND VPWR VPWR _8969_/X sky130_fd_sc_hd__mux2_4
XFILLER_102_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4650_ _4994_/A VGND VGND VPWR VPWR _4651_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_174_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput10 mask_rev_in[15] VGND VGND VPWR VPWR _6085_/A sky130_fd_sc_hd__clkbuf_1
Xinput21 mask_rev_in[25] VGND VGND VPWR VPWR _6831_/A sky130_fd_sc_hd__clkbuf_1
Xinput54 mgmt_gpio_in[26] VGND VGND VPWR VPWR _6680_/A sky130_fd_sc_hd__clkbuf_1
Xinput43 mgmt_gpio_in[16] VGND VGND VPWR VPWR _4754_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_162_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6320_ _9325_/Q VGND VGND VPWR VPWR _6320_/Y sky130_fd_sc_hd__clkinv_2
X_4581_ _9746_/Q _4579_/A _8845_/X _4579_/Y VGND VGND VPWR VPWR _9746_/D sky130_fd_sc_hd__a22o_1
Xinput32 mask_rev_in[6] VGND VGND VPWR VPWR _6153_/A sky130_fd_sc_hd__clkbuf_1
Xinput65 mgmt_gpio_in[36] VGND VGND VPWR VPWR _8817_/A sky130_fd_sc_hd__buf_4
Xinput87 spimemio_flash_io1_do VGND VGND VPWR VPWR _8816_/A sky130_fd_sc_hd__buf_6
XFILLER_155_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput76 qspi_enabled VGND VGND VPWR VPWR _8835_/S sky130_fd_sc_hd__buf_6
Xinput98 sram_ro_data[14] VGND VGND VPWR VPWR _6221_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_170_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6251_ _6251_/A VGND VGND VPWR VPWR _6251_/Y sky130_fd_sc_hd__inv_4
XFILLER_170_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5202_ _6134_/A _6322_/A _5259_/A _8977_/X VGND VGND VPWR VPWR _5203_/A sky130_fd_sc_hd__a211o_4
XFILLER_115_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6182_ _9224_/Q VGND VGND VPWR VPWR _6182_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_69_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5133_ _5133_/A _8977_/S VGND VGND VPWR VPWR _5156_/B sky130_fd_sc_hd__or2_4
XFILLER_111_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5064_ _8968_/X _9666_/Q _5078_/S VGND VGND VPWR VPWR _5065_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8823_ _9150_/Q _9790_/Q _9787_/Q VGND VGND VPWR VPWR _8823_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8754_ _8754_/A VGND VGND VPWR VPWR _8754_/X sky130_fd_sc_hd__clkbuf_1
X_5966_ _9102_/Q _5962_/A _5966_/B1 _5962_/Y VGND VGND VPWR VPWR _9102_/D sky130_fd_sc_hd__a22o_1
XFILLER_178_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5897_ _5960_/A _5897_/B VGND VGND VPWR VPWR _5898_/A sky130_fd_sc_hd__or2_1
X_8685_ _8685_/A _8685_/B VGND VGND VPWR VPWR _8686_/B sky130_fd_sc_hd__or2_1
XFILLER_40_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7705_ _7705_/A VGND VGND VPWR VPWR _7706_/A sky130_fd_sc_hd__clkbuf_1
X_4917_ _4917_/A _4931_/B VGND VGND VPWR VPWR _5382_/B sky130_fd_sc_hd__or2_4
XFILLER_193_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4848_ _9411_/Q VGND VGND VPWR VPWR _4848_/Y sky130_fd_sc_hd__clkinv_2
X_7636_ _6935_/Y _7441_/X _6824_/Y _7443_/X _7635_/X VGND VGND VPWR VPWR _7643_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4779_ _9231_/Q VGND VGND VPWR VPWR _4779_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_148_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7567_ _6288_/Y _7465_/X _6244_/Y _7467_/X VGND VGND VPWR VPWR _7567_/X sky130_fd_sc_hd__o22a_1
X_9306_ _9440_/CLK _9306_/D _9685_/SET_B VGND VGND VPWR VPWR _9306_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_134_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7498_ _6889_/Y _7471_/X _7150_/A _7473_/X _7497_/X VGND VGND VPWR VPWR _7499_/D
+ sky130_fd_sc_hd__o221a_1
X_6518_ _6516_/Y _5960_/B _6517_/Y _5089_/B VGND VGND VPWR VPWR _6518_/X sky130_fd_sc_hd__o22a_1
XFILLER_180_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9237_ _9596_/CLK _9237_/D _9528_/SET_B VGND VGND VPWR VPWR _9237_/Q sky130_fd_sc_hd__dfrtp_1
X_6449_ _9736_/Q VGND VGND VPWR VPWR _6449_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_161_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9168_ _9203_/CLK _9168_/D _9633_/SET_B VGND VGND VPWR VPWR _9168_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_40_csclk clkbuf_2_1_0_csclk/X VGND VGND VPWR VPWR _9785_/CLK sky130_fd_sc_hd__clkbuf_16
X_8119_ _8119_/A VGND VGND VPWR VPWR _8546_/A sky130_fd_sc_hd__inv_2
X_9099_ _9344_/CLK _9099_/D _9647_/SET_B VGND VGND VPWR VPWR _9099_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_0_0_csclk clkbuf_2_1_0_csclk/A VGND VGND VPWR VPWR _9329_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_57_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5820_ _5820_/A VGND VGND VPWR VPWR _5820_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5751_ _9280_/Q _9279_/Q _5751_/C _9277_/Q VGND VGND VPWR VPWR _5753_/B sky130_fd_sc_hd__or4_2
XFILLER_34_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8470_ _8470_/A _8470_/B _8698_/A VGND VGND VPWR VPWR _8474_/A sky130_fd_sc_hd__or3_1
X_4702_ _4917_/A _4843_/B VGND VGND VPWR VPWR _5013_/B sky130_fd_sc_hd__or2_4
X_5682_ _9263_/Q _5681_/A _8846_/X _5681_/Y VGND VGND VPWR VPWR _9263_/D sky130_fd_sc_hd__a22o_1
XFILLER_147_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7421_ _7421_/A VGND VGND VPWR VPWR _7421_/X sky130_fd_sc_hd__buf_6
XFILLER_163_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4633_ _9050_/Q VGND VGND VPWR VPWR _4964_/B sky130_fd_sc_hd__inv_2
XFILLER_162_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7352_ _7352_/A _7352_/B _7352_/C _7352_/D VGND VGND VPWR VPWR _7353_/C sky130_fd_sc_hd__and4_1
X_4564_ _5960_/A _4564_/B VGND VGND VPWR VPWR _4565_/A sky130_fd_sc_hd__or2_1
XFILLER_143_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6303_ _9098_/Q VGND VGND VPWR VPWR _6303_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_116_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7283_ _6072_/Y _5728_/X _6059_/Y _7040_/A _7282_/X VGND VGND VPWR VPWR _7286_/C
+ sky130_fd_sc_hd__o221a_1
X_9022_ _9027_/CLK _9022_/D VGND VGND VPWR VPWR _9022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4495_ _9784_/Q _4493_/A _8845_/X _4493_/Y VGND VGND VPWR VPWR _9784_/D sky130_fd_sc_hd__a22o_1
X_6234_ _6232_/Y _5045_/B _6233_/Y _4861_/X VGND VGND VPWR VPWR _6234_/X sky130_fd_sc_hd__o22a_1
XFILLER_97_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6165_ _6165_/A VGND VGND VPWR VPWR _8955_/S sky130_fd_sc_hd__clkinv_8
X_6096_ _6096_/A _6096_/B _6096_/C _6096_/D VGND VGND VPWR VPWR _6145_/B sky130_fd_sc_hd__and4_2
X_5116_ _9636_/Q _5112_/A _5963_/B1 _5112_/Y VGND VGND VPWR VPWR _9636_/D sky130_fd_sc_hd__a22o_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5047_ _5047_/A VGND VGND VPWR VPWR _5047_/Y sky130_fd_sc_hd__inv_2
XFILLER_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9786_ _9788_/CLK _9786_/D _9295_/SET_B VGND VGND VPWR VPWR _9786_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_80_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8806_ _8806_/A VGND VGND VPWR VPWR _8806_/X sky130_fd_sc_hd__clkbuf_1
X_6998_ _5691_/A _6991_/Y _6996_/Y _6999_/A VGND VGND VPWR VPWR _9055_/D sky130_fd_sc_hd__o22ai_1
XFILLER_159_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5949_ _6052_/A _5949_/B VGND VGND VPWR VPWR _5950_/A sky130_fd_sc_hd__or2_1
X_8737_ _8137_/B _8554_/B _8736_/X _8628_/X VGND VGND VPWR VPWR _8737_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_13_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8668_ _8668_/A _8668_/B _8668_/C _8668_/D VGND VGND VPWR VPWR _8699_/D sky130_fd_sc_hd__or4_4
XFILLER_21_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8599_ _8599_/A _8599_/B _8599_/C _8599_/D VGND VGND VPWR VPWR _8696_/A sky130_fd_sc_hd__or4_4
X_7619_ _4660_/Y _7455_/X _4823_/Y _7457_/X VGND VGND VPWR VPWR _7619_/X sky130_fd_sc_hd__o22a_1
XFILLER_181_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput200 wb_sel_i[2] VGND VGND VPWR VPWR _7733_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7970_ _7970_/A VGND VGND VPWR VPWR _8098_/A sky130_fd_sc_hd__buf_6
XFILLER_94_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6921_ _9689_/Q VGND VGND VPWR VPWR _6921_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9640_ _4450_/A1 _9640_/D _6146_/A VGND VGND VPWR VPWR _9640_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_120_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6852_ _6843_/Y _5328_/B _6846_/X _6851_/X VGND VGND VPWR VPWR _6878_/C sky130_fd_sc_hd__o211a_1
X_5803_ _9208_/Q _5799_/A _8925_/A1 _5799_/Y VGND VGND VPWR VPWR _9208_/D sky130_fd_sc_hd__a22o_1
X_9571_ _9613_/CLK _9571_/D _9646_/SET_B VGND VGND VPWR VPWR _9571_/Q sky130_fd_sc_hd__dfrtp_1
X_8522_ _8064_/C _8064_/B _8521_/Y _8016_/B VGND VGND VPWR VPWR _8527_/B sky130_fd_sc_hd__a31o_1
X_6783_ _6783_/A _6783_/B _6783_/C _6783_/D VGND VGND VPWR VPWR _6784_/D sky130_fd_sc_hd__and4_2
XFILLER_50_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5734_ _7037_/A _5731_/Y _5724_/B _7096_/B VGND VGND VPWR VPWR _9248_/D sky130_fd_sc_hd__o22ai_1
XFILLER_50_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5665_ _9274_/Q _5662_/A _8844_/X _5662_/Y VGND VGND VPWR VPWR _9274_/D sky130_fd_sc_hd__a22o_1
XFILLER_129_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8453_ _8665_/A _8453_/B _8453_/C _8607_/C VGND VGND VPWR VPWR _8455_/A sky130_fd_sc_hd__or4_1
XFILLER_30_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8384_ _8384_/A _8651_/B VGND VGND VPWR VPWR _8385_/B sky130_fd_sc_hd__nor2_1
XFILLER_148_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7404_ _7466_/A _7476_/C _9255_/Q VGND VGND VPWR VPWR _7405_/A sky130_fd_sc_hd__or3_1
X_4616_ _9725_/Q _4615_/A _5963_/B1 _4615_/Y VGND VGND VPWR VPWR _9725_/D sky130_fd_sc_hd__a22o_1
XFILLER_190_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5596_ _5596_/A VGND VGND VPWR VPWR _5596_/Y sky130_fd_sc_hd__inv_2
X_7335_ _6732_/Y _7040_/C _6743_/Y _7059_/C VGND VGND VPWR VPWR _7335_/X sky130_fd_sc_hd__o22a_1
X_4547_ _8810_/A _8812_/A _8813_/A VGND VGND VPWR VPWR _4548_/A sky130_fd_sc_hd__and3_1
XFILLER_116_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7266_ _6113_/Y _7086_/X _6074_/Y _7088_/X VGND VGND VPWR VPWR _7266_/X sky130_fd_sc_hd__o22a_1
X_4478_ _4478_/A VGND VGND VPWR VPWR _9789_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9005_ _9598_/Q _8787_/A VGND VGND VPWR VPWR mgmt_gpio_out[28] sky130_fd_sc_hd__ebufn_8
XFILLER_131_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7197_ _8769_/A _7124_/X _6485_/Y _7068_/B _7196_/X VGND VGND VPWR VPWR _7198_/D
+ sky130_fd_sc_hd__o221a_1
X_6217_ _6212_/Y _5872_/B _6213_/Y _6251_/A _6216_/X VGND VGND VPWR VPWR _6236_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_58_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6148_ _6148_/A VGND VGND VPWR VPWR _6149_/A sky130_fd_sc_hd__clkbuf_4
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6079_ _9527_/Q VGND VGND VPWR VPWR _6079_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_73_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9769_ _9769_/CLK _9769_/D _4628_/A VGND VGND VPWR VPWR _9769_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_110_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5450_ _5671_/A _5450_/B VGND VGND VPWR VPWR _5451_/A sky130_fd_sc_hd__or2_1
XFILLER_145_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5381_ _9458_/Q _5376_/A _8839_/X _5376_/Y VGND VGND VPWR VPWR _9458_/D sky130_fd_sc_hd__a22o_1
XFILLER_125_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7120_ _4687_/Y _7059_/D _4877_/Y _7116_/X _7119_/X VGND VGND VPWR VPWR _7131_/B
+ sky130_fd_sc_hd__o221a_1
Xclkbuf_3_2_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A VGND VGND VPWR VPWR _9280_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_140_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7051_ _9248_/Q _7056_/B _7127_/A VGND VGND VPWR VPWR _7085_/B sky130_fd_sc_hd__or3_1
XFILLER_101_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6002_ _9087_/Q _5995_/A _8912_/X _5995_/Y VGND VGND VPWR VPWR _9087_/D sky130_fd_sc_hd__a22o_1
XFILLER_27_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7953_ _8195_/A _8632_/A VGND VGND VPWR VPWR _7954_/A sky130_fd_sc_hd__or2_1
X_6904_ _9355_/Q VGND VGND VPWR VPWR _6904_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7884_ _7903_/C _8193_/A _8583_/A VGND VGND VPWR VPWR _7885_/B sky130_fd_sc_hd__or3_2
XFILLER_23_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6835_ _6833_/Y _5100_/B _6834_/Y _4590_/B VGND VGND VPWR VPWR _6835_/X sky130_fd_sc_hd__o22a_1
X_9623_ _9674_/CLK _9623_/D _9633_/SET_B VGND VGND VPWR VPWR _9623_/Q sky130_fd_sc_hd__dfrtp_1
X_9554_ _9755_/CLK _9554_/D _9633_/SET_B VGND VGND VPWR VPWR _9554_/Q sky130_fd_sc_hd__dfrtp_1
X_6766_ _6766_/A VGND VGND VPWR VPWR _6766_/Y sky130_fd_sc_hd__inv_2
XFILLER_148_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8505_ _8597_/D _8599_/D _8657_/C _8504_/X VGND VGND VPWR VPWR _8509_/A sky130_fd_sc_hd__or4b_4
XFILLER_10_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5717_ _9246_/Q VGND VGND VPWR VPWR _5737_/A sky130_fd_sc_hd__inv_2
XFILLER_136_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6697_ _6692_/Y _4491_/B _6693_/Y _5545_/B _6696_/X VGND VGND VPWR VPWR _6716_/A
+ sky130_fd_sc_hd__o221a_1
X_9485_ _9774_/CLK _9485_/D _7011_/B VGND VGND VPWR VPWR _9485_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_40_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8436_ _8436_/A _8436_/B VGND VGND VPWR VPWR _8487_/A sky130_fd_sc_hd__nand2_1
X_5648_ _9280_/Q VGND VGND VPWR VPWR _5649_/A sky130_fd_sc_hd__inv_2
XFILLER_40_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5579_ _9323_/Q _5574_/A _8929_/A1 _5574_/Y VGND VGND VPWR VPWR _9323_/D sky130_fd_sc_hd__a22o_1
X_8367_ _8367_/A _8367_/B VGND VGND VPWR VPWR _8578_/C sky130_fd_sc_hd__or2_1
X_8298_ _8298_/A VGND VGND VPWR VPWR _8600_/A sky130_fd_sc_hd__inv_2
X_7318_ _6802_/Y _7059_/B _6840_/Y _7068_/C _7317_/X VGND VGND VPWR VPWR _7321_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_2_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7249_ _6169_/Y _7097_/X _6168_/Y _7099_/X VGND VGND VPWR VPWR _7249_/X sky130_fd_sc_hd__o22a_1
XFILLER_49_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_124 _7015_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_113 input86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_102 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_157 _8765_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_146 _6356_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_135 _7626_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_179 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_168 _7021_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput8 mask_rev_in[13] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4950_ _9092_/Q _9091_/Q _6022_/C VGND VGND VPWR VPWR _4951_/B sky130_fd_sc_hd__and3_1
X_4881_ _4874_/Y _4602_/B _4875_/Y _5110_/B _4880_/X VGND VGND VPWR VPWR _4896_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_51_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6620_ _6615_/Y _5336_/B _8793_/A _5393_/B _6619_/X VGND VGND VPWR VPWR _6627_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_158_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6551_ _9644_/Q VGND VGND VPWR VPWR _6551_/Y sky130_fd_sc_hd__inv_2
X_5502_ _9376_/Q _5498_/A _8925_/A1 _5498_/Y VGND VGND VPWR VPWR _9376_/D sky130_fd_sc_hd__a22o_1
XFILLER_185_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9270_ _9535_/CLK _9270_/D _9528_/SET_B VGND VGND VPWR VPWR _9270_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_118_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6482_ _6477_/Y _5768_/B _8757_/A _5679_/B _6481_/X VGND VGND VPWR VPWR _6501_/A
+ sky130_fd_sc_hd__o221a_1
X_5433_ _5433_/A VGND VGND VPWR VPWR _5433_/Y sky130_fd_sc_hd__inv_2
XFILLER_173_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8221_ _8510_/A _8498_/A _8640_/A VGND VGND VPWR VPWR _8223_/A sky130_fd_sc_hd__or3_1
Xoutput301 _9044_/Q VGND VGND VPWR VPWR pwr_ctrl_out[0] sky130_fd_sc_hd__buf_2
X_5364_ _9469_/Q _5357_/A _8840_/X _5357_/Y VGND VGND VPWR VPWR _9469_/D sky130_fd_sc_hd__a22o_1
Xoutput334 _9019_/Q VGND VGND VPWR VPWR wb_dat_o[15] sky130_fd_sc_hd__buf_2
Xoutput312 _8804_/X VGND VGND VPWR VPWR spi_sdi sky130_fd_sc_hd__buf_2
X_8152_ _8152_/A _8674_/A VGND VGND VPWR VPWR _8154_/A sky130_fd_sc_hd__or2_1
Xoutput323 _9768_/Q VGND VGND VPWR VPWR sram_ro_addr[6] sky130_fd_sc_hd__buf_2
Xoutput345 _9037_/Q VGND VGND VPWR VPWR wb_dat_o[25] sky130_fd_sc_hd__buf_2
X_7103_ _4732_/Y _7059_/B _4744_/Y _7068_/C _7102_/X VGND VGND VPWR VPWR _7108_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_126_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput356 _9026_/Q VGND VGND VPWR VPWR wb_dat_o[6] sky130_fd_sc_hd__buf_2
X_8083_ _8185_/A _8187_/A _8083_/C VGND VGND VPWR VPWR _8086_/A sky130_fd_sc_hd__and3_1
X_5295_ _9517_/Q _5292_/A _5965_/B1 _5292_/Y VGND VGND VPWR VPWR _9517_/D sky130_fd_sc_hd__a22o_1
XFILLER_87_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7034_ _7125_/A _7111_/C VGND VGND VPWR VPWR _7115_/B sky130_fd_sc_hd__or2_1
XFILLER_95_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8985_ _8985_/A _8747_/A VGND VGND VPWR VPWR mgmt_gpio_out[8] sky130_fd_sc_hd__ebufn_8
XFILLER_55_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7936_ _8476_/A _7936_/B VGND VGND VPWR VPWR _7936_/X sky130_fd_sc_hd__or2_1
XFILLER_70_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7867_ _7959_/A _8528_/A _8583_/A _7894_/B VGND VGND VPWR VPWR _7868_/A sky130_fd_sc_hd__or4_4
X_9606_ _9617_/CLK _9606_/D _9295_/SET_B VGND VGND VPWR VPWR _9606_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_143_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6818_ _9443_/Q VGND VGND VPWR VPWR _6818_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_168_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7798_ _8510_/A _8188_/B VGND VGND VPWR VPWR _8651_/A sky130_fd_sc_hd__nor2_2
XFILLER_149_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6749_ _9046_/Q VGND VGND VPWR VPWR _6749_/Y sky130_fd_sc_hd__clkinv_4
X_9537_ _9768_/CLK _9537_/D _4628_/A VGND VGND VPWR VPWR _9537_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9468_ _9535_/CLK _9468_/D _9528_/SET_B VGND VGND VPWR VPWR _9468_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_191_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8419_ _8552_/A _8401_/B _8415_/X _8418_/Y VGND VGND VPWR VPWR _8419_/X sky130_fd_sc_hd__o211a_1
XFILLER_151_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9399_ _9758_/CLK _9399_/D _7011_/B VGND VGND VPWR VPWR _9399_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_151_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8815__379 VGND VGND VPWR VPWR _9057_/D _8815__379/LO sky130_fd_sc_hd__conb_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5080_ _5259_/A _5080_/B VGND VGND VPWR VPWR _5081_/A sky130_fd_sc_hd__or2_1
XFILLER_96_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8770_ _8770_/A VGND VGND VPWR VPWR _8770_/X sky130_fd_sc_hd__clkbuf_1
X_5982_ _9092_/Q _5981_/X _7008_/A _5985_/B VGND VGND VPWR VPWR _9092_/D sky130_fd_sc_hd__o22a_1
X_4933_ _4924_/Y _5366_/B _4926_/Y _5306_/B _4932_/X VGND VGND VPWR VPWR _4934_/D
+ sky130_fd_sc_hd__o221a_1
X_7721_ _7721_/A VGND VGND VPWR VPWR _7722_/B sky130_fd_sc_hd__inv_2
XANTENNA_13 _7397_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4864_ _4864_/A _4864_/B _4864_/C _4864_/D VGND VGND VPWR VPWR _4935_/B sky130_fd_sc_hd__and4_1
X_7652_ _6731_/Y _7425_/X _7649_/X _7651_/X VGND VGND VPWR VPWR _7662_/C sky130_fd_sc_hd__o211a_1
X_6603_ _9479_/Q VGND VGND VPWR VPWR _8775_/A sky130_fd_sc_hd__clkinv_8
XFILLER_177_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_24 _4481_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7583_ _6154_/Y _7455_/X _6157_/Y _7457_/X VGND VGND VPWR VPWR _7583_/X sky130_fd_sc_hd__o22a_1
XANTENNA_35 _4922_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_57 _6716_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4795_ _9627_/Q VGND VGND VPWR VPWR _4795_/Y sky130_fd_sc_hd__inv_2
XANTENNA_46 _6280_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9322_ _9352_/CLK _9322_/D _9646_/SET_B VGND VGND VPWR VPWR _9322_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_68 _7343_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6534_ _9047_/Q VGND VGND VPWR VPWR _6534_/Y sky130_fd_sc_hd__inv_2
XANTENNA_79 _8831_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6465_ _6463_/Y _5045_/B _6464_/Y _5080_/B VGND VGND VPWR VPWR _6465_/X sky130_fd_sc_hd__o22a_1
X_9253_ _9681_/CLK _9253_/D _9633_/SET_B VGND VGND VPWR VPWR _9253_/Q sky130_fd_sc_hd__dfrtp_2
X_8204_ _8204_/A _8640_/A VGND VGND VPWR VPWR _8678_/A sky130_fd_sc_hd__nor2_1
XFILLER_133_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5416_ _9435_/Q _5414_/A _5964_/B1 _5414_/Y VGND VGND VPWR VPWR _9435_/D sky130_fd_sc_hd__a22o_1
X_6396_ _9480_/Q VGND VGND VPWR VPWR _6396_/Y sky130_fd_sc_hd__clkinv_4
X_9184_ _9613_/CLK _9184_/D _9646_/SET_B VGND VGND VPWR VPWR _9184_/Q sky130_fd_sc_hd__dfrtp_1
X_5347_ _9483_/Q _5346_/A _8846_/X _5346_/Y VGND VGND VPWR VPWR _9483_/D sky130_fd_sc_hd__a22o_1
XFILLER_161_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8135_ _8137_/B _8378_/B VGND VGND VPWR VPWR _8359_/A sky130_fd_sc_hd__nor2_1
X_5278_ _5545_/A _5278_/B VGND VGND VPWR VPWR _5279_/A sky130_fd_sc_hd__or2_1
X_8066_ _8282_/B _8518_/A _8282_/C VGND VGND VPWR VPWR _8539_/A sky130_fd_sc_hd__and3_1
XFILLER_87_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7017_ _7017_/A VGND VGND VPWR VPWR _7017_/Y sky130_fd_sc_hd__inv_2
X_8968_ _7751_/X _8968_/A1 _8975_/S VGND VGND VPWR VPWR _8968_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7919_ _8521_/B _8254_/B VGND VGND VPWR VPWR _8320_/A sky130_fd_sc_hd__or2_1
XFILLER_168_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8899_ _7712_/X _9083_/Q _9051_/Q VGND VGND VPWR VPWR _8899_/X sky130_fd_sc_hd__mux2_1
XFILLER_168_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4580_ _9747_/Q _4579_/A _8846_/X _4579_/Y VGND VGND VPWR VPWR _9747_/D sky130_fd_sc_hd__a22o_1
Xinput11 mask_rev_in[16] VGND VGND VPWR VPWR _4906_/A sky130_fd_sc_hd__clkbuf_1
Xinput22 mask_rev_in[26] VGND VGND VPWR VPWR _6726_/A sky130_fd_sc_hd__clkbuf_1
Xinput55 mgmt_gpio_in[27] VGND VGND VPWR VPWR _6531_/A sky130_fd_sc_hd__clkbuf_1
Xinput44 mgmt_gpio_in[17] VGND VGND VPWR VPWR _6903_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_162_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput33 mask_rev_in[7] VGND VGND VPWR VPWR _6087_/A sky130_fd_sc_hd__clkbuf_1
Xinput66 mgmt_gpio_in[37] VGND VGND VPWR VPWR _8818_/A sky130_fd_sc_hd__buf_4
Xinput88 spimemio_flash_io1_oeb VGND VGND VPWR VPWR _7015_/B sky130_fd_sc_hd__buf_6
Xinput77 ser_tx VGND VGND VPWR VPWR input77/X sky130_fd_sc_hd__buf_4
XFILLER_115_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6250_ _9637_/Q VGND VGND VPWR VPWR _6250_/Y sky130_fd_sc_hd__inv_2
Xinput99 sram_ro_data[15] VGND VGND VPWR VPWR _6099_/A sky130_fd_sc_hd__clkbuf_1
X_6181_ _9300_/Q VGND VGND VPWR VPWR _7260_/A sky130_fd_sc_hd__inv_2
X_5201_ _9578_/Q _5193_/Y _8849_/X _5193_/A VGND VGND VPWR VPWR _9578_/D sky130_fd_sc_hd__o22a_1
X_5132_ _7022_/B VGND VGND VPWR VPWR _8977_/S sky130_fd_sc_hd__inv_8
X_5063_ _5063_/A VGND VGND VPWR VPWR _5078_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_123_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8822_ _9176_/Q _9079_/Q _9787_/Q VGND VGND VPWR VPWR _8822_/X sky130_fd_sc_hd__mux2_4
XFILLER_25_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8753_ _8753_/A VGND VGND VPWR VPWR _8754_/A sky130_fd_sc_hd__clkbuf_1
X_5965_ _9103_/Q _5962_/A _5965_/B1 _5962_/Y VGND VGND VPWR VPWR _9103_/D sky130_fd_sc_hd__a22o_1
XFILLER_40_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4916_ _9450_/Q VGND VGND VPWR VPWR _4916_/Y sky130_fd_sc_hd__inv_2
X_8684_ _8115_/Y _8625_/B _8405_/A _8683_/X _8629_/B VGND VGND VPWR VPWR _8689_/A
+ sky130_fd_sc_hd__a2111o_2
XFILLER_21_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5896_ _8924_/X _6997_/A _5895_/Y _5849_/A _9138_/Q VGND VGND VPWR VPWR _9138_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_52_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7704_ _7704_/A VGND VGND VPWR VPWR _7704_/X sky130_fd_sc_hd__clkbuf_1
X_4847_ _4876_/B _4931_/B VGND VGND VPWR VPWR _5267_/B sky130_fd_sc_hd__or2_4
X_7635_ _6867_/Y _7445_/X _6872_/Y _7447_/X VGND VGND VPWR VPWR _7635_/X sky130_fd_sc_hd__o22a_1
XFILLER_193_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4778_ _4769_/Y _5089_/B _4771_/Y _5583_/B _4777_/X VGND VGND VPWR VPWR _4790_/C
+ sky130_fd_sc_hd__o221a_1
X_7566_ _6298_/Y _7451_/X _6274_/Y _7453_/X _7565_/X VGND VGND VPWR VPWR _7571_/B
+ sky130_fd_sc_hd__o221a_1
X_9305_ _9440_/CLK _9305_/D _9685_/SET_B VGND VGND VPWR VPWR _9305_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6517_ _9649_/Q VGND VGND VPWR VPWR _6517_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7497_ _6823_/Y _7475_/X _6926_/Y _7477_/X VGND VGND VPWR VPWR _7497_/X sky130_fd_sc_hd__o22a_1
XFILLER_164_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9236_ _9371_/CLK _9236_/D _9295_/SET_B VGND VGND VPWR VPWR _9236_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_161_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6448_ _6434_/Y _5864_/B _6437_/X _6443_/X _6447_/X VGND VGND VPWR VPWR _6474_/C
+ sky130_fd_sc_hd__o2111a_1
XFILLER_134_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6379_ _9268_/Q VGND VGND VPWR VPWR _6379_/Y sky130_fd_sc_hd__clkinv_2
X_9167_ _9203_/CLK _9167_/D _9633_/SET_B VGND VGND VPWR VPWR _9167_/Q sky130_fd_sc_hd__dfrtp_1
X_8118_ _8394_/A _8379_/B _8117_/A VGND VGND VPWR VPWR _8118_/X sky130_fd_sc_hd__or3b_1
XFILLER_121_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9098_ _9344_/CLK _9098_/D _9647_/SET_B VGND VGND VPWR VPWR _9098_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8049_ _8097_/B _8554_/A _8048_/Y VGND VGND VPWR VPWR _8053_/A sky130_fd_sc_hd__o21ba_1
XFILLER_102_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5750_ _9056_/Q _8819_/X VGND VGND VPWR VPWR _5750_/Y sky130_fd_sc_hd__nor2_1
X_5681_ _5681_/A VGND VGND VPWR VPWR _5681_/Y sky130_fd_sc_hd__clkinv_2
X_4701_ _9688_/Q VGND VGND VPWR VPWR _4701_/Y sky130_fd_sc_hd__inv_2
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4632_ _9697_/Q VGND VGND VPWR VPWR _5214_/A sky130_fd_sc_hd__inv_2
X_7420_ _7474_/C _7466_/A _7474_/D VGND VGND VPWR VPWR _7421_/A sky130_fd_sc_hd__or3_1
XFILLER_175_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4563_ _4891_/A _6158_/A VGND VGND VPWR VPWR _4564_/B sky130_fd_sc_hd__or2_4
X_7351_ _6700_/Y _7124_/X _6701_/Y _7068_/B _7350_/X VGND VGND VPWR VPWR _7352_/D
+ sky130_fd_sc_hd__o221a_2
XFILLER_162_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7282_ _7282_/A _7392_/B VGND VGND VPWR VPWR _7282_/X sky130_fd_sc_hd__or2_1
X_6302_ _9156_/Q VGND VGND VPWR VPWR _6302_/Y sky130_fd_sc_hd__clkinv_2
X_4494_ _9785_/Q _4493_/A _8846_/X _4493_/Y VGND VGND VPWR VPWR _9785_/D sky130_fd_sc_hd__a22o_1
X_9021_ _9027_/CLK _9021_/D VGND VGND VPWR VPWR _9021_/Q sky130_fd_sc_hd__dfxtp_1
X_6233_ _6233_/A VGND VGND VPWR VPWR _6233_/Y sky130_fd_sc_hd__clkinv_4
X_6164_ _9404_/Q VGND VGND VPWR VPWR _6164_/Y sky130_fd_sc_hd__inv_2
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6095_ _6090_/Y _5458_/B _6091_/Y _5496_/B _6094_/X VGND VGND VPWR VPWR _6096_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_69_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5115_ _9637_/Q _5112_/A _8844_/X _5112_/Y VGND VGND VPWR VPWR _9637_/D sky130_fd_sc_hd__a22o_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5046_ _5046_/A VGND VGND VPWR VPWR _5047_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_27_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8805_ _8805_/A input1/X VGND VGND VPWR VPWR _8806_/A sky130_fd_sc_hd__and2_1
X_6997_ _6997_/A _8819_/X _6997_/C VGND VGND VPWR VPWR _6999_/A sky130_fd_sc_hd__or3_1
X_9785_ _9785_/CLK _9785_/D _9779_/SET_B VGND VGND VPWR VPWR _9785_/Q sky130_fd_sc_hd__dfrtp_1
X_8736_ _8164_/A _8550_/A _8029_/X _8411_/Y VGND VGND VPWR VPWR _8736_/X sky130_fd_sc_hd__o211a_1
X_5948_ _9114_/Q _5943_/A _5967_/B1 _5943_/Y VGND VGND VPWR VPWR _9114_/D sky130_fd_sc_hd__a22o_1
XFILLER_40_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5879_ _9154_/Q _5874_/A _8929_/A1 _5874_/Y VGND VGND VPWR VPWR _9154_/D sky130_fd_sc_hd__a22o_1
X_8667_ _8667_/A _8667_/B VGND VGND VPWR VPWR _8668_/B sky130_fd_sc_hd__or2_1
XFILLER_21_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8598_ _8695_/D _8659_/C _8727_/A _8657_/D VGND VGND VPWR VPWR _8601_/A sky130_fd_sc_hd__or4_2
X_7618_ _4722_/Y _7441_/X _4865_/Y _7443_/X _7617_/X VGND VGND VPWR VPWR _7625_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_181_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7549_ _6367_/Y _7465_/X _6427_/Y _7467_/X VGND VGND VPWR VPWR _7549_/X sky130_fd_sc_hd__o22a_1
XFILLER_5_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9219_ _9695_/CLK _9219_/D _9779_/SET_B VGND VGND VPWR VPWR _9219_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_122_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput201 wb_sel_i[3] VGND VGND VPWR VPWR _7734_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6920_ _9178_/Q VGND VGND VPWR VPWR _6920_/Y sky130_fd_sc_hd__clkinv_2
X_6851_ _6847_/Y _4868_/X _6848_/Y _5298_/B _6850_/X VGND VGND VPWR VPWR _6851_/X
+ sky130_fd_sc_hd__o221a_1
X_5802_ _9209_/Q _5799_/A _8844_/X _5799_/Y VGND VGND VPWR VPWR _9209_/D sky130_fd_sc_hd__a22o_1
X_9570_ _9613_/CLK _9570_/D _9646_/SET_B VGND VGND VPWR VPWR _9570_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_62_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8521_ _8521_/A _8521_/B VGND VGND VPWR VPWR _8521_/Y sky130_fd_sc_hd__nand2_1
XFILLER_22_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6782_ _6778_/Y _4893_/X _4949_/Y _6165_/A _6781_/X VGND VGND VPWR VPWR _6783_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_188_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5733_ _9248_/Q _7056_/B _7104_/A VGND VGND VPWR VPWR _7096_/B sky130_fd_sc_hd__or3_2
X_5664_ _9275_/Q _5662_/A _8845_/X _5662_/Y VGND VGND VPWR VPWR _9275_/D sky130_fd_sc_hd__a22o_1
XFILLER_148_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8452_ _8238_/A _7864_/X _8097_/B _8130_/B VGND VGND VPWR VPWR _8607_/C sky130_fd_sc_hd__o22ai_1
X_8383_ _8636_/A _8514_/A VGND VGND VPWR VPWR _8651_/B sky130_fd_sc_hd__or2_1
XFILLER_148_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5595_ _5595_/A VGND VGND VPWR VPWR _5596_/A sky130_fd_sc_hd__clkbuf_2
X_4615_ _4615_/A VGND VGND VPWR VPWR _4615_/Y sky130_fd_sc_hd__inv_2
X_7403_ _7413_/A _7406_/B VGND VGND VPWR VPWR _7476_/C sky130_fd_sc_hd__or2_4
X_4546_ _9068_/Q VGND VGND VPWR VPWR _8813_/A sky130_fd_sc_hd__inv_2
X_7334_ _6730_/Y _7082_/X _6705_/Y _7084_/X _7333_/X VGND VGND VPWR VPWR _7353_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_190_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7265_ _7265_/A _7265_/B _7265_/C VGND VGND VPWR VPWR _7265_/Y sky130_fd_sc_hd__nand3_4
X_4477_ _8839_/X _9789_/Q _4477_/S VGND VGND VPWR VPWR _4478_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9004_ _9597_/Q _8785_/A VGND VGND VPWR VPWR mgmt_gpio_out[27] sky130_fd_sc_hd__ebufn_8
X_7196_ _8783_/A _7126_/X _8781_/A _7128_/X VGND VGND VPWR VPWR _7196_/X sky130_fd_sc_hd__o22a_1
X_6216_ _6214_/Y _4577_/B _6215_/Y _5013_/B VGND VGND VPWR VPWR _6216_/X sky130_fd_sc_hd__o22a_1
X_6147_ _6974_/B _6147_/B VGND VGND VPWR VPWR _6148_/A sky130_fd_sc_hd__or2_1
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6078_ _9483_/Q VGND VGND VPWR VPWR _6078_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5029_ _9685_/Q _5026_/A _8841_/X _5026_/Y VGND VGND VPWR VPWR _9685_/D sky130_fd_sc_hd__a22o_1
XFILLER_72_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9768_ _9768_/CLK _9768_/D _4628_/A VGND VGND VPWR VPWR _9768_/Q sky130_fd_sc_hd__dfrtp_4
X_8719_ _8719_/A _8719_/B _8719_/C VGND VGND VPWR VPWR _8731_/C sky130_fd_sc_hd__or3_2
XFILLER_70_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9699_ _9709_/CLK _9699_/D _4995_/X VGND VGND VPWR VPWR _9699_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5380_ _9459_/Q _5376_/A _8930_/A1 _5376_/Y VGND VGND VPWR VPWR _9459_/D sky130_fd_sc_hd__a22o_1
XFILLER_132_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7050_ _7050_/A VGND VGND VPWR VPWR _7059_/A sky130_fd_sc_hd__buf_8
XFILLER_101_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6001_ _6001_/A VGND VGND VPWR VPWR _6001_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_140_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7952_ _7952_/A VGND VGND VPWR VPWR _8437_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_131_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6903_ _6903_/A VGND VGND VPWR VPWR _6903_/Y sky130_fd_sc_hd__inv_2
X_7883_ _8397_/A VGND VGND VPWR VPWR _7886_/B sky130_fd_sc_hd__inv_2
X_9622_ _9674_/CLK _9622_/D _9633_/SET_B VGND VGND VPWR VPWR _9622_/Q sky130_fd_sc_hd__dfrtp_1
X_6834_ _9733_/Q VGND VGND VPWR VPWR _6834_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6765_ _6760_/Y _5306_/B _6761_/Y _5240_/B _6764_/X VGND VGND VPWR VPWR _6783_/A
+ sky130_fd_sc_hd__o221a_1
X_9553_ _9639_/CLK _9553_/D _9757_/SET_B VGND VGND VPWR VPWR _9553_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8504_ _8501_/X _8504_/B _8504_/C VGND VGND VPWR VPWR _8504_/X sky130_fd_sc_hd__and3b_1
X_9484_ _9777_/CLK _9484_/D _9633_/SET_B VGND VGND VPWR VPWR _9484_/Q sky130_fd_sc_hd__dfrtp_1
X_5716_ _9249_/Q VGND VGND VPWR VPWR _5725_/B sky130_fd_sc_hd__inv_2
XFILLER_148_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8435_ _8636_/B _8435_/B VGND VGND VPWR VPWR _8436_/B sky130_fd_sc_hd__or2_1
XFILLER_136_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6696_ _6694_/Y _5267_/B _6695_/Y _5442_/B VGND VGND VPWR VPWR _6696_/X sky130_fd_sc_hd__o22a_1
XFILLER_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5647_ _5647_/A _5658_/A _5751_/C VGND VGND VPWR VPWR _5647_/X sky130_fd_sc_hd__or3_1
XFILLER_40_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5578_ _9324_/Q _5574_/A _8925_/A1 _5574_/Y VGND VGND VPWR VPWR _9324_/D sky130_fd_sc_hd__a22o_1
X_8366_ _8685_/B _8493_/B VGND VGND VPWR VPWR _8675_/A sky130_fd_sc_hd__or2_1
XFILLER_144_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8297_ _8651_/A _8606_/B VGND VGND VPWR VPWR _8673_/A sky130_fd_sc_hd__or2_1
X_7317_ _6826_/Y _7079_/B _6928_/Y _7059_/A VGND VGND VPWR VPWR _7317_/X sky130_fd_sc_hd__o22a_1
X_4529_ _9767_/Q _4526_/A _8844_/X _4526_/Y VGND VGND VPWR VPWR _9767_/D sky130_fd_sc_hd__a22o_1
XFILLER_116_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7248_ _6175_/Y _7048_/B _6215_/Y _7077_/A _7247_/X VGND VGND VPWR VPWR _7255_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_172_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7179_ _8757_/A _7077_/C _6491_/Y _7077_/D _7178_/X VGND VGND VPWR VPWR _7179_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_114 input86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_125 _7015_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_103 input86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_158 _8767_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_147 _6363_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_136 _7698_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_169 _7021_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput9 mask_rev_in[14] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__clkbuf_1
XFILLER_91_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4880_ _4877_/Y _5496_/B _4879_/Y _4517_/A VGND VGND VPWR VPWR _4880_/X sky130_fd_sc_hd__o22a_2
XFILLER_32_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6550_ _9539_/Q VGND VGND VPWR VPWR _6550_/Y sky130_fd_sc_hd__inv_2
XFILLER_192_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5501_ _9377_/Q _5498_/A _8844_/X _5498_/Y VGND VGND VPWR VPWR _9377_/D sky130_fd_sc_hd__a22o_1
X_6481_ _6479_/Y _5916_/B _6480_/Y _5564_/B VGND VGND VPWR VPWR _6481_/X sky130_fd_sc_hd__o22a_1
X_5432_ _5432_/A VGND VGND VPWR VPWR _5433_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_145_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8220_ _8566_/B _8214_/Y _8217_/Y _8110_/C _8219_/Y VGND VGND VPWR VPWR _8224_/C
+ sky130_fd_sc_hd__o32a_2
XFILLER_10_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput313 _7019_/X VGND VGND VPWR VPWR spimemio_flash_io0_di sky130_fd_sc_hd__buf_2
X_5363_ _9470_/Q _5357_/A _8841_/X _5357_/Y VGND VGND VPWR VPWR _9470_/D sky130_fd_sc_hd__a22o_1
XFILLER_145_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput335 _9028_/Q VGND VGND VPWR VPWR wb_dat_o[16] sky130_fd_sc_hd__buf_2
XFILLER_133_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8151_ _8552_/A _8640_/B VGND VGND VPWR VPWR _8674_/A sky130_fd_sc_hd__nor2_1
Xoutput324 _9769_/Q VGND VGND VPWR VPWR sram_ro_addr[7] sky130_fd_sc_hd__buf_2
Xoutput302 _9045_/Q VGND VGND VPWR VPWR pwr_ctrl_out[1] sky130_fd_sc_hd__buf_2
Xoutput346 _9038_/Q VGND VGND VPWR VPWR wb_dat_o[26] sky130_fd_sc_hd__buf_2
X_7102_ _4833_/Y _7079_/B _4726_/Y _7059_/A VGND VGND VPWR VPWR _7102_/X sky130_fd_sc_hd__o22a_1
Xoutput357 _9027_/Q VGND VGND VPWR VPWR wb_dat_o[7] sky130_fd_sc_hd__buf_2
XFILLER_126_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8082_ _8082_/A _8186_/A VGND VGND VPWR VPWR _8083_/C sky130_fd_sc_hd__and2_1
XFILLER_87_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5294_ _9518_/Q _5292_/A _5964_/B1 _5292_/Y VGND VGND VPWR VPWR _9518_/D sky130_fd_sc_hd__a22o_1
XFILLER_101_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7033_ _7033_/A VGND VGND VPWR VPWR _7040_/B sky130_fd_sc_hd__buf_8
XFILLER_142_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8984_ _9585_/Q _7699_/A VGND VGND VPWR VPWR mgmt_gpio_out[7] sky130_fd_sc_hd__ebufn_8
X_7935_ _8376_/A _7935_/B VGND VGND VPWR VPWR _7936_/B sky130_fd_sc_hd__or2_1
XFILLER_82_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7866_ _7866_/A VGND VGND VPWR VPWR _8319_/A sky130_fd_sc_hd__buf_2
X_9605_ _9617_/CLK _9605_/D _9295_/SET_B VGND VGND VPWR VPWR _9605_/Q sky130_fd_sc_hd__dfrtp_1
X_6817_ _6817_/A VGND VGND VPWR VPWR _6817_/Y sky130_fd_sc_hd__clkinv_2
X_7797_ _7797_/A VGND VGND VPWR VPWR _8188_/B sky130_fd_sc_hd__buf_2
XFILLER_23_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9536_ _9768_/CLK _9536_/D _4628_/A VGND VGND VPWR VPWR _9536_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_183_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6748_ _9288_/Q VGND VGND VPWR VPWR _6748_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9467_ _9514_/CLK _9467_/D _4628_/A VGND VGND VPWR VPWR _9467_/Q sky130_fd_sc_hd__dfrtp_1
X_6679_ _6679_/A VGND VGND VPWR VPWR _6679_/Y sky130_fd_sc_hd__inv_4
X_8418_ _8686_/A VGND VGND VPWR VPWR _8418_/Y sky130_fd_sc_hd__inv_2
X_9398_ _9758_/CLK _9398_/D _7011_/B VGND VGND VPWR VPWR _9398_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_164_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8349_ _8640_/A _8349_/B VGND VGND VPWR VPWR _8352_/B sky130_fd_sc_hd__or2_2
XFILLER_124_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5981_ _9090_/Q _5981_/B _9091_/Q VGND VGND VPWR VPWR _5981_/X sky130_fd_sc_hd__and3_1
X_4932_ _4928_/Y _5458_/B _4930_/Y _5328_/B VGND VGND VPWR VPWR _4932_/X sky130_fd_sc_hd__o22a_1
XFILLER_17_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7720_ _9087_/Q _7719_/B _7721_/A VGND VGND VPWR VPWR _7720_/X sky130_fd_sc_hd__o21a_1
XFILLER_178_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7651_ _6743_/Y _7430_/X _6725_/Y _7432_/X _7650_/X VGND VGND VPWR VPWR _7651_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA_14 _7500_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6602_ _6587_/Y _5480_/B _6590_/X _6596_/X _6601_/X VGND VGND VPWR VPWR _6628_/C
+ sky130_fd_sc_hd__o2111a_1
X_4863_ _4855_/Y _5317_/B _4857_/Y _4491_/B _4862_/X VGND VGND VPWR VPWR _4864_/D
+ sky130_fd_sc_hd__o221a_1
X_7582_ _6183_/Y _7441_/X _6195_/Y _7443_/X _7581_/X VGND VGND VPWR VPWR _7589_/A
+ sky130_fd_sc_hd__o221a_1
XANTENNA_25 _6165_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4794_ _4911_/A _4929_/A VGND VGND VPWR VPWR _5240_/B sky130_fd_sc_hd__or2_4
XANTENNA_47 _6291_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_36 _4935_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9321_ _9352_/CLK _9321_/D _9646_/SET_B VGND VGND VPWR VPWR _9321_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA_69 _7352_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_58 _6706_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6533_ _9657_/Q VGND VGND VPWR VPWR _6533_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9252_ _9279_/CLK _9252_/D _9633_/SET_B VGND VGND VPWR VPWR _9252_/Q sky130_fd_sc_hd__dfstp_1
X_6464_ _9658_/Q VGND VGND VPWR VPWR _6464_/Y sky130_fd_sc_hd__inv_2
X_8203_ _8203_/A VGND VGND VPWR VPWR _8476_/B sky130_fd_sc_hd__inv_2
XFILLER_146_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5415_ _9436_/Q _5414_/A _8843_/X _5414_/Y VGND VGND VPWR VPWR _9436_/D sky130_fd_sc_hd__a22o_1
XFILLER_161_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9183_ _9613_/CLK _9183_/D _9646_/SET_B VGND VGND VPWR VPWR _9183_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6395_ _6390_/Y _5355_/B _6391_/Y _5374_/B _6394_/X VGND VGND VPWR VPWR _6408_/B
+ sky130_fd_sc_hd__o221a_1
X_5346_ _5346_/A VGND VGND VPWR VPWR _5346_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8134_ _8137_/B _8640_/B VGND VGND VPWR VPWR _8642_/A sky130_fd_sc_hd__nor2_1
X_5277_ _9528_/Q _5269_/A _8839_/X _5269_/Y VGND VGND VPWR VPWR _9528_/D sky130_fd_sc_hd__a22o_1
X_8065_ _8065_/A _8703_/C VGND VGND VPWR VPWR _8067_/A sky130_fd_sc_hd__or2_1
XFILLER_114_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7016_ _7016_/A VGND VGND VPWR VPWR _7017_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_55_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8967_ _7749_/X _8967_/A1 _8975_/S VGND VGND VPWR VPWR _8967_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7918_ _8515_/B _8254_/B VGND VGND VPWR VPWR _8492_/A sky130_fd_sc_hd__or2_1
X_8898_ _9617_/Q _8846_/X _8930_/S VGND VGND VPWR VPWR _8898_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7849_ _8379_/D _8379_/B _8394_/C _8195_/A VGND VGND VPWR VPWR _7850_/A sky130_fd_sc_hd__or4_1
XFILLER_178_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9519_ _9771_/CLK _9519_/D _4628_/A VGND VGND VPWR VPWR _9519_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_109_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_1_0_mgmt_gpio_in[4] clkbuf_2_1_0_mgmt_gpio_in[4]/A VGND VGND VPWR VPWR _9709_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput12 mask_rev_in[17] VGND VGND VPWR VPWR _6794_/A sky130_fd_sc_hd__clkbuf_1
Xinput45 mgmt_gpio_in[18] VGND VGND VPWR VPWR input45/X sky130_fd_sc_hd__buf_2
Xinput34 mask_rev_in[8] VGND VGND VPWR VPWR input34/X sky130_fd_sc_hd__buf_2
Xinput23 mask_rev_in[27] VGND VGND VPWR VPWR _6624_/A sky130_fd_sc_hd__clkbuf_1
Xinput56 mgmt_gpio_in[28] VGND VGND VPWR VPWR input56/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput89 spimemio_flash_io2_do VGND VGND VPWR VPWR input89/X sky130_fd_sc_hd__clkbuf_4
XFILLER_143_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput78 spi_csb VGND VGND VPWR VPWR input78/X sky130_fd_sc_hd__buf_6
XFILLER_6_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput67 mgmt_gpio_in[3] VGND VGND VPWR VPWR _4629_/C sky130_fd_sc_hd__buf_12
XFILLER_170_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6180_ _6178_/Y _5679_/B _6179_/Y _5660_/B VGND VGND VPWR VPWR _6187_/B sky130_fd_sc_hd__o22a_1
X_5200_ _9579_/Q _5193_/Y _8903_/X _5193_/A VGND VGND VPWR VPWR _9579_/D sky130_fd_sc_hd__o22a_1
XFILLER_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5131_ _9048_/Q _4951_/B _9708_/Q _9626_/Q _4951_/Y VGND VGND VPWR VPWR _9626_/D
+ sky130_fd_sc_hd__a32o_1
X_5062_ _5062_/A _5062_/B _5062_/C _5062_/D VGND VGND VPWR VPWR _5063_/A sky130_fd_sc_hd__or4_1
X_8821_ _9057_/Q _9078_/Q _9787_/Q VGND VGND VPWR VPWR _8821_/X sky130_fd_sc_hd__mux2_1
X_8752_ _8752_/A VGND VGND VPWR VPWR _8752_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5964_ _9104_/Q _5962_/A _5964_/B1 _5962_/Y VGND VGND VPWR VPWR _9104_/D sky130_fd_sc_hd__a22o_1
X_7703_ _7703_/A VGND VGND VPWR VPWR _7704_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_178_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8683_ _8683_/A _8683_/B VGND VGND VPWR VPWR _8683_/X sky130_fd_sc_hd__or2_1
X_4915_ _6086_/B _4931_/B VGND VGND VPWR VPWR _5420_/B sky130_fd_sc_hd__or2_4
X_5895_ _8959_/X VGND VGND VPWR VPWR _5895_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4846_ _9528_/Q VGND VGND VPWR VPWR _4846_/Y sky130_fd_sc_hd__inv_2
X_7634_ _6929_/Y _7425_/X _7631_/X _7633_/X VGND VGND VPWR VPWR _7644_/C sky130_fd_sc_hd__o211a_1
XFILLER_32_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7565_ _6277_/Y _7455_/X _6314_/Y _7457_/X VGND VGND VPWR VPWR _7565_/X sky130_fd_sc_hd__o22a_1
X_9304_ _9440_/CLK _9304_/D _9685_/SET_B VGND VGND VPWR VPWR _9304_/Q sky130_fd_sc_hd__dfrtp_1
X_4777_ _4773_/Y _5045_/B _4775_/Y _5916_/B VGND VGND VPWR VPWR _4777_/X sky130_fd_sc_hd__o22a_2
X_6516_ _9104_/Q VGND VGND VPWR VPWR _6516_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_134_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7496_ _6920_/Y _7461_/X _6832_/Y _7463_/X _7495_/X VGND VGND VPWR VPWR _7499_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9235_ _9508_/CLK _9235_/D _9528_/SET_B VGND VGND VPWR VPWR _9235_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_161_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6447_ _6444_/Y _4832_/X _6445_/Y _5100_/B _6446_/Y VGND VGND VPWR VPWR _6447_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_164_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6378_ _9285_/Q VGND VGND VPWR VPWR _7392_/A sky130_fd_sc_hd__clkinv_2
X_9166_ _9203_/CLK _9166_/D _9633_/SET_B VGND VGND VPWR VPWR _9166_/Q sky130_fd_sc_hd__dfrtp_1
X_8117_ _8117_/A _8117_/B VGND VGND VPWR VPWR _8393_/A sky130_fd_sc_hd__nand2_2
XFILLER_102_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5329_ _5329_/A VGND VGND VPWR VPWR _5330_/A sky130_fd_sc_hd__clkbuf_2
X_9097_ _9501_/CLK _9097_/D _9647_/SET_B VGND VGND VPWR VPWR _9097_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_102_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8048_ _8554_/A _8389_/A _8047_/X VGND VGND VPWR VPWR _8048_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_57_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5680_ _5680_/A VGND VGND VPWR VPWR _5681_/A sky130_fd_sc_hd__clkbuf_4
X_4700_ _4931_/A _4843_/B VGND VGND VPWR VPWR _5897_/B sky130_fd_sc_hd__or2_4
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4631_ _6050_/A VGND VGND VPWR VPWR _4994_/A sky130_fd_sc_hd__buf_12
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4562_ _4562_/A VGND VGND VPWR VPWR _9756_/D sky130_fd_sc_hd__clkbuf_1
X_7350_ _6652_/Y _7126_/X _6762_/Y _7128_/X VGND VGND VPWR VPWR _7350_/X sky130_fd_sc_hd__o22a_1
X_7281_ _6127_/Y _7059_/D _6091_/Y _7116_/X _7280_/X VGND VGND VPWR VPWR _7286_/B
+ sky130_fd_sc_hd__o221a_1
X_6301_ _9223_/Q VGND VGND VPWR VPWR _6301_/Y sky130_fd_sc_hd__inv_2
X_4493_ _4493_/A VGND VGND VPWR VPWR _4493_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9020_ _9027_/CLK _9020_/D VGND VGND VPWR VPWR _9020_/Q sky130_fd_sc_hd__dfxtp_1
X_6232_ _9673_/Q VGND VGND VPWR VPWR _6232_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_170_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6163_ _9318_/Q VGND VGND VPWR VPWR _6163_/Y sky130_fd_sc_hd__inv_2
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6094_ _6092_/Y _4577_/B _6093_/Y _4907_/X VGND VGND VPWR VPWR _6094_/X sky130_fd_sc_hd__o22a_2
X_5114_ _9638_/Q _5112_/A _8845_/X _5112_/Y VGND VGND VPWR VPWR _9638_/D sky130_fd_sc_hd__a22o_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5045_ _5960_/A _5045_/B VGND VGND VPWR VPWR _5046_/A sky130_fd_sc_hd__or2_1
XFILLER_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8804_ _8804_/A VGND VGND VPWR VPWR _8804_/X sky130_fd_sc_hd__clkbuf_1
X_9784_ _9785_/CLK _9784_/D _9779_/SET_B VGND VGND VPWR VPWR _9784_/Q sky130_fd_sc_hd__dfrtp_1
X_6996_ _7075_/A _7094_/B VGND VGND VPWR VPWR _6996_/Y sky130_fd_sc_hd__nor2_2
X_8735_ _8735_/A _8735_/B _8735_/C _8735_/D VGND VGND VPWR VPWR _8735_/X sky130_fd_sc_hd__or4_1
X_5947_ _9115_/Q _5943_/A _8930_/A1 _5943_/Y VGND VGND VPWR VPWR _9115_/D sky130_fd_sc_hd__a22o_1
XFILLER_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8666_ _8666_/A _8666_/B _8666_/C _8666_/D VGND VGND VPWR VPWR _8735_/D sky130_fd_sc_hd__or4_2
XFILLER_33_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5878_ _9155_/Q _5874_/A _8925_/A1 _5874_/Y VGND VGND VPWR VPWR _9155_/D sky130_fd_sc_hd__a22o_1
X_7617_ _4848_/Y _7445_/X _4918_/Y _7447_/X VGND VGND VPWR VPWR _7617_/X sky130_fd_sc_hd__o22a_1
XFILLER_193_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4829_ _4821_/Y _4822_/X _4823_/Y _5100_/B _4828_/X VGND VGND VPWR VPWR _4830_/D
+ sky130_fd_sc_hd__o221a_1
X_8597_ _8597_/A _8597_/B _8597_/C _8597_/D VGND VGND VPWR VPWR _8657_/D sky130_fd_sc_hd__or4_4
XFILLER_193_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7548_ _6353_/Y _7451_/X _6415_/Y _7453_/X _7547_/X VGND VGND VPWR VPWR _7553_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_181_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7479_ _4668_/Y _7471_/X _7121_/A _7473_/X _7478_/X VGND VGND VPWR VPWR _7480_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_4_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9218_ _9379_/CLK _9218_/D _9646_/SET_B VGND VGND VPWR VPWR _9218_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_134_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput202 wb_stb_i VGND VGND VPWR VPWR input202/X sky130_fd_sc_hd__clkbuf_4
XFILLER_108_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9149_ _9280_/CLK _9149_/D _9757_/SET_B VGND VGND VPWR VPWR _9149_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_102_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1 hold1/A VGND VGND VPWR VPWR hold1/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_82_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6850_ _9787_/Q _6251_/Y _6849_/Y _6086_/X VGND VGND VPWR VPWR _6850_/X sky130_fd_sc_hd__o2bb2a_2
XFILLER_35_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5801_ _9210_/Q _5799_/A _8845_/X _5799_/Y VGND VGND VPWR VPWR _9210_/D sky130_fd_sc_hd__a22o_1
X_6781_ _6779_/Y _5290_/B _6780_/Y _5328_/B VGND VGND VPWR VPWR _6781_/X sky130_fd_sc_hd__o22a_1
X_8520_ _8472_/Y _8517_/Y _8518_/X _8444_/B VGND VGND VPWR VPWR _8612_/B sky130_fd_sc_hd__a31o_1
X_5732_ _9249_/Q _5731_/Y _5724_/Y VGND VGND VPWR VPWR _9249_/D sky130_fd_sc_hd__o21ba_1
Xclkbuf_1_1_1_mgmt_gpio_in[4] clkbuf_1_1_1_mgmt_gpio_in[4]/A VGND VGND VPWR VPWR clkbuf_2_3_0_mgmt_gpio_in[4]/A
+ sky130_fd_sc_hd__clkbuf_2
X_5663_ _9276_/Q _5662_/A _8846_/X _5662_/Y VGND VGND VPWR VPWR _9276_/D sky130_fd_sc_hd__a22o_1
X_8451_ _8451_/A _8683_/A VGND VGND VPWR VPWR _8453_/C sky130_fd_sc_hd__or2_1
X_8382_ _8705_/A _8382_/B VGND VGND VPWR VPWR _8384_/A sky130_fd_sc_hd__or2_1
XFILLER_135_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5594_ _5671_/A _5594_/B VGND VGND VPWR VPWR _5595_/A sky130_fd_sc_hd__or2_1
X_4614_ _4614_/A VGND VGND VPWR VPWR _4615_/A sky130_fd_sc_hd__clkbuf_2
X_7402_ _9254_/Q VGND VGND VPWR VPWR _7413_/A sky130_fd_sc_hd__inv_2
X_4545_ _9067_/Q VGND VGND VPWR VPWR _8812_/A sky130_fd_sc_hd__inv_2
XFILLER_163_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7333_ _6645_/Y _7077_/C _6756_/Y _7077_/D _7332_/X VGND VGND VPWR VPWR _7333_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_190_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9003_ _9596_/Q _8783_/A VGND VGND VPWR VPWR mgmt_gpio_out[26] sky130_fd_sc_hd__ebufn_8
X_4476_ _4787_/A _4891_/A _5259_/A VGND VGND VPWR VPWR _4477_/S sky130_fd_sc_hd__or3_1
XFILLER_116_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7264_ _7264_/A _7264_/B _7264_/C _7264_/D VGND VGND VPWR VPWR _7265_/C sky130_fd_sc_hd__and4_1
XFILLER_131_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7195_ _8793_/A _5728_/X _7705_/A _7040_/A _7194_/X VGND VGND VPWR VPWR _7198_/C
+ sky130_fd_sc_hd__o221a_1
X_6215_ _9694_/Q VGND VGND VPWR VPWR _6215_/Y sky130_fd_sc_hd__inv_2
X_6146_ _6146_/A VGND VGND VPWR VPWR _6974_/B sky130_fd_sc_hd__inv_2
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6077_ _6072_/Y _5393_/B _6073_/Y _5317_/B _6076_/X VGND VGND VPWR VPWR _6096_/A
+ sky130_fd_sc_hd__o221a_1
X_5028_ _9686_/Q _5026_/A _8842_/X _5026_/Y VGND VGND VPWR VPWR _9686_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6979_ _6326_/Y _6976_/A _9017_/Q _6976_/Y VGND VGND VPWR VPWR _9017_/D sky130_fd_sc_hd__o22a_1
X_9767_ _9769_/CLK _9767_/D _9757_/SET_B VGND VGND VPWR VPWR _9767_/Q sky130_fd_sc_hd__dfrtp_2
X_8718_ _8347_/X _8717_/X _8223_/B _8312_/D VGND VGND VPWR VPWR _8719_/B sky130_fd_sc_hd__o211ai_1
XFILLER_110_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9698_ _9709_/CLK _9698_/D _5000_/X VGND VGND VPWR VPWR _9698_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_166_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8649_ _8722_/A _8681_/B _8720_/B VGND VGND VPWR VPWR _8649_/Y sky130_fd_sc_hd__nor3_1
XFILLER_186_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6000_ _6040_/A VGND VGND VPWR VPWR _6001_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7951_ _8525_/A _8538_/B _8538_/C _8084_/A VGND VGND VPWR VPWR _7952_/A sky130_fd_sc_hd__or4_1
X_6902_ _9684_/Q VGND VGND VPWR VPWR _6902_/Y sky130_fd_sc_hd__inv_4
X_7882_ _8394_/D _8097_/B VGND VGND VPWR VPWR _8397_/A sky130_fd_sc_hd__or2_4
XFILLER_23_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6833_ _9642_/Q VGND VGND VPWR VPWR _6833_/Y sky130_fd_sc_hd__clkinv_2
X_9621_ _9674_/CLK _9621_/D _9633_/SET_B VGND VGND VPWR VPWR _9621_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6764_ _6762_/Y _5251_/B _6763_/Y _5393_/B VGND VGND VPWR VPWR _6764_/X sky130_fd_sc_hd__o22a_1
X_9552_ _9639_/CLK _9552_/D _9633_/SET_B VGND VGND VPWR VPWR _9552_/Q sky130_fd_sc_hd__dfrtp_1
X_9483_ _9483_/CLK _9483_/D _9685_/SET_B VGND VGND VPWR VPWR _9483_/Q sky130_fd_sc_hd__dfrtp_1
X_6695_ _9413_/Q VGND VGND VPWR VPWR _6695_/Y sky130_fd_sc_hd__clkinv_2
X_8503_ _8341_/A _8239_/B _8238_/A _8498_/B _7910_/X VGND VGND VPWR VPWR _8504_/C
+ sky130_fd_sc_hd__o221a_1
X_5715_ _9250_/Q VGND VGND VPWR VPWR _6994_/A sky130_fd_sc_hd__inv_2
XFILLER_50_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8434_ _8434_/A _8636_/C VGND VGND VPWR VPWR _8435_/B sky130_fd_sc_hd__nor2_1
X_5646_ _9278_/Q VGND VGND VPWR VPWR _5751_/C sky130_fd_sc_hd__inv_2
XFILLER_163_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5577_ _9325_/Q _5574_/A _8844_/X _5574_/Y VGND VGND VPWR VPWR _9325_/D sky130_fd_sc_hd__a22o_1
X_8365_ _8551_/A _8378_/B _8250_/A VGND VGND VPWR VPWR _8577_/C sky130_fd_sc_hd__o21ai_1
XFILLER_163_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8296_ _8296_/A _8296_/B VGND VGND VPWR VPWR _8296_/Y sky130_fd_sc_hd__nand2_1
XFILLER_104_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7316_ _6866_/Y _7095_/X _6935_/Y _7068_/D _7315_/X VGND VGND VPWR VPWR _7321_/B
+ sky130_fd_sc_hd__o221a_1
X_4528_ _9768_/Q _4526_/A _8845_/X _4526_/Y VGND VGND VPWR VPWR _9768_/D sky130_fd_sc_hd__a22o_1
X_7247_ _6232_/Y _7040_/C _6224_/Y _7059_/C VGND VGND VPWR VPWR _7247_/X sky130_fd_sc_hd__o22a_1
X_4459_ _4459_/A VGND VGND VPWR VPWR _6111_/A sky130_fd_sc_hd__clkbuf_8
X_7178_ _8773_/A _7086_/X _8771_/A _7088_/X VGND VGND VPWR VPWR _7178_/X sky130_fd_sc_hd__o22a_1
XFILLER_58_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6129_ _9674_/Q VGND VGND VPWR VPWR _6129_/Y sky130_fd_sc_hd__clkinv_2
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_104 input86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_115 _8816_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_126 input91/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_137 _5960_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_148 _6584_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_159 _8791_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5500_ _9378_/Q _5498_/A _8845_/X _5498_/Y VGND VGND VPWR VPWR _9378_/D sky130_fd_sc_hd__a22o_1
XFILLER_185_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6480_ _9331_/Q VGND VGND VPWR VPWR _6480_/Y sky130_fd_sc_hd__inv_2
X_5431_ _5545_/A _5431_/B VGND VGND VPWR VPWR _5432_/A sky130_fd_sc_hd__or2_1
XFILLER_145_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput314 _7021_/X VGND VGND VPWR VPWR spimemio_flash_io1_di sky130_fd_sc_hd__buf_2
X_5362_ _9471_/Q _5357_/A _8842_/X _5357_/Y VGND VGND VPWR VPWR _9471_/D sky130_fd_sc_hd__a22o_1
XFILLER_114_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8150_ _8150_/A _8685_/B VGND VGND VPWR VPWR _8152_/A sky130_fd_sc_hd__or2_1
Xoutput325 _9760_/Q VGND VGND VPWR VPWR sram_ro_clk sky130_fd_sc_hd__buf_2
Xoutput303 _9046_/Q VGND VGND VPWR VPWR pwr_ctrl_out[2] sky130_fd_sc_hd__buf_2
Xoutput347 _9039_/Q VGND VGND VPWR VPWR wb_dat_o[27] sky130_fd_sc_hd__buf_2
X_8081_ _8188_/B _8640_/B VGND VGND VPWR VPWR _8186_/A sky130_fd_sc_hd__or2_1
Xoutput336 _9029_/Q VGND VGND VPWR VPWR wb_dat_o[17] sky130_fd_sc_hd__buf_2
Xoutput358 _9012_/Q VGND VGND VPWR VPWR wb_dat_o[8] sky130_fd_sc_hd__buf_2
X_7101_ _4897_/Y _7095_/X _4779_/Y _7068_/D _7100_/X VGND VGND VPWR VPWR _7108_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_99_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7032_ _7073_/C _7109_/B VGND VGND VPWR VPWR _7033_/A sky130_fd_sc_hd__or2_1
X_5293_ _9519_/Q _5292_/A _5963_/B1 _5292_/Y VGND VGND VPWR VPWR _9519_/D sky130_fd_sc_hd__a22o_1
XFILLER_59_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8983_ _8983_/A _7701_/A VGND VGND VPWR VPWR mgmt_gpio_out[6] sky130_fd_sc_hd__ebufn_8
X_7934_ _8282_/C _7836_/C _7831_/Y _7933_/X VGND VGND VPWR VPWR _7935_/B sky130_fd_sc_hd__a31o_1
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7865_ _7959_/A _8528_/A _8525_/A _8189_/A VGND VGND VPWR VPWR _7866_/A sky130_fd_sc_hd__or4_4
XFILLER_63_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9604_ _9617_/CLK _9604_/D _9295_/SET_B VGND VGND VPWR VPWR _9604_/Q sky130_fd_sc_hd__dfrtp_1
X_7796_ _8084_/A _8085_/A VGND VGND VPWR VPWR _7797_/A sky130_fd_sc_hd__or2_1
X_6816_ _6811_/Y _4613_/B _6812_/Y _4504_/B _6815_/X VGND VGND VPWR VPWR _6829_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9535_ _9535_/CLK _9535_/D _9528_/SET_B VGND VGND VPWR VPWR _9535_/Q sky130_fd_sc_hd__dfrtp_1
X_6747_ _6742_/Y _5110_/B _6743_/Y _5916_/B _6746_/X VGND VGND VPWR VPWR _6759_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_149_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6678_ _6673_/Y _5968_/B _6674_/Y _5864_/B _6677_/X VGND VGND VPWR VPWR _6690_/B
+ sky130_fd_sc_hd__o221a_1
X_9466_ _9514_/CLK _9466_/D _4628_/A VGND VGND VPWR VPWR _9466_/Q sky130_fd_sc_hd__dfrtp_1
X_9397_ _9509_/CLK _9397_/D _9528_/SET_B VGND VGND VPWR VPWR _9397_/Q sky130_fd_sc_hd__dfrtp_1
X_5629_ _9288_/Q _5623_/A _8955_/A1 _5623_/Y VGND VGND VPWR VPWR _9288_/D sky130_fd_sc_hd__a22o_1
XFILLER_109_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8417_ _8667_/B _8577_/A VGND VGND VPWR VPWR _8686_/A sky130_fd_sc_hd__or2_1
XFILLER_191_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8348_ _8378_/B _8347_/X _8216_/X VGND VGND VPWR VPWR _8349_/B sky130_fd_sc_hd__o21a_1
XFILLER_104_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8279_ _8279_/A _8378_/B _8279_/C VGND VGND VPWR VPWR _8280_/C sky130_fd_sc_hd__or3_1
XFILLER_104_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5980_ _5980_/A VGND VGND VPWR VPWR _5980_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_17_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4931_ _4931_/A _4931_/B VGND VGND VPWR VPWR _5328_/B sky130_fd_sc_hd__or2_4
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4862_ _4858_/Y _5374_/B _4860_/Y _4861_/X VGND VGND VPWR VPWR _4862_/X sky130_fd_sc_hd__o22a_1
X_7650_ _6779_/Y _7434_/X _6780_/Y _7436_/X VGND VGND VPWR VPWR _7650_/X sky130_fd_sc_hd__o22a_1
XFILLER_177_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6601_ _6597_/Y _5232_/B _8785_/A _5240_/B _6600_/X VGND VGND VPWR VPWR _6601_/X
+ sky130_fd_sc_hd__o221a_1
X_9320_ _9613_/CLK _9320_/D _9646_/SET_B VGND VGND VPWR VPWR _9320_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA_26 _4777_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_48 _6294_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7581_ _6225_/Y _7445_/X _6164_/Y _7447_/X VGND VGND VPWR VPWR _7581_/X sky130_fd_sc_hd__o22a_1
XANTENNA_37 _6096_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4793_ _9546_/Q VGND VGND VPWR VPWR _4793_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_20_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_15 _7518_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6532_ _9154_/Q VGND VGND VPWR VPWR _7699_/A sky130_fd_sc_hd__clkinv_4
XANTENNA_59 _6787_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9251_ _9279_/CLK _9251_/D _9633_/SET_B VGND VGND VPWR VPWR _9251_/Q sky130_fd_sc_hd__dfrtp_4
X_6463_ _9671_/Q VGND VGND VPWR VPWR _6463_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_173_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8202_ _8202_/A _8213_/A VGND VGND VPWR VPWR _8721_/A sky130_fd_sc_hd__nor2_4
XFILLER_161_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9182_ _9652_/CLK _9182_/D _9646_/SET_B VGND VGND VPWR VPWR _9182_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5414_ _5414_/A VGND VGND VPWR VPWR _5414_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6394_ _6392_/Y _6081_/B _6393_/Y _5602_/B VGND VGND VPWR VPWR _6394_/X sky130_fd_sc_hd__o22a_1
X_8133_ _8133_/A VGND VGND VPWR VPWR _8358_/A sky130_fd_sc_hd__inv_2
X_5345_ _5345_/A VGND VGND VPWR VPWR _5346_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_87_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5276_ _9529_/Q _5269_/A _8930_/A1 _5269_/Y VGND VGND VPWR VPWR _9529_/D sky130_fd_sc_hd__a22o_1
X_8064_ _8518_/A _8064_/B _8064_/C VGND VGND VPWR VPWR _8703_/C sky130_fd_sc_hd__and3_1
XFILLER_114_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7015_ _9586_/Q _7015_/B VGND VGND VPWR VPWR _7016_/A sky130_fd_sc_hd__or2_1
XFILLER_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8966_ _7747_/X _8966_/A1 _8975_/S VGND VGND VPWR VPWR _8966_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7917_ _8734_/A _7917_/B _8317_/A _8597_/A VGND VGND VPWR VPWR _7917_/Y sky130_fd_sc_hd__nor4_1
XFILLER_169_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8897_ _8896_/X _9149_/Q _9054_/Q VGND VGND VPWR VPWR _8897_/X sky130_fd_sc_hd__mux2_1
X_7848_ _7848_/A _8077_/A VGND VGND VPWR VPWR _7929_/A sky130_fd_sc_hd__or2_1
XFILLER_11_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7779_ _7832_/A _7837_/B _5934_/X VGND VGND VPWR VPWR _8218_/B sky130_fd_sc_hd__o21ai_2
XFILLER_178_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9518_ _9545_/CLK _9518_/D _4628_/A VGND VGND VPWR VPWR _9518_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_149_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9449_ _9785_/CLK _9449_/D _9779_/SET_B VGND VGND VPWR VPWR _9449_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_191_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput13 mask_rev_in[18] VGND VGND VPWR VPWR _6766_/A sky130_fd_sc_hd__clkbuf_1
Xinput46 mgmt_gpio_in[19] VGND VGND VPWR VPWR _6521_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_128_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput35 mask_rev_in[9] VGND VGND VPWR VPWR _6849_/A sky130_fd_sc_hd__clkbuf_1
Xinput24 mask_rev_in[28] VGND VGND VPWR VPWR _6411_/A sky130_fd_sc_hd__clkbuf_1
Xinput57 mgmt_gpio_in[29] VGND VGND VPWR VPWR input57/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput79 spi_enabled VGND VGND VPWR VPWR _8833_/S sky130_fd_sc_hd__buf_6
Xinput68 mgmt_gpio_in[5] VGND VGND VPWR VPWR _8801_/A sky130_fd_sc_hd__buf_4
XFILLER_170_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5130_ _5130_/A VGND VGND VPWR VPWR _5130_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5061_ _8812_/A _5058_/X _8811_/A _5060_/X VGND VGND VPWR VPWR _5062_/C sky130_fd_sc_hd__o22ai_1
XFILLER_151_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8820_ _9217_/Q _9069_/Q _9787_/Q VGND VGND VPWR VPWR _8820_/X sky130_fd_sc_hd__mux2_1
X_8751_ _8751_/A VGND VGND VPWR VPWR _8752_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_92_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5963_ _9105_/Q _5962_/A _5963_/B1 _5962_/Y VGND VGND VPWR VPWR _9105_/D sky130_fd_sc_hd__a22o_1
X_4914_ _9424_/Q VGND VGND VPWR VPWR _4914_/Y sky130_fd_sc_hd__clkinv_2
X_7702_ _7702_/A VGND VGND VPWR VPWR _7702_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_opt_4_0_csclk clkbuf_2_1_0_csclk/X VGND VGND VPWR VPWR clkbuf_opt_4_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_16
X_8682_ _8720_/B _8722_/A _8722_/B _8723_/A VGND VGND VPWR VPWR _8682_/X sky130_fd_sc_hd__or4_4
X_5894_ _5849_/A _8875_/X _8924_/X _9139_/Q VGND VGND VPWR VPWR _9139_/D sky130_fd_sc_hd__o22a_1
XFILLER_178_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7633_ _6922_/Y _7430_/X _6805_/Y _7432_/X _7632_/X VGND VGND VPWR VPWR _7633_/X
+ sky130_fd_sc_hd__o221a_1
X_4845_ _4840_/Y _4841_/X _4842_/Y _5968_/B _4844_/X VGND VGND VPWR VPWR _4864_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_193_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7564_ _6308_/Y _7441_/X _6256_/Y _7443_/X _7563_/X VGND VGND VPWR VPWR _7571_/A
+ sky130_fd_sc_hd__o221a_1
X_4776_ _4925_/A _4843_/B VGND VGND VPWR VPWR _5916_/B sky130_fd_sc_hd__or2_4
X_6515_ _9272_/Q VGND VGND VPWR VPWR _8759_/A sky130_fd_sc_hd__inv_4
X_9303_ _9440_/CLK _9303_/D _9685_/SET_B VGND VGND VPWR VPWR _9303_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_173_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7495_ _6879_/Y _7465_/X _6825_/Y _7467_/X VGND VGND VPWR VPWR _7495_/X sky130_fd_sc_hd__o22a_1
XFILLER_106_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6446_ input56/X _6322_/Y _8817_/A _4680_/Y VGND VGND VPWR VPWR _6446_/Y sky130_fd_sc_hd__a22oi_4
X_9234_ _9371_/CLK _9234_/D _9295_/SET_B VGND VGND VPWR VPWR _9234_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_134_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6377_ _9273_/Q VGND VGND VPWR VPWR _6377_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9165_ _9203_/CLK _9165_/D _9633_/SET_B VGND VGND VPWR VPWR _9165_/Q sky130_fd_sc_hd__dfrtp_1
X_9096_ _9501_/CLK _9096_/D _9647_/SET_B VGND VGND VPWR VPWR _9096_/Q sky130_fd_sc_hd__dfrtp_4
X_8116_ _8116_/A _8116_/B VGND VGND VPWR VPWR _8117_/B sky130_fd_sc_hd__or2_2
XFILLER_0_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5328_ _5671_/A _5328_/B VGND VGND VPWR VPWR _5329_/A sky130_fd_sc_hd__or2_1
XFILLER_114_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8047_ _8047_/A _8467_/A VGND VGND VPWR VPWR _8047_/X sky130_fd_sc_hd__and2_1
XFILLER_87_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5259_ _5259_/A _5259_/B VGND VGND VPWR VPWR _5260_/A sky130_fd_sc_hd__or2_1
XFILLER_68_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8949_ _9713_/Q _6629_/Y _8957_/S VGND VGND VPWR VPWR _8949_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4630_ _6052_/B _7022_/B VGND VGND VPWR VPWR _6050_/A sky130_fd_sc_hd__nor2_8
XFILLER_175_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6300_ _6296_/Y _5621_/B _6297_/Y _5013_/B _6299_/X VGND VGND VPWR VPWR _6307_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_8_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4561_ _5967_/B1 _9756_/Q _4561_/S VGND VGND VPWR VPWR _4562_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7280_ _6109_/Y _7118_/X _6068_/Y _7048_/C VGND VGND VPWR VPWR _7280_/X sky130_fd_sc_hd__o22a_1
X_4492_ _4492_/A VGND VGND VPWR VPWR _4493_/A sky130_fd_sc_hd__buf_2
XFILLER_170_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6231_ _9638_/Q VGND VGND VPWR VPWR _6231_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6162_ _6157_/Y _5089_/B _6158_/X _6161_/X VGND VGND VPWR VPWR _6174_/B sky130_fd_sc_hd__o211a_1
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5113_ _9639_/Q _5112_/A _8846_/X _5112_/Y VGND VGND VPWR VPWR _9639_/D sky130_fd_sc_hd__a22o_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6093_ _6093_/A VGND VGND VPWR VPWR _6093_/Y sky130_fd_sc_hd__inv_2
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5044_ _8969_/X _4551_/B _9675_/Q _5062_/D VGND VGND VPWR VPWR _9675_/D sky130_fd_sc_hd__a22o_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8803_ _8803_/A _8833_/S VGND VGND VPWR VPWR _8804_/A sky130_fd_sc_hd__and2_1
XFILLER_38_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9783_ _9785_/CLK _9783_/D _9779_/SET_B VGND VGND VPWR VPWR _9783_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_53_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6995_ _9248_/Q _7056_/B _7125_/A VGND VGND VPWR VPWR _7094_/B sky130_fd_sc_hd__or3_1
X_8734_ _8734_/A _8734_/B _8734_/C _8734_/D VGND VGND VPWR VPWR _8735_/B sky130_fd_sc_hd__or4_1
XFILLER_80_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5946_ _9116_/Q _5943_/A _5965_/B1 _5943_/Y VGND VGND VPWR VPWR _9116_/D sky130_fd_sc_hd__a22o_1
XFILLER_139_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5877_ _9156_/Q _5874_/A _8844_/X _5874_/Y VGND VGND VPWR VPWR _9156_/D sky130_fd_sc_hd__a22o_1
X_8665_ _8665_/A _8665_/B _7877_/X VGND VGND VPWR VPWR _8666_/B sky130_fd_sc_hd__or3b_1
XFILLER_193_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7616_ _4765_/Y _7425_/X _7613_/X _7615_/X VGND VGND VPWR VPWR _7626_/C sky130_fd_sc_hd__o211a_1
X_4828_ _8807_/A _5227_/B _4827_/Y _6251_/A VGND VGND VPWR VPWR _4828_/X sky130_fd_sc_hd__o22a_1
XFILLER_178_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8596_ _8077_/A _8239_/B _8236_/A _8304_/Y _8504_/B VGND VGND VPWR VPWR _8727_/A
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_193_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4759_ _9294_/Q VGND VGND VPWR VPWR _7121_/A sky130_fd_sc_hd__clkinv_4
XFILLER_153_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7547_ _6398_/Y _7455_/X _6439_/Y _7457_/X VGND VGND VPWR VPWR _7547_/X sky130_fd_sc_hd__o22a_1
XFILLER_175_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7478_ _4814_/Y _7475_/X _4726_/Y _7477_/X VGND VGND VPWR VPWR _7478_/X sky130_fd_sc_hd__o22a_1
XFILLER_107_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9217_ _9280_/CLK _9217_/D _9757_/SET_B VGND VGND VPWR VPWR _9217_/Q sky130_fd_sc_hd__dfrtp_1
X_6429_ _9777_/Q VGND VGND VPWR VPWR _6429_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_134_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9148_ _9280_/CLK _9148_/D _9757_/SET_B VGND VGND VPWR VPWR _9148_/Q sky130_fd_sc_hd__dfrtp_1
Xinput203 wb_we_i VGND VGND VPWR VPWR _7734_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_88_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9079_ _9790_/CLK _9079_/D _9757_/SET_B VGND VGND VPWR VPWR _9079_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2 hold2/A VGND VGND VPWR VPWR hold2/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_58_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5800_ _9211_/Q _5799_/A _8846_/X _5799_/Y VGND VGND VPWR VPWR _9211_/D sky130_fd_sc_hd__a22o_1
X_6780_ _9491_/Q VGND VGND VPWR VPWR _6780_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_22_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5731_ _9055_/Q _7041_/A _5713_/Y VGND VGND VPWR VPWR _5731_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_188_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5662_ _5662_/A VGND VGND VPWR VPWR _5662_/Y sky130_fd_sc_hd__inv_2
X_8450_ _8450_/A VGND VGND VPWR VPWR _8683_/A sky130_fd_sc_hd__inv_2
X_8381_ _8722_/A _8381_/B VGND VGND VPWR VPWR _8382_/B sky130_fd_sc_hd__or2_1
X_5593_ _9312_/Q _5585_/A _8839_/X _5585_/Y VGND VGND VPWR VPWR _9312_/D sky130_fd_sc_hd__a22o_1
X_4613_ _5259_/A _4613_/B VGND VGND VPWR VPWR _4614_/A sky130_fd_sc_hd__or2_1
XFILLER_30_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7401_ _9252_/Q _7401_/B VGND VGND VPWR VPWR _7466_/A sky130_fd_sc_hd__or2_4
X_4544_ _9066_/Q VGND VGND VPWR VPWR _8810_/A sky130_fd_sc_hd__inv_2
XFILLER_163_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7332_ _6723_/Y _7086_/X _6695_/Y _7088_/X VGND VGND VPWR VPWR _7332_/X sky130_fd_sc_hd__o22a_1
XFILLER_190_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7263_ _6164_/Y _7124_/X _6163_/Y _7068_/B _7262_/X VGND VGND VPWR VPWR _7264_/D
+ sky130_fd_sc_hd__o221a_1
X_9002_ _9595_/Q _8781_/A VGND VGND VPWR VPWR mgmt_gpio_out[25] sky130_fd_sc_hd__ebufn_8
XFILLER_171_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4475_ _6052_/A VGND VGND VPWR VPWR _5259_/A sky130_fd_sc_hd__buf_12
XFILLER_104_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6214_ _9746_/Q VGND VGND VPWR VPWR _6214_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_143_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7194_ _8761_/A _7392_/B VGND VGND VPWR VPWR _7194_/X sky130_fd_sc_hd__or2_1
X_6145_ _6071_/Y _6145_/B _6145_/C _6145_/D VGND VGND VPWR VPWR _6145_/Y sky130_fd_sc_hd__nand4b_4
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6076_ _6074_/Y _5420_/B _6075_/Y _4861_/X VGND VGND VPWR VPWR _6076_/X sky130_fd_sc_hd__o22a_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5027_ _9687_/Q _5026_/A _8925_/A1 _5026_/Y VGND VGND VPWR VPWR _9687_/D sky130_fd_sc_hd__a22o_1
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9766_ _9769_/CLK _9766_/D _9757_/SET_B VGND VGND VPWR VPWR _9766_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_26_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6978_ _6237_/Y _6976_/A _9018_/Q _6976_/Y VGND VGND VPWR VPWR _9018_/D sky130_fd_sc_hd__o22a_1
X_8717_ _8640_/A _8164_/A _8640_/A _8640_/B VGND VGND VPWR VPWR _8717_/X sky130_fd_sc_hd__o22a_1
X_5929_ _7781_/A _7781_/B VGND VGND VPWR VPWR _7837_/C sky130_fd_sc_hd__or2_1
XFILLER_179_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9697_ _9709_/CLK _9697_/D _5004_/X VGND VGND VPWR VPWR _9697_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_166_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8648_ _8566_/B _8214_/Y _8340_/C VGND VGND VPWR VPWR _8681_/B sky130_fd_sc_hd__o21a_1
XFILLER_139_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8579_ _8708_/B _8579_/B _8579_/C VGND VGND VPWR VPWR _8716_/A sky130_fd_sc_hd__or3_2
XFILLER_181_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7950_ _8394_/D _8515_/B _8660_/C VGND VGND VPWR VPWR _8187_/A sky130_fd_sc_hd__or3_1
XFILLER_82_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7881_ _7881_/A VGND VGND VPWR VPWR _8566_/A sky130_fd_sc_hd__inv_2
X_6901_ _6901_/A _6901_/B _6901_/C _6901_/D VGND VGND VPWR VPWR _6945_/A sky130_fd_sc_hd__and4_1
X_6832_ _9521_/Q VGND VGND VPWR VPWR _6832_/Y sky130_fd_sc_hd__inv_6
XFILLER_35_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9620_ _9620_/CLK _9620_/D _9633_/SET_B VGND VGND VPWR VPWR _9620_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9551_ _9639_/CLK _9551_/D _9757_/SET_B VGND VGND VPWR VPWR _9551_/Q sky130_fd_sc_hd__dfrtp_1
X_6763_ _9444_/Q VGND VGND VPWR VPWR _6763_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9482_ _9483_/CLK _9482_/D _9685_/SET_B VGND VGND VPWR VPWR _9482_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_176_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6694_ _9530_/Q VGND VGND VPWR VPWR _6694_/Y sky130_fd_sc_hd__inv_2
X_8502_ _8230_/A _8498_/B _7877_/X _8233_/A VGND VGND VPWR VPWR _8504_/B sky130_fd_sc_hd__o211a_1
X_5714_ _7401_/B _9055_/Q _9251_/Q _5713_/Y VGND VGND VPWR VPWR _9251_/D sky130_fd_sc_hd__a22o_1
XFILLER_50_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8433_ _8514_/A _8433_/B VGND VGND VPWR VPWR _8636_/C sky130_fd_sc_hd__or2_1
X_5645_ _6997_/A _5643_/Y _5724_/B _9054_/Q _8819_/X VGND VGND VPWR VPWR _5658_/A
+ sky130_fd_sc_hd__a32o_2
XFILLER_40_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5576_ _9326_/Q _5574_/A _8845_/X _5574_/Y VGND VGND VPWR VPWR _9326_/D sky130_fd_sc_hd__a22o_1
X_8364_ _8364_/A _8730_/C _8575_/C _8364_/D VGND VGND VPWR VPWR _8368_/A sky130_fd_sc_hd__or4_1
X_8295_ _8295_/A _8295_/B VGND VGND VPWR VPWR _8296_/B sky130_fd_sc_hd__and2_1
XFILLER_116_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7315_ _6843_/Y _7097_/X _6845_/Y _7099_/X VGND VGND VPWR VPWR _7315_/X sky130_fd_sc_hd__o22a_1
X_4527_ _9769_/Q _4526_/A _8846_/X _4526_/Y VGND VGND VPWR VPWR _9769_/D sky130_fd_sc_hd__a22o_1
XFILLER_131_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7246_ _6160_/Y _7082_/X _6195_/Y _7084_/X _7245_/X VGND VGND VPWR VPWR _7265_/A
+ sky130_fd_sc_hd__o221a_1
X_4458_ _4661_/C _8938_/X _4665_/C VGND VGND VPWR VPWR _4459_/A sky130_fd_sc_hd__or3_1
X_7177_ _7177_/A _7177_/B _7177_/C VGND VGND VPWR VPWR _7177_/Y sky130_fd_sc_hd__nand3_4
XFILLER_77_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6128_ _9158_/Q VGND VGND VPWR VPWR _6128_/Y sky130_fd_sc_hd__inv_2
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6059_ _9100_/Q VGND VGND VPWR VPWR _6059_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_105 input86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_116 _8816_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_127 input91/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_138 _5259_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_149 _6787_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9749_ _9777_/CLK _9749_/D _9757_/SET_B VGND VGND VPWR VPWR _9749_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_41_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5430_ _9424_/Q _5422_/A _8839_/X _5422_/Y VGND VGND VPWR VPWR _9424_/D sky130_fd_sc_hd__a22o_1
XFILLER_145_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput315 _8817_/X VGND VGND VPWR VPWR spimemio_flash_io2_di sky130_fd_sc_hd__buf_2
X_5361_ _9472_/Q _5357_/A _8925_/A1 _5357_/Y VGND VGND VPWR VPWR _9472_/D sky130_fd_sc_hd__a22o_1
XFILLER_160_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput326 _9761_/Q VGND VGND VPWR VPWR sram_ro_csb sky130_fd_sc_hd__buf_2
Xoutput304 _9047_/Q VGND VGND VPWR VPWR pwr_ctrl_out[3] sky130_fd_sc_hd__buf_2
X_8080_ _8080_/A VGND VGND VPWR VPWR _8640_/B sky130_fd_sc_hd__buf_8
Xoutput348 _9040_/Q VGND VGND VPWR VPWR wb_dat_o[28] sky130_fd_sc_hd__buf_2
Xoutput337 _9030_/Q VGND VGND VPWR VPWR wb_dat_o[18] sky130_fd_sc_hd__buf_2
Xoutput359 _9013_/Q VGND VGND VPWR VPWR wb_dat_o[9] sky130_fd_sc_hd__buf_2
X_7100_ _4926_/Y _7097_/X _4910_/Y _7099_/X VGND VGND VPWR VPWR _7100_/X sky130_fd_sc_hd__o22a_1
XFILLER_99_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5292_ _5292_/A VGND VGND VPWR VPWR _5292_/Y sky130_fd_sc_hd__inv_2
X_7031_ _7127_/A _7111_/C VGND VGND VPWR VPWR _7109_/B sky130_fd_sc_hd__or2_1
XFILLER_101_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8982_ _9583_/Q _8745_/A VGND VGND VPWR VPWR mgmt_gpio_out[5] sky130_fd_sc_hd__ebufn_8
X_7933_ _8662_/A _7933_/B VGND VGND VPWR VPWR _7933_/X sky130_fd_sc_hd__or2_1
XFILLER_82_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7864_ _7864_/A VGND VGND VPWR VPWR _7864_/X sky130_fd_sc_hd__buf_6
XFILLER_23_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9603_ _9617_/CLK _9603_/D _9295_/SET_B VGND VGND VPWR VPWR _9603_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7795_ _8538_/C _8516_/B VGND VGND VPWR VPWR _8085_/A sky130_fd_sc_hd__or2_2
X_6815_ _6813_/Y _4870_/X _6814_/Y _4623_/B VGND VGND VPWR VPWR _6815_/X sky130_fd_sc_hd__o22a_1
X_9534_ _9534_/CLK _9534_/D _9647_/SET_B VGND VGND VPWR VPWR _9534_/Q sky130_fd_sc_hd__dfrtp_1
X_6746_ _6744_/Y _4841_/X _6745_/Y _5100_/B VGND VGND VPWR VPWR _6746_/X sky130_fd_sc_hd__o22a_1
XFILLER_50_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9465_ _9514_/CLK _9465_/D _4628_/A VGND VGND VPWR VPWR _9465_/Q sky130_fd_sc_hd__dfstp_1
X_6677_ _6675_/Y _4613_/B _6676_/Y _4868_/X VGND VGND VPWR VPWR _6677_/X sky130_fd_sc_hd__o22a_2
X_9396_ _9509_/CLK _9396_/D _9528_/SET_B VGND VGND VPWR VPWR _9396_/Q sky130_fd_sc_hd__dfrtp_1
X_5628_ _9289_/Q _5623_/A _8842_/X _5623_/Y VGND VGND VPWR VPWR _9289_/D sky130_fd_sc_hd__a22o_1
XFILLER_164_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8416_ _8416_/A VGND VGND VPWR VPWR _8667_/B sky130_fd_sc_hd__inv_2
X_8347_ _8377_/B _8350_/C VGND VGND VPWR VPWR _8347_/X sky130_fd_sc_hd__or2_2
XFILLER_164_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5559_ _9337_/Q _5558_/A _8843_/X _5558_/Y VGND VGND VPWR VPWR _9337_/D sky130_fd_sc_hd__a22o_1
XFILLER_117_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8278_ _8345_/A _8583_/C _8345_/B VGND VGND VPWR VPWR _8279_/A sky130_fd_sc_hd__or3b_1
X_7229_ _6264_/Y _7079_/B _6316_/Y _7059_/A VGND VGND VPWR VPWR _7229_/X sky130_fd_sc_hd__o22a_1
XFILLER_132_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_1_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A VGND VGND VPWR VPWR _9681_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_187_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4930_ _9489_/Q VGND VGND VPWR VPWR _4930_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_178_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4861_ _6111_/A _4925_/A VGND VGND VPWR VPWR _4861_/X sky130_fd_sc_hd__or2_4
X_6600_ _9069_/Q _6251_/Y _6599_/Y _4602_/B VGND VGND VPWR VPWR _6600_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_32_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_27 _4788_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_38 _6119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7580_ _6218_/Y _7425_/X _7577_/X _7579_/X VGND VGND VPWR VPWR _7590_/C sky130_fd_sc_hd__o211a_1
X_4792_ _9748_/Q VGND VGND VPWR VPWR _4792_/Y sky130_fd_sc_hd__inv_2
XANTENNA_16 _7536_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6531_ _6531_/A VGND VGND VPWR VPWR _6531_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_158_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_49 _6367_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6462_ _9692_/Q VGND VGND VPWR VPWR _6462_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9250_ _9279_/CLK _9250_/D _9633_/SET_B VGND VGND VPWR VPWR _9250_/Q sky130_fd_sc_hd__dfrtp_1
X_8201_ _8377_/C VGND VGND VPWR VPWR _8340_/C sky130_fd_sc_hd__inv_2
X_9181_ _9613_/CLK _9181_/D _9646_/SET_B VGND VGND VPWR VPWR _9181_/Q sky130_fd_sc_hd__dfrtp_1
X_6393_ _9306_/Q VGND VGND VPWR VPWR _6393_/Y sky130_fd_sc_hd__inv_2
X_5413_ _5413_/A VGND VGND VPWR VPWR _5414_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_173_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5344_ _5545_/A _5344_/B VGND VGND VPWR VPWR _5345_/A sky130_fd_sc_hd__or2_1
XFILLER_161_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8132_ _8164_/A _8137_/B VGND VGND VPWR VPWR _8133_/A sky130_fd_sc_hd__or2_1
X_5275_ _9530_/Q _5269_/A _8841_/X _5269_/Y VGND VGND VPWR VPWR _9530_/D sky130_fd_sc_hd__a22o_1
XFILLER_99_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8063_ _8077_/A VGND VGND VPWR VPWR _8518_/A sky130_fd_sc_hd__clkinv_4
X_7014_ _7014_/A VGND VGND VPWR VPWR _7014_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8965_ _7745_/X _8965_/A1 _8975_/S VGND VGND VPWR VPWR _8965_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8896_ _7397_/Y _9631_/Q _8959_/S VGND VGND VPWR VPWR _8896_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7916_ _8077_/A _8254_/B VGND VGND VPWR VPWR _8597_/A sky130_fd_sc_hd__nor2_1
XFILLER_169_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7847_ _7847_/A VGND VGND VPWR VPWR _8077_/A sky130_fd_sc_hd__buf_12
XFILLER_178_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7778_ _7756_/B _7777_/Y _7837_/B _7777_/A VGND VGND VPWR VPWR _7897_/A sky130_fd_sc_hd__o22a_1
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6729_ _9465_/Q VGND VGND VPWR VPWR _6729_/Y sky130_fd_sc_hd__clkinv_2
X_9517_ _9545_/CLK _9517_/D _4628_/A VGND VGND VPWR VPWR _9517_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_183_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9448_ _9785_/CLK _9448_/D _9779_/SET_B VGND VGND VPWR VPWR _9448_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_152_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9379_ _9379_/CLK _9379_/D _9779_/SET_B VGND VGND VPWR VPWR _9379_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_11_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput36 mgmt_gpio_in[0] VGND VGND VPWR VPWR _8805_/A sky130_fd_sc_hd__buf_8
Xinput14 mask_rev_in[19] VGND VGND VPWR VPWR _6570_/A sky130_fd_sc_hd__clkbuf_1
Xinput25 mask_rev_in[29] VGND VGND VPWR VPWR _6245_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_128_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput69 mgmt_gpio_in[6] VGND VGND VPWR VPWR input69/X sky130_fd_sc_hd__buf_2
Xinput47 mgmt_gpio_in[1] VGND VGND VPWR VPWR input47/X sky130_fd_sc_hd__clkbuf_4
Xinput58 mgmt_gpio_in[2] VGND VGND VPWR VPWR _4949_/A sky130_fd_sc_hd__buf_12
XFILLER_6_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5060_ _5060_/A VGND VGND VPWR VPWR _5060_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8750_ _8750_/A VGND VGND VPWR VPWR _8750_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_92_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5962_ _5962_/A VGND VGND VPWR VPWR _5962_/Y sky130_fd_sc_hd__inv_2
X_7701_ _7701_/A VGND VGND VPWR VPWR _7702_/A sky130_fd_sc_hd__clkbuf_1
X_4913_ _4906_/Y _4907_/X _4908_/Y _4577_/B _4912_/X VGND VGND VPWR VPWR _4934_/B
+ sky130_fd_sc_hd__o221a_2
XFILLER_18_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8681_ _8681_/A _8681_/B _8681_/C VGND VGND VPWR VPWR _8723_/A sky130_fd_sc_hd__or3_1
X_5893_ _5849_/A _8877_/X _8924_/X _9140_/Q VGND VGND VPWR VPWR _9140_/D sky130_fd_sc_hd__o22a_1
X_7632_ _6874_/Y _7434_/X _6843_/Y _7436_/X VGND VGND VPWR VPWR _7632_/X sky130_fd_sc_hd__o22a_1
X_4844_ _4919_/A _6158_/A VGND VGND VPWR VPWR _4844_/X sky130_fd_sc_hd__or2_1
XFILLER_193_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7563_ _6239_/Y _7445_/X _6269_/Y _7447_/X VGND VGND VPWR VPWR _7563_/X sky130_fd_sc_hd__o22a_1
X_4775_ _9120_/Q VGND VGND VPWR VPWR _4775_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_193_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9302_ _9440_/CLK _9302_/D _9685_/SET_B VGND VGND VPWR VPWR _9302_/Q sky130_fd_sc_hd__dfrtp_1
X_6514_ _9193_/Q VGND VGND VPWR VPWR _8749_/A sky130_fd_sc_hd__clkinv_4
X_9233_ _9508_/CLK _9233_/D _9647_/SET_B VGND VGND VPWR VPWR _9233_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_119_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7494_ _6933_/Y _7451_/X _6853_/Y _7453_/X _7493_/X VGND VGND VPWR VPWR _7499_/B
+ sky130_fd_sc_hd__o221a_1
X_6445_ _9645_/Q VGND VGND VPWR VPWR _6445_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6376_ _6371_/Y _5679_/B _6372_/Y _5776_/B _6375_/X VGND VGND VPWR VPWR _6376_/X
+ sky130_fd_sc_hd__o221a_1
X_9164_ _9203_/CLK _9164_/D _9633_/SET_B VGND VGND VPWR VPWR _9164_/Q sky130_fd_sc_hd__dfrtp_1
X_9095_ _9508_/CLK _9095_/D _9295_/SET_B VGND VGND VPWR VPWR _9095_/Q sky130_fd_sc_hd__dfrtp_1
X_5327_ _9494_/Q _5319_/A _8839_/X _5319_/Y VGND VGND VPWR VPWR _9494_/D sky130_fd_sc_hd__a22o_1
X_8115_ _8401_/A VGND VGND VPWR VPWR _8115_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8046_ _8624_/B _8554_/A VGND VGND VPWR VPWR _8467_/A sky130_fd_sc_hd__or2_1
XFILLER_75_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5258_ _9541_/Q _5253_/A _5967_/B1 _5253_/Y VGND VGND VPWR VPWR _9541_/D sky130_fd_sc_hd__a22o_1
X_5189_ _6040_/A VGND VGND VPWR VPWR _5190_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_113_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8948_ hold1/X _6237_/Y _8957_/S VGND VGND VPWR VPWR _8948_/X sky130_fd_sc_hd__mux2_1
XFILLER_188_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8879_ _8878_/X _9140_/Q _9054_/Q VGND VGND VPWR VPWR _8879_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4560_ _4560_/A VGND VGND VPWR VPWR _9757_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4491_ _5960_/A _4491_/B VGND VGND VPWR VPWR _4492_/A sky130_fd_sc_hd__or2_1
X_6230_ _9099_/Q VGND VGND VPWR VPWR _6230_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6161_ _6159_/Y _5382_/B _6160_/Y _5317_/B VGND VGND VPWR VPWR _6161_/X sky130_fd_sc_hd__o22a_1
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5112_ _5112_/A VGND VGND VPWR VPWR _5112_/Y sky130_fd_sc_hd__inv_2
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6092_ _9747_/Q VGND VGND VPWR VPWR _6092_/Y sky130_fd_sc_hd__inv_2
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5043_ _8970_/X _4551_/B _9676_/Q _5062_/D VGND VGND VPWR VPWR _9676_/D sky130_fd_sc_hd__a22o_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8802_ _8802_/A VGND VGND VPWR VPWR _8802_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9782_ _9785_/CLK _9782_/D _9779_/SET_B VGND VGND VPWR VPWR _9782_/Q sky130_fd_sc_hd__dfrtp_1
X_6994_ _6994_/A _9249_/Q VGND VGND VPWR VPWR _7075_/A sky130_fd_sc_hd__or2_4
X_8733_ _8733_/A VGND VGND VPWR VPWR _8733_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5945_ _9117_/Q _5943_/A _5964_/B1 _5943_/Y VGND VGND VPWR VPWR _9117_/D sky130_fd_sc_hd__a22o_1
XFILLER_25_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8664_ _8664_/A VGND VGND VPWR VPWR _8664_/X sky130_fd_sc_hd__clkbuf_1
X_5876_ _9157_/Q _5874_/A _8845_/X _5874_/Y VGND VGND VPWR VPWR _9157_/D sky130_fd_sc_hd__a22o_1
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7615_ _4775_/Y _7430_/X _4836_/Y _7432_/X _7614_/X VGND VGND VPWR VPWR _7615_/X
+ sky130_fd_sc_hd__o221a_1
X_4827_ _9203_/Q VGND VGND VPWR VPWR _4827_/Y sky130_fd_sc_hd__clkinv_2
X_8595_ _8595_/A _8595_/B _8595_/C _7902_/X VGND VGND VPWR VPWR _8659_/C sky130_fd_sc_hd__or4b_1
XFILLER_21_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4758_ _4749_/Y _5602_/B _4751_/Y _5545_/B _4757_/X VGND VGND VPWR VPWR _4790_/A
+ sky130_fd_sc_hd__o221a_1
X_7546_ _6368_/Y _7441_/X _6390_/Y _7443_/X _7545_/X VGND VGND VPWR VPWR _7553_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_5_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7477_ _7477_/A VGND VGND VPWR VPWR _7477_/X sky130_fd_sc_hd__buf_6
X_4689_ _6086_/B _4843_/B VGND VGND VPWR VPWR _5949_/B sky130_fd_sc_hd__or2_4
X_6428_ _9420_/Q VGND VGND VPWR VPWR _6428_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9216_ _9655_/CLK _9216_/D _9779_/SET_B VGND VGND VPWR VPWR _9216_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_68_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9147_ _9280_/CLK _9147_/D _9757_/SET_B VGND VGND VPWR VPWR _9147_/Q sky130_fd_sc_hd__dfrtp_1
X_6359_ _6359_/A1 _6165_/A _6356_/Y _5621_/B _6358_/X VGND VGND VPWR VPWR _6359_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_130_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9078_ _9790_/CLK _9078_/D _9757_/SET_B VGND VGND VPWR VPWR _9078_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_88_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8029_ _8624_/B _8550_/A VGND VGND VPWR VPWR _8029_/X sky130_fd_sc_hd__or2_1
XFILLER_29_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5730_ _5730_/A VGND VGND VPWR VPWR _9250_/D sky130_fd_sc_hd__inv_2
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5661_ _5661_/A VGND VGND VPWR VPWR _5662_/A sky130_fd_sc_hd__clkbuf_4
X_7400_ _7400_/A VGND VGND VPWR VPWR _7400_/X sky130_fd_sc_hd__buf_6
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8380_ _8380_/A _8380_/B _8720_/C _8585_/A VGND VGND VPWR VPWR _8381_/B sky130_fd_sc_hd__or4_1
X_5592_ _9313_/Q _5585_/A _8930_/A1 _5585_/Y VGND VGND VPWR VPWR _9313_/D sky130_fd_sc_hd__a22o_1
X_4612_ _6111_/A _6158_/B VGND VGND VPWR VPWR _4613_/B sky130_fd_sc_hd__or2_4
X_4543_ _9064_/Q VGND VGND VPWR VPWR _8811_/A sky130_fd_sc_hd__inv_2
X_7331_ _7331_/A _7331_/B _7331_/C VGND VGND VPWR VPWR _7331_/Y sky130_fd_sc_hd__nand3_4
XFILLER_190_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7262_ _6188_/Y _7126_/X _6189_/Y _7128_/X VGND VGND VPWR VPWR _7262_/X sky130_fd_sc_hd__o22a_1
X_9001_ _9594_/Q _8779_/A VGND VGND VPWR VPWR mgmt_gpio_out[24] sky130_fd_sc_hd__ebufn_8
XFILLER_171_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6213_ _8823_/X VGND VGND VPWR VPWR _6213_/Y sky130_fd_sc_hd__clkinv_2
X_4474_ _4729_/A _4729_/B _4669_/A _4729_/D VGND VGND VPWR VPWR _4891_/A sky130_fd_sc_hd__or4_4
X_7193_ _7703_/A _7059_/D _8767_/A _7116_/X _7192_/X VGND VGND VPWR VPWR _7198_/B
+ sky130_fd_sc_hd__o221a_1
X_6144_ _6144_/A _6144_/B _6144_/C _6144_/D VGND VGND VPWR VPWR _6145_/D sky130_fd_sc_hd__and4_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6075_ _6075_/A VGND VGND VPWR VPWR _6075_/Y sky130_fd_sc_hd__clkinv_4
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5026_ _5026_/A VGND VGND VPWR VPWR _5026_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6977_ _6145_/Y _6976_/A _9019_/Q _6976_/Y VGND VGND VPWR VPWR _9019_/D sky130_fd_sc_hd__o22a_1
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9765_ _9768_/CLK _9765_/D _4628_/A VGND VGND VPWR VPWR _9765_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_26_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5928_ _7774_/C _7774_/D _5928_/C VGND VGND VPWR VPWR _5936_/C sky130_fd_sc_hd__or3_1
X_8716_ _8716_/A _8716_/B _8716_/C _8716_/D VGND VGND VPWR VPWR _8729_/A sky130_fd_sc_hd__or4_1
XFILLER_179_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9696_ _8837_/A1 _9696_/D _5010_/X VGND VGND VPWR VPWR _9696_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_186_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8647_ _8647_/A _8716_/C _8678_/C _8721_/C VGND VGND VPWR VPWR _8647_/Y sky130_fd_sc_hd__nor4_1
XFILLER_21_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5859_ _5849_/X _8855_/X _8924_/X _9167_/Q VGND VGND VPWR VPWR _9167_/D sky130_fd_sc_hd__o22a_1
XFILLER_166_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8578_ _8578_/A _8578_/B _8578_/C VGND VGND VPWR VPWR _8645_/D sky130_fd_sc_hd__or3_1
XFILLER_147_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7529_ _8765_/A _7455_/X _6517_/Y _7457_/X VGND VGND VPWR VPWR _7529_/X sky130_fd_sc_hd__o22a_1
XFILLER_5_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7880_ _8394_/D _8272_/A VGND VGND VPWR VPWR _7881_/A sky130_fd_sc_hd__or2_2
X_6900_ _6895_/Y _5572_/B _6896_/Y _5897_/B _6899_/X VGND VGND VPWR VPWR _6901_/D
+ sky130_fd_sc_hd__o221a_1
X_6831_ _6831_/A VGND VGND VPWR VPWR _6831_/Y sky130_fd_sc_hd__clkinv_2
X_9550_ _9655_/CLK _9550_/D _9633_/SET_B VGND VGND VPWR VPWR _9550_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8501_ _8594_/A _8695_/C _8501_/C _8501_/D VGND VGND VPWR VPWR _8501_/X sky130_fd_sc_hd__or4_2
XFILLER_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6762_ _9543_/Q VGND VGND VPWR VPWR _6762_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_50_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9481_ _9527_/CLK _9481_/D _9685_/SET_B VGND VGND VPWR VPWR _9481_/Q sky130_fd_sc_hd__dfrtp_1
X_6693_ _9340_/Q VGND VGND VPWR VPWR _6693_/Y sky130_fd_sc_hd__clkinv_2
X_5713_ _5713_/A VGND VGND VPWR VPWR _5713_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_176_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8432_ _8562_/A _8672_/C _8432_/C VGND VGND VPWR VPWR _8434_/A sky130_fd_sc_hd__or3_1
X_5644_ _9055_/Q VGND VGND VPWR VPWR _5724_/B sky130_fd_sc_hd__clkinv_4
XFILLER_148_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8363_ _8627_/B _8490_/B VGND VGND VPWR VPWR _8364_/D sky130_fd_sc_hd__or2_1
XFILLER_156_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5575_ _9327_/Q _5574_/A _8846_/X _5574_/Y VGND VGND VPWR VPWR _9327_/D sky130_fd_sc_hd__a22o_1
X_7314_ _6883_/Y _7048_/B _6800_/Y _7077_/A _7313_/X VGND VGND VPWR VPWR _7321_/A
+ sky130_fd_sc_hd__o221a_1
X_8294_ _8294_/A _8650_/C VGND VGND VPWR VPWR _8295_/B sky130_fd_sc_hd__or2_1
XFILLER_116_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4526_ _4526_/A VGND VGND VPWR VPWR _4526_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7245_ _6178_/Y _7077_/C _6151_/Y _7077_/D _7244_/X VGND VGND VPWR VPWR _7245_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_116_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4457_ _4456_/Y _8942_/X _8941_/X VGND VGND VPWR VPWR _4665_/C sky130_fd_sc_hd__a21o_1
XFILLER_172_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7176_ _7176_/A _7176_/B _7176_/C _7176_/D VGND VGND VPWR VPWR _7177_/C sky130_fd_sc_hd__and4_1
X_6127_ _9113_/Q VGND VGND VPWR VPWR _6127_/Y sky130_fd_sc_hd__inv_2
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6058_ _9044_/Q _6054_/A _8916_/A1 _6054_/Y VGND VGND VPWR VPWR _9044_/D sky130_fd_sc_hd__a22o_1
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_106 input86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5009_ _6040_/A VGND VGND VPWR VPWR _5010_/A sky130_fd_sc_hd__clkbuf_1
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_128 mgmt_gpio_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_139 _4590_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_117 _8816_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9748_ _9755_/CLK _9748_/D _9757_/SET_B VGND VGND VPWR VPWR _9748_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_139_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9679_ _9681_/CLK _9679_/D _6146_/A VGND VGND VPWR VPWR _9679_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_182_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput316 _8818_/X VGND VGND VPWR VPWR spimemio_flash_io3_di sky130_fd_sc_hd__buf_2
X_5360_ _9473_/Q _5357_/A _8844_/X _5357_/Y VGND VGND VPWR VPWR _9473_/D sky130_fd_sc_hd__a22o_1
Xoutput305 _4808_/A VGND VGND VPWR VPWR reset sky130_fd_sc_hd__buf_2
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput349 _9041_/Q VGND VGND VPWR VPWR wb_dat_o[29] sky130_fd_sc_hd__buf_2
XFILLER_160_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput338 _9031_/Q VGND VGND VPWR VPWR wb_dat_o[19] sky130_fd_sc_hd__buf_2
XFILLER_126_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput327 _9119_/Q VGND VGND VPWR VPWR wb_ack_o sky130_fd_sc_hd__buf_2
X_5291_ _5291_/A VGND VGND VPWR VPWR _5292_/A sky130_fd_sc_hd__clkbuf_2
X_7030_ _7030_/A VGND VGND VPWR VPWR _7040_/A sky130_fd_sc_hd__buf_8
XFILLER_113_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8981_ _9582_/Q _7703_/A VGND VGND VPWR VPWR mgmt_gpio_out[4] sky130_fd_sc_hd__ebufn_8
X_7932_ _8394_/B _8298_/A _7931_/X VGND VGND VPWR VPWR _7933_/B sky130_fd_sc_hd__o21ai_1
XFILLER_82_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7863_ _8496_/A _8305_/A VGND VGND VPWR VPWR _7864_/A sky130_fd_sc_hd__or2_1
XFILLER_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9602_ _9617_/CLK _9602_/D _9295_/SET_B VGND VGND VPWR VPWR _9602_/Q sky130_fd_sc_hd__dfrtp_1
X_7794_ _7823_/A _7823_/B _8538_/B VGND VGND VPWR VPWR _8516_/B sky130_fd_sc_hd__o21ai_2
X_6814_ _9720_/Q VGND VGND VPWR VPWR _6814_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9533_ _9535_/CLK _9533_/D _9528_/SET_B VGND VGND VPWR VPWR _9533_/Q sky130_fd_sc_hd__dfrtp_1
X_6745_ _9643_/Q VGND VGND VPWR VPWR _6745_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_50_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9464_ _9514_/CLK _9464_/D _4628_/A VGND VGND VPWR VPWR _9464_/Q sky130_fd_sc_hd__dfrtp_1
X_6676_ _6676_/A VGND VGND VPWR VPWR _6676_/Y sky130_fd_sc_hd__inv_4
XFILLER_176_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8415_ _8551_/A _8401_/B _8412_/X _8414_/Y VGND VGND VPWR VPWR _8415_/X sky130_fd_sc_hd__o211a_1
XFILLER_191_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9395_ _9509_/CLK _9395_/D _9528_/SET_B VGND VGND VPWR VPWR _9395_/Q sky130_fd_sc_hd__dfrtp_1
X_5627_ _9290_/Q _5623_/A _8925_/A1 _5623_/Y VGND VGND VPWR VPWR _9290_/D sky130_fd_sc_hd__a22o_1
XFILLER_164_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8346_ _8346_/A _8346_/B _8196_/X VGND VGND VPWR VPWR _8350_/C sky130_fd_sc_hd__or3b_1
X_5558_ _5558_/A VGND VGND VPWR VPWR _5558_/Y sky130_fd_sc_hd__inv_2
X_8277_ _8525_/A _8189_/A _8213_/A _8583_/A _8189_/Y VGND VGND VPWR VPWR _8345_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_132_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4509_ _9775_/Q _4506_/A _5965_/B1 _4506_/Y VGND VGND VPWR VPWR _9775_/D sky130_fd_sc_hd__a22o_1
XFILLER_132_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7228_ _6290_/Y _7095_/X _6308_/Y _7068_/D _7227_/X VGND VGND VPWR VPWR _7233_/B
+ sky130_fd_sc_hd__o221a_1
X_5489_ _5489_/A VGND VGND VPWR VPWR _5490_/A sky130_fd_sc_hd__clkbuf_2
X_7159_ _6667_/Y _7040_/C _6754_/Y _7059_/C VGND VGND VPWR VPWR _7159_/X sky130_fd_sc_hd__o22a_1
XFILLER_86_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4860_ _4860_/A VGND VGND VPWR VPWR _4860_/Y sky130_fd_sc_hd__inv_2
X_4791_ _4791_/A _4791_/B _4791_/C _4791_/D VGND VGND VPWR VPWR _4936_/B sky130_fd_sc_hd__and4_1
XANTENNA_39 _6107_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6530_ _6528_/Y _5897_/B _6529_/Y _5024_/B VGND VGND VPWR VPWR _6530_/X sky130_fd_sc_hd__o22a_2
XANTENNA_17 _7572_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_28 _4833_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6461_ _9342_/Q VGND VGND VPWR VPWR _6461_/Y sky130_fd_sc_hd__inv_2
X_6392_ _9394_/Q VGND VGND VPWR VPWR _6392_/Y sky130_fd_sc_hd__inv_2
X_8200_ _8218_/A _8200_/B _8200_/C VGND VGND VPWR VPWR _8377_/C sky130_fd_sc_hd__or3_2
XFILLER_173_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9180_ _9613_/CLK _9180_/D _9646_/SET_B VGND VGND VPWR VPWR _9180_/Q sky130_fd_sc_hd__dfrtp_4
X_5412_ _5671_/A _5412_/B VGND VGND VPWR VPWR _5413_/A sky130_fd_sc_hd__or2_1
X_8131_ _8131_/A _8676_/A _8357_/A _8573_/A VGND VGND VPWR VPWR _8136_/A sky130_fd_sc_hd__or4_1
X_5343_ _9484_/Q _5338_/A _5967_/B1 _5338_/Y VGND VGND VPWR VPWR _9484_/D sky130_fd_sc_hd__a22o_1
XFILLER_99_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5274_ _9531_/Q _5269_/A _8929_/A1 _5269_/Y VGND VGND VPWR VPWR _9531_/D sky130_fd_sc_hd__a22o_1
X_8062_ _8062_/A _8062_/B VGND VGND VPWR VPWR _8065_/A sky130_fd_sc_hd__or2_1
XFILLER_114_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7013_ _7013_/A VGND VGND VPWR VPWR _7014_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8964_ _7743_/X _8964_/A1 _8975_/S VGND VGND VPWR VPWR _8964_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8895_ _8894_/X _9148_/Q _9054_/Q VGND VGND VPWR VPWR _8895_/X sky130_fd_sc_hd__mux2_1
X_7915_ _8226_/C _8319_/A VGND VGND VPWR VPWR _8254_/B sky130_fd_sc_hd__or2_1
X_7846_ _8394_/A _8394_/B _8394_/C _8195_/A VGND VGND VPWR VPWR _7847_/A sky130_fd_sc_hd__or4_1
XFILLER_70_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7777_ _7777_/A VGND VGND VPWR VPWR _7777_/Y sky130_fd_sc_hd__inv_2
XFILLER_184_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4989_ _9091_/Q _9090_/Q _9092_/Q VGND VGND VPWR VPWR _4989_/X sky130_fd_sc_hd__o21a_1
XFILLER_134_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6728_ _6723_/Y _5404_/B _6724_/Y _5496_/B _6727_/X VGND VGND VPWR VPWR _6741_/B
+ sky130_fd_sc_hd__o221a_1
X_9516_ _9771_/CLK _9516_/D _4628_/A VGND VGND VPWR VPWR _9516_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_7_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6659_ _4921_/A _6158_/A _6658_/Y _4481_/B _6158_/X VGND VGND VPWR VPWR _6659_/X
+ sky130_fd_sc_hd__o221a_1
X_9447_ _9791_/CLK _9447_/D _9633_/SET_B VGND VGND VPWR VPWR _9447_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_164_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9378_ _9378_/CLK _9378_/D _9646_/SET_B VGND VGND VPWR VPWR _9378_/Q sky130_fd_sc_hd__dfrtp_1
X_8329_ _8662_/A _8600_/A _8329_/C VGND VGND VPWR VPWR _8331_/A sky130_fd_sc_hd__or3_1
XFILLER_127_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput37 mgmt_gpio_in[10] VGND VGND VPWR VPWR input37/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput15 mask_rev_in[1] VGND VGND VPWR VPWR _6813_/A sky130_fd_sc_hd__clkbuf_1
Xinput26 mask_rev_in[2] VGND VGND VPWR VPWR _6706_/A sky130_fd_sc_hd__clkbuf_1
Xinput59 mgmt_gpio_in[30] VGND VGND VPWR VPWR _6193_/A sky130_fd_sc_hd__clkbuf_1
Xinput48 mgmt_gpio_in[20] VGND VGND VPWR VPWR _6450_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_143_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5961_ _5961_/A VGND VGND VPWR VPWR _5962_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8680_ _8716_/D _8731_/D _8680_/C _8720_/A VGND VGND VPWR VPWR _8680_/Y sky130_fd_sc_hd__nor4_2
X_7700_ _7700_/A VGND VGND VPWR VPWR _7700_/X sky130_fd_sc_hd__clkbuf_1
X_4912_ _6158_/A _4925_/A _4909_/Y _4910_/Y _5278_/B VGND VGND VPWR VPWR _4912_/X
+ sky130_fd_sc_hd__o32a_1
X_7631_ _6856_/Y _7427_/X _6938_/Y _5699_/X VGND VGND VPWR VPWR _7631_/X sky130_fd_sc_hd__o22a_1
X_5892_ _5849_/A _8879_/X _8924_/X _9141_/Q VGND VGND VPWR VPWR _9141_/D sky130_fd_sc_hd__o22a_1
XFILLER_33_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4843_ _4929_/A _4843_/B VGND VGND VPWR VPWR _5968_/B sky130_fd_sc_hd__or2_4
X_7562_ _6315_/Y _7425_/X _7559_/X _7561_/X VGND VGND VPWR VPWR _7572_/C sky130_fd_sc_hd__o211a_1
X_4774_ _6158_/B _4843_/B VGND VGND VPWR VPWR _5045_/B sky130_fd_sc_hd__or2_4
XFILLER_165_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9301_ _9788_/CLK _9301_/D _9295_/SET_B VGND VGND VPWR VPWR _9301_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_119_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7493_ _6793_/Y _7455_/X _6908_/Y _7457_/X VGND VGND VPWR VPWR _7493_/X sky130_fd_sc_hd__o22a_1
X_6513_ _6508_/Y _5556_/B _8763_/A _5572_/B _6512_/X VGND VGND VPWR VPWR _6526_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_20_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9232_ _9508_/CLK _9232_/D _9528_/SET_B VGND VGND VPWR VPWR _9232_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_146_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6444_ _6444_/A VGND VGND VPWR VPWR _6444_/Y sky130_fd_sc_hd__inv_2
X_9163_ _9532_/CLK _9163_/D _9647_/SET_B VGND VGND VPWR VPWR _9163_/Q sky130_fd_sc_hd__dfrtp_1
X_6375_ _6373_/Y _5789_/B _6374_/Y _5768_/B VGND VGND VPWR VPWR _6375_/X sky130_fd_sc_hd__o22a_1
X_9094_ _9501_/CLK _9094_/D _9647_/SET_B VGND VGND VPWR VPWR _9094_/Q sky130_fd_sc_hd__dfstp_1
X_5326_ _9495_/Q _5319_/A _8930_/A1 _5319_/Y VGND VGND VPWR VPWR _9495_/D sky130_fd_sc_hd__a22o_1
XFILLER_114_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8114_ _8164_/A VGND VGND VPWR VPWR _8114_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8045_ _8045_/A _8615_/B VGND VGND VPWR VPWR _8047_/A sky130_fd_sc_hd__nor2_1
X_5257_ _9542_/Q _5253_/A _5966_/B1 _5253_/Y VGND VGND VPWR VPWR _9542_/D sky130_fd_sc_hd__a22o_1
XFILLER_180_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5188_ _9587_/Q _5939_/A _5108_/X _4551_/X VGND VGND VPWR VPWR _9587_/D sky130_fd_sc_hd__a211o_1
XFILLER_68_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8947_ _9715_/Q _6326_/Y _8957_/S VGND VGND VPWR VPWR _8947_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8878_ _7199_/Y _9635_/Q _8959_/S VGND VGND VPWR VPWR _8878_/X sky130_fd_sc_hd__mux2_1
XFILLER_169_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7829_ _7829_/A VGND VGND VPWR VPWR _8376_/A sky130_fd_sc_hd__inv_2
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4490_ _4911_/A _4805_/A VGND VGND VPWR VPWR _4491_/B sky130_fd_sc_hd__or2_4
XFILLER_143_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6160_ _9500_/Q VGND VGND VPWR VPWR _6160_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5111_ _5111_/A VGND VGND VPWR VPWR _5112_/A sky130_fd_sc_hd__clkbuf_4
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6091_ _9379_/Q VGND VGND VPWR VPWR _6091_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_69_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5042_ _8971_/X _4551_/B _9677_/Q _5062_/D VGND VGND VPWR VPWR _9677_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8801_ _8801_/A _8801_/B VGND VGND VPWR VPWR _8802_/A sky130_fd_sc_hd__and2_1
XFILLER_65_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6993_ _9054_/Q _8819_/X _9054_/Q _6997_/C _9055_/Q VGND VGND VPWR VPWR _9054_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_25_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_51_csclk _9329_/CLK VGND VGND VPWR VPWR _9768_/CLK sky130_fd_sc_hd__clkbuf_16
X_9781_ _9785_/CLK _9781_/D _9779_/SET_B VGND VGND VPWR VPWR _9781_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_53_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8732_ _8732_/A VGND VGND VPWR VPWR _8732_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5944_ _9118_/Q _5943_/A _5963_/B1 _5943_/Y VGND VGND VPWR VPWR _9118_/D sky130_fd_sc_hd__a22o_1
XFILLER_18_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8663_ _8696_/C _8727_/C _8663_/C _8721_/A VGND VGND VPWR VPWR _8664_/A sky130_fd_sc_hd__or4_1
X_5875_ _9158_/Q _5874_/A _8846_/X _5874_/Y VGND VGND VPWR VPWR _9158_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8594_ _8594_/A _8594_/B _7896_/X VGND VGND VPWR VPWR _8595_/A sky130_fd_sc_hd__or3b_1
X_7614_ _4800_/Y _7434_/X _4930_/Y _7436_/X VGND VGND VPWR VPWR _7614_/X sky130_fd_sc_hd__o22a_1
XFILLER_21_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4826_ _6111_/A _4927_/A VGND VGND VPWR VPWR _5227_/B sky130_fd_sc_hd__or2_1
XFILLER_119_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7545_ _6357_/Y _7445_/X _6328_/Y _7447_/X VGND VGND VPWR VPWR _7545_/X sky130_fd_sc_hd__o22a_1
XFILLER_193_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4757_ _4787_/A _4891_/A _4753_/Y _4754_/Y _6135_/A VGND VGND VPWR VPWR _4757_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_119_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7476_ _7476_/A _9251_/Q _7476_/C _9255_/Q VGND VGND VPWR VPWR _7477_/A sky130_fd_sc_hd__or4_1
XFILLER_4_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4688_ _4729_/A _8944_/X _8934_/X _4729_/D VGND VGND VPWR VPWR _6086_/B sky130_fd_sc_hd__or4_4
XFILLER_146_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6427_ _9498_/Q VGND VGND VPWR VPWR _6427_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_108_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9215_ _9758_/CLK _9215_/D _9779_/SET_B VGND VGND VPWR VPWR _9215_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_161_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6358_ _9772_/Q _6251_/Y _6357_/Y _5420_/B VGND VGND VPWR VPWR _6358_/X sky130_fd_sc_hd__o2bb2a_1
X_9146_ _9280_/CLK _9146_/D _9757_/SET_B VGND VGND VPWR VPWR _9146_/Q sky130_fd_sc_hd__dfrtp_1
X_5309_ _9509_/Q _5308_/A _8846_/X _5308_/Y VGND VGND VPWR VPWR _9509_/D sky130_fd_sc_hd__a22o_1
XFILLER_102_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9077_ _9687_/CLK _9077_/D _9685_/SET_B VGND VGND VPWR VPWR _9077_/Q sky130_fd_sc_hd__dfrtp_1
X_6289_ _9753_/Q VGND VGND VPWR VPWR _6289_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_102_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8028_ _8521_/A _8550_/A VGND VGND VPWR VPWR _8410_/A sky130_fd_sc_hd__or2_1
XFILLER_124_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_19_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR _9509_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_17_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5660_ _6052_/A _5660_/B VGND VGND VPWR VPWR _5661_/A sky130_fd_sc_hd__or2_1
XFILLER_15_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4611_ _8934_/X _8932_/X _4729_/A _8944_/X VGND VGND VPWR VPWR _6158_/B sky130_fd_sc_hd__or4_4
XFILLER_175_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5591_ _9314_/Q _5585_/A _8841_/X _5585_/Y VGND VGND VPWR VPWR _9314_/D sky130_fd_sc_hd__a22o_1
X_4542_ _9065_/Q VGND VGND VPWR VPWR _7731_/A sky130_fd_sc_hd__clkinv_2
X_7330_ _7330_/A _7330_/B _7330_/C _7330_/D VGND VGND VPWR VPWR _7331_/C sky130_fd_sc_hd__and4_1
XFILLER_143_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7261_ _6200_/Y _5728_/X _6230_/Y _7040_/A _7260_/X VGND VGND VPWR VPWR _7264_/C
+ sky130_fd_sc_hd__o221a_1
X_4473_ _8932_/X VGND VGND VPWR VPWR _4729_/D sky130_fd_sc_hd__clkinv_2
X_9000_ _9568_/Q _8777_/A VGND VGND VPWR VPWR mgmt_gpio_out[23] sky130_fd_sc_hd__ebufn_8
X_6212_ _9157_/Q VGND VGND VPWR VPWR _6212_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_131_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7192_ _8779_/A _7118_/X _8799_/A _7048_/C VGND VGND VPWR VPWR _7192_/X sky130_fd_sc_hd__o22a_1
X_6143_ _7282_/A _5610_/B _6139_/Y _5679_/B _6142_/X VGND VGND VPWR VPWR _6144_/D
+ sky130_fd_sc_hd__o221a_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6074_ _9431_/Q VGND VGND VPWR VPWR _6074_/Y sky130_fd_sc_hd__clkinv_4
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5025_ _5025_/A VGND VGND VPWR VPWR _5026_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_85_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6976_ _6976_/A VGND VGND VPWR VPWR _6976_/Y sky130_fd_sc_hd__clkinv_2
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9764_ _9770_/CLK _9764_/D _7011_/B VGND VGND VPWR VPWR _9764_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_26_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5927_ _7771_/A _7771_/B _7771_/C _7771_/D VGND VGND VPWR VPWR _5928_/C sky130_fd_sc_hd__or4_1
XFILLER_110_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8715_ _8715_/A _8715_/B _8715_/C VGND VGND VPWR VPWR _8716_/B sky130_fd_sc_hd__or3_1
X_9695_ _9695_/CLK _9695_/D _9779_/SET_B VGND VGND VPWR VPWR _9695_/Q sky130_fd_sc_hd__dfrtp_1
X_8646_ _8646_/A _8646_/B VGND VGND VPWR VPWR _8678_/C sky130_fd_sc_hd__or2_1
XFILLER_139_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5858_ _5849_/X _8857_/X _8924_/X _9168_/Q VGND VGND VPWR VPWR _9168_/D sky130_fd_sc_hd__o22a_1
X_8577_ _8577_/A _8577_/B _8577_/C VGND VGND VPWR VPWR _8675_/C sky130_fd_sc_hd__or3_1
X_4809_ _9541_/Q VGND VGND VPWR VPWR _4809_/Y sky130_fd_sc_hd__clkinv_2
X_5789_ _5960_/A _5789_/B VGND VGND VPWR VPWR _5790_/A sky130_fd_sc_hd__or2_1
XFILLER_154_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7528_ _8755_/A _7441_/X _8791_/A _7443_/X _7527_/X VGND VGND VPWR VPWR _7535_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_5_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7459_ _4740_/Y _7451_/X _4916_/Y _7453_/X _7458_/X VGND VGND VPWR VPWR _7480_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_119_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9129_ _9129_/CLK _9129_/D _9779_/SET_B VGND VGND VPWR VPWR _9129_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6830_ _6830_/A _6830_/B _6830_/C _6830_/D VGND VGND VPWR VPWR _6946_/A sky130_fd_sc_hd__and4_1
XFILLER_62_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6761_ _9548_/Q VGND VGND VPWR VPWR _6761_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8500_ _8695_/A _8659_/A _8594_/B _7892_/X VGND VGND VPWR VPWR _8501_/D sky130_fd_sc_hd__or4b_1
X_5712_ _5724_/B _5704_/Y _5710_/Y _9252_/Q _5713_/A VGND VGND VPWR VPWR _9252_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_188_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9480_ _9527_/CLK _9480_/D _9685_/SET_B VGND VGND VPWR VPWR _9480_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_176_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6692_ _9780_/Q VGND VGND VPWR VPWR _6692_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8431_ _8431_/A _8431_/B VGND VGND VPWR VPWR _8432_/C sky130_fd_sc_hd__or2_1
X_5643_ _9056_/Q VGND VGND VPWR VPWR _5643_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5574_ _5574_/A VGND VGND VPWR VPWR _5574_/Y sky130_fd_sc_hd__inv_2
X_8362_ _8362_/A _8362_/B VGND VGND VPWR VPWR _8575_/C sky130_fd_sc_hd__or2_1
XFILLER_191_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7313_ _6940_/Y _7040_/C _6922_/Y _7059_/C VGND VGND VPWR VPWR _7313_/X sky130_fd_sc_hd__o22a_1
X_4525_ _4525_/A VGND VGND VPWR VPWR _4526_/A sky130_fd_sc_hd__clkbuf_4
X_8293_ _8377_/C _8204_/A _9067_/Q VGND VGND VPWR VPWR _8650_/C sky130_fd_sc_hd__o21ai_2
XFILLER_171_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7244_ _6159_/Y _7086_/X _6225_/Y _7088_/X VGND VGND VPWR VPWR _7244_/X sky130_fd_sc_hd__o22a_1
XFILLER_104_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4456_ _9587_/Q VGND VGND VPWR VPWR _4456_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7175_ _6767_/Y _7124_/X _6738_/Y _7068_/B _7174_/X VGND VGND VPWR VPWR _7176_/D
+ sky130_fd_sc_hd__o221a_1
X_6126_ _9225_/Q VGND VGND VPWR VPWR _6126_/Y sky130_fd_sc_hd__clkinv_2
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6057_ _9045_/Q _6054_/A _8930_/A1 _6054_/Y VGND VGND VPWR VPWR _9045_/D sky130_fd_sc_hd__a22o_1
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_107 input86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5008_ _5008_/A VGND VGND VPWR VPWR _9697_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_129 _6485_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_118 _8816_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6959_ _6946_/Y _6952_/A _9029_/Q _6952_/Y VGND VGND VPWR VPWR _9029_/D sky130_fd_sc_hd__o22a_1
X_9747_ _9777_/CLK _9747_/D _9757_/SET_B VGND VGND VPWR VPWR _9747_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_53_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9678_ _9681_/CLK _9678_/D _6146_/A VGND VGND VPWR VPWR _9678_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8629_ _8710_/A _8629_/B _8686_/D _8628_/X VGND VGND VPWR VPWR _8633_/A sky130_fd_sc_hd__or4b_2
XFILLER_182_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput306 _8802_/X VGND VGND VPWR VPWR ser_rx sky130_fd_sc_hd__buf_2
Xoutput317 _9762_/Q VGND VGND VPWR VPWR sram_ro_addr[0] sky130_fd_sc_hd__buf_2
XFILLER_126_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput339 _9021_/Q VGND VGND VPWR VPWR wb_dat_o[1] sky130_fd_sc_hd__buf_2
Xoutput328 _9020_/Q VGND VGND VPWR VPWR wb_dat_o[0] sky130_fd_sc_hd__buf_2
X_5290_ _5671_/A _5290_/B VGND VGND VPWR VPWR _5291_/A sky130_fd_sc_hd__or2_1
XFILLER_141_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8980_ _9581_/Q _7705_/A VGND VGND VPWR VPWR mgmt_gpio_out[3] sky130_fd_sc_hd__ebufn_8
X_7931_ _7931_/A _7931_/B VGND VGND VPWR VPWR _7931_/X sky130_fd_sc_hd__and2_1
XFILLER_82_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9601_ _9601_/CLK _9601_/D _9295_/SET_B VGND VGND VPWR VPWR _9601_/Q sky130_fd_sc_hd__dfrtp_1
X_7862_ _8260_/A VGND VGND VPWR VPWR _7862_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7793_ _8189_/A _7791_/B _7792_/B VGND VGND VPWR VPWR _8538_/B sky130_fd_sc_hd__a21o_2
XFILLER_90_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6813_ _6813_/A VGND VGND VPWR VPWR _6813_/Y sky130_fd_sc_hd__inv_2
X_9532_ _9532_/CLK _9532_/D _9647_/SET_B VGND VGND VPWR VPWR _9532_/Q sky130_fd_sc_hd__dfrtp_1
X_6744_ _6744_/A VGND VGND VPWR VPWR _6744_/Y sky130_fd_sc_hd__inv_2
XFILLER_167_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9463_ _9514_/CLK _9463_/D _4628_/A VGND VGND VPWR VPWR _9463_/Q sky130_fd_sc_hd__dfrtp_1
X_6675_ _9723_/Q VGND VGND VPWR VPWR _6675_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5626_ _9291_/Q _5623_/A _8844_/X _5623_/Y VGND VGND VPWR VPWR _9291_/D sky130_fd_sc_hd__a22o_1
XFILLER_164_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8414_ _8627_/C VGND VGND VPWR VPWR _8414_/Y sky130_fd_sc_hd__inv_2
X_9394_ _9483_/CLK _9394_/D _9528_/SET_B VGND VGND VPWR VPWR _9394_/Q sky130_fd_sc_hd__dfrtp_1
X_8345_ _8345_/A _8345_/B VGND VGND VPWR VPWR _8377_/B sky130_fd_sc_hd__or2_1
X_5557_ _5557_/A VGND VGND VPWR VPWR _5558_/A sky130_fd_sc_hd__clkbuf_2
X_8276_ _8660_/A _8660_/B _8496_/A VGND VGND VPWR VPWR _8280_/B sky130_fd_sc_hd__or3_2
X_5488_ _5671_/A _5488_/B VGND VGND VPWR VPWR _5489_/A sky130_fd_sc_hd__or2_1
X_4508_ _9776_/Q _4506_/A _5964_/B1 _4506_/Y VGND VGND VPWR VPWR _9776_/D sky130_fd_sc_hd__a22o_1
XFILLER_132_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7227_ _6240_/Y _7097_/X _6271_/Y _7099_/X VGND VGND VPWR VPWR _7227_/X sky130_fd_sc_hd__o22a_1
XFILLER_116_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7158_ _6717_/Y _7082_/X _6704_/Y _7084_/X _7157_/X VGND VGND VPWR VPWR _7177_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_98_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6109_ _9535_/Q VGND VGND VPWR VPWR _6109_/Y sky130_fd_sc_hd__inv_2
X_7089_ _4916_/Y _7086_/X _4914_/Y _7088_/X VGND VGND VPWR VPWR _7089_/X sky130_fd_sc_hd__o22a_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4790_ _4790_/A _4790_/B _4790_/C _4790_/D VGND VGND VPWR VPWR _4791_/D sky130_fd_sc_hd__and4_1
XANTENNA_18 _7608_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_29 _4835_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6460_ _8808_/B _6134_/A _6456_/Y _5949_/B _6459_/X VGND VGND VPWR VPWR _6473_/B
+ sky130_fd_sc_hd__o221a_1
X_6391_ _9462_/Q VGND VGND VPWR VPWR _6391_/Y sky130_fd_sc_hd__inv_2
X_5411_ _9437_/Q _5406_/A _5967_/B1 _5406_/Y VGND VGND VPWR VPWR _9437_/D sky130_fd_sc_hd__a22o_1
XFILLER_161_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8130_ _8213_/A _8130_/B VGND VGND VPWR VPWR _8573_/A sky130_fd_sc_hd__nor2_1
X_5342_ _9485_/Q _5338_/A _5966_/B1 _5338_/Y VGND VGND VPWR VPWR _9485_/D sky130_fd_sc_hd__a22o_1
X_8061_ _8061_/A _8064_/B _8061_/C VGND VGND VPWR VPWR _8062_/B sky130_fd_sc_hd__and3_1
XFILLER_99_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5273_ _9532_/Q _5269_/A _8843_/X _5269_/Y VGND VGND VPWR VPWR _9532_/D sky130_fd_sc_hd__a22o_1
XFILLER_114_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7012_ _9626_/Q input86/X VGND VGND VPWR VPWR _7013_/A sky130_fd_sc_hd__or2b_1
XFILLER_68_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8963_ _7741_/X _8963_/A1 _8975_/S VGND VGND VPWR VPWR _8963_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8894_ _7375_/Y _9630_/Q _8959_/S VGND VGND VPWR VPWR _8894_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7914_ _8521_/B _8246_/B VGND VGND VPWR VPWR _8317_/A sky130_fd_sc_hd__nor2_1
X_7845_ _7845_/A VGND VGND VPWR VPWR _8305_/A sky130_fd_sc_hd__buf_8
XFILLER_169_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7776_ _8189_/A _7791_/B _7966_/A _7966_/C VGND VGND VPWR VPWR _7777_/A sky130_fd_sc_hd__or4_1
XFILLER_178_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4988_ _9700_/Q _9699_/Q VGND VGND VPWR VPWR _5992_/B sky130_fd_sc_hd__nor2_1
XFILLER_51_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9515_ _9545_/CLK _9515_/D _4628_/A VGND VGND VPWR VPWR _9515_/Q sky130_fd_sc_hd__dfrtp_1
X_6727_ _6725_/Y _5232_/B _6726_/Y _4822_/X VGND VGND VPWR VPWR _6727_/X sky130_fd_sc_hd__o22a_2
XFILLER_176_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6658_ _9788_/Q VGND VGND VPWR VPWR _6658_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_127_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9446_ _9791_/CLK _9446_/D _9779_/SET_B VGND VGND VPWR VPWR _9446_/Q sky130_fd_sc_hd__dfrtp_1
X_5609_ _9302_/Q _5604_/A _5967_/B1 _5604_/Y VGND VGND VPWR VPWR _9302_/D sky130_fd_sc_hd__a22o_1
X_9377_ _9378_/CLK _9377_/D _9646_/SET_B VGND VGND VPWR VPWR _9377_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_152_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8328_ _7848_/A _8300_/B _8327_/Y VGND VGND VPWR VPWR _8329_/C sky130_fd_sc_hd__o21ai_1
X_6589_ _9466_/Q VGND VGND VPWR VPWR _6589_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8259_ _8259_/A _8367_/B VGND VGND VPWR VPWR _8261_/A sky130_fd_sc_hd__or2_1
XFILLER_120_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput16 mask_rev_in[20] VGND VGND VPWR VPWR _6385_/A sky130_fd_sc_hd__clkbuf_1
Xinput27 mask_rev_in[30] VGND VGND VPWR VPWR _6207_/A sky130_fd_sc_hd__clkbuf_1
Xinput49 mgmt_gpio_in[21] VGND VGND VPWR VPWR input49/X sky130_fd_sc_hd__clkbuf_4
Xinput38 mgmt_gpio_in[11] VGND VGND VPWR VPWR _6505_/A sky130_fd_sc_hd__buf_6
XFILLER_182_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5960_ _5960_/A _5960_/B VGND VGND VPWR VPWR _5961_/A sky130_fd_sc_hd__or2_1
XFILLER_93_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5891_ _5849_/A _8881_/X _8924_/X _9142_/Q VGND VGND VPWR VPWR _9142_/D sky130_fd_sc_hd__o22a_1
X_4911_ _4911_/A _6086_/B VGND VGND VPWR VPWR _5278_/B sky130_fd_sc_hd__or2_4
X_7630_ _6932_/Y _7415_/X _6800_/Y _7417_/X _7629_/X VGND VGND VPWR VPWR _7644_/B
+ sky130_fd_sc_hd__o221a_1
X_4842_ _9093_/Q VGND VGND VPWR VPWR _4842_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_119_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7561_ _6304_/Y _7430_/X _6263_/Y _7432_/X _7560_/X VGND VGND VPWR VPWR _7561_/X
+ sky130_fd_sc_hd__o221a_1
X_4773_ _9667_/Q VGND VGND VPWR VPWR _4773_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9300_ _9788_/CLK _9300_/D _9295_/SET_B VGND VGND VPWR VPWR _9300_/Q sky130_fd_sc_hd__dfrtp_1
X_7492_ _6939_/Y _7441_/X _6787_/Y _7443_/X _7491_/X VGND VGND VPWR VPWR _7499_/A
+ sky130_fd_sc_hd__o221a_1
X_6512_ _6510_/Y _5671_/B _8753_/A _5776_/B VGND VGND VPWR VPWR _6512_/X sky130_fd_sc_hd__o22a_1
X_9231_ _9508_/CLK _9231_/D _9528_/SET_B VGND VGND VPWR VPWR _9231_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_119_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6443_ _6438_/Y _4841_/X _6439_/Y _5089_/B _6442_/X VGND VGND VPWR VPWR _6443_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_106_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9162_ _9358_/CLK _9162_/D _9685_/SET_B VGND VGND VPWR VPWR _9162_/Q sky130_fd_sc_hd__dfrtp_1
X_6374_ _9230_/Q VGND VGND VPWR VPWR _6374_/Y sky130_fd_sc_hd__inv_2
XFILLER_142_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9093_ _9501_/CLK _9093_/D _9647_/SET_B VGND VGND VPWR VPWR _9093_/Q sky130_fd_sc_hd__dfstp_1
X_5325_ _9496_/Q _5319_/A _8841_/X _5319_/Y VGND VGND VPWR VPWR _9496_/D sky130_fd_sc_hd__a22o_1
XFILLER_102_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8113_ _8401_/A _8378_/B VGND VGND VPWR VPWR _8354_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8044_ _8521_/A _8554_/A VGND VGND VPWR VPWR _8615_/B sky130_fd_sc_hd__nor2_1
X_5256_ _9543_/Q _5253_/A _5965_/B1 _5253_/Y VGND VGND VPWR VPWR _9543_/D sky130_fd_sc_hd__a22o_1
XFILLER_102_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5187_ _9059_/Q VGND VGND VPWR VPWR _5939_/A sky130_fd_sc_hd__inv_2
XFILLER_68_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8946_ _8945_/X _9676_/Q _9587_/Q VGND VGND VPWR VPWR _8946_/X sky130_fd_sc_hd__mux2_4
XFILLER_56_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8877_ _8876_/X _9139_/Q _9054_/Q VGND VGND VPWR VPWR _8877_/X sky130_fd_sc_hd__mux2_1
X_7828_ _8097_/B _8660_/B _8660_/C VGND VGND VPWR VPWR _7829_/A sky130_fd_sc_hd__or3_1
X_7759_ _8525_/A _7894_/B _7903_/C _8528_/A VGND VGND VPWR VPWR _8394_/D sky130_fd_sc_hd__or4_4
XFILLER_11_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9429_ _9508_/CLK _9429_/D _9295_/SET_B VGND VGND VPWR VPWR _9429_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_137_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5110_ _5545_/A _5110_/B VGND VGND VPWR VPWR _5111_/A sky130_fd_sc_hd__or2_1
X_6090_ _9405_/Q VGND VGND VPWR VPWR _6090_/Y sky130_fd_sc_hd__inv_2
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5041_ _8972_/X _4551_/B _9678_/Q _5062_/D VGND VGND VPWR VPWR _9678_/D sky130_fd_sc_hd__a22o_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8800_ _8800_/A VGND VGND VPWR VPWR _8800_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0_wb_clk_i wb_clk_i VGND VGND VPWR VPWR clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_65_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9780_ _9785_/CLK _9780_/D _9779_/SET_B VGND VGND VPWR VPWR _9780_/Q sky130_fd_sc_hd__dfrtp_1
X_8731_ _8731_/A _8731_/B _8731_/C _8731_/D VGND VGND VPWR VPWR _8731_/X sky130_fd_sc_hd__or4_1
XFILLER_80_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6992_ _5643_/Y _5753_/B _9053_/Q _6991_/Y VGND VGND VPWR VPWR _9053_/D sky130_fd_sc_hd__a2bb2o_1
X_5943_ _5943_/A VGND VGND VPWR VPWR _5943_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8662_ _8662_/A _8662_/B _8662_/C _8661_/X VGND VGND VPWR VPWR _8663_/C sky130_fd_sc_hd__or4b_2
X_5874_ _5874_/A VGND VGND VPWR VPWR _5874_/Y sky130_fd_sc_hd__inv_2
X_8593_ _7836_/B _8591_/Y _8641_/A _8501_/C VGND VGND VPWR VPWR _8695_/D sky130_fd_sc_hd__a211o_1
X_7613_ _4858_/Y _7427_/X _4718_/Y _5699_/X VGND VGND VPWR VPWR _7613_/X sky130_fd_sc_hd__o22a_2
X_4825_ _9559_/Q VGND VGND VPWR VPWR _8807_/A sky130_fd_sc_hd__inv_2
XFILLER_193_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7544_ _6456_/Y _7425_/X _7541_/X _7543_/X VGND VGND VPWR VPWR _7554_/C sky130_fd_sc_hd__o211a_1
XFILLER_193_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4756_ _4756_/A VGND VGND VPWR VPWR _6135_/A sky130_fd_sc_hd__buf_8
XFILLER_162_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4687_ _9106_/Q VGND VGND VPWR VPWR _4687_/Y sky130_fd_sc_hd__clkinv_2
X_7475_ _7475_/A VGND VGND VPWR VPWR _7475_/X sky130_fd_sc_hd__buf_8
XFILLER_161_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6426_ _6421_/Y _5496_/B _6422_/Y _5393_/B _6425_/X VGND VGND VPWR VPWR _6433_/C
+ sky130_fd_sc_hd__o221a_1
X_9214_ _9655_/CLK _9214_/D _9779_/SET_B VGND VGND VPWR VPWR _9214_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_161_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6357_ _9428_/Q VGND VGND VPWR VPWR _6357_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9145_ _9203_/CLK _9145_/D _9633_/SET_B VGND VGND VPWR VPWR _9145_/Q sky130_fd_sc_hd__dfrtp_1
X_5308_ _5308_/A VGND VGND VPWR VPWR _5308_/Y sky130_fd_sc_hd__inv_2
XFILLER_161_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9076_ _9687_/CLK _9076_/D _9685_/SET_B VGND VGND VPWR VPWR _9076_/Q sky130_fd_sc_hd__dfrtp_1
X_6288_ _9209_/Q VGND VGND VPWR VPWR _6288_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8027_ _8389_/A _8137_/B _8097_/B _8137_/B _8026_/X VGND VGND VPWR VPWR _8027_/X
+ sky130_fd_sc_hd__o221a_1
X_5239_ _9554_/Q _5234_/A _5967_/B1 _5234_/Y VGND VGND VPWR VPWR _9554_/D sky130_fd_sc_hd__a22o_1
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8929_ _9613_/Q _8929_/A1 _8930_/S VGND VGND VPWR VPWR _8929_/X sky130_fd_sc_hd__mux2_1
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4610_ _9726_/Q _4604_/A _5967_/B1 _4604_/Y VGND VGND VPWR VPWR _9726_/D sky130_fd_sc_hd__a22o_1
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5590_ _9315_/Q _5585_/A _8929_/A1 _5585_/Y VGND VGND VPWR VPWR _9315_/D sky130_fd_sc_hd__a22o_1
XFILLER_30_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4541_ _4541_/A VGND VGND VPWR VPWR _9760_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7260_ _7260_/A _7392_/B VGND VGND VPWR VPWR _7260_/X sky130_fd_sc_hd__or2_1
X_4472_ _8934_/X VGND VGND VPWR VPWR _4669_/A sky130_fd_sc_hd__clkinv_2
X_6211_ _6211_/A _6211_/B _6211_/C _6211_/D VGND VGND VPWR VPWR _6237_/C sky130_fd_sc_hd__and4_1
XFILLER_104_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7191_ _8747_/A _7040_/D _8765_/A _7110_/X _7190_/X VGND VGND VPWR VPWR _7198_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_143_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6142_ _6140_/Y _5818_/B _6141_/Y _5572_/B VGND VGND VPWR VPWR _6142_/X sky130_fd_sc_hd__o22a_1
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6073_ _9501_/Q VGND VGND VPWR VPWR _6073_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _5259_/A _5024_/B VGND VGND VPWR VPWR _5025_/A sky130_fd_sc_hd__or2_2
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6975_ _6975_/A VGND VGND VPWR VPWR _6976_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9763_ _9770_/CLK _9763_/D _7011_/B VGND VGND VPWR VPWR _9763_/Q sky130_fd_sc_hd__dfrtp_2
X_5926_ _7770_/A _7770_/B _7768_/A _7768_/B VGND VGND VPWR VPWR _5936_/B sky130_fd_sc_hd__or4_1
X_8714_ _8714_/A _8714_/B _8714_/C _8714_/D VGND VGND VPWR VPWR _8739_/A sky130_fd_sc_hd__or4_1
XFILLER_80_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9694_ _9695_/CLK _9694_/D _9779_/SET_B VGND VGND VPWR VPWR _9694_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_34_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8645_ _8645_/A _8645_/B _8645_/C _8645_/D VGND VGND VPWR VPWR _8716_/C sky130_fd_sc_hd__or4_4
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5857_ _5849_/X _8859_/X _8924_/X _9169_/Q VGND VGND VPWR VPWR _9169_/D sky130_fd_sc_hd__o22a_1
XFILLER_186_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8576_ _8576_/A _8642_/D _8730_/D _8576_/D VGND VGND VPWR VPWR _8580_/A sky130_fd_sc_hd__or4_1
X_5788_ _9277_/Q _9056_/Q _5787_/Y _9217_/Q _5755_/A VGND VGND VPWR VPWR _9217_/D
+ sky130_fd_sc_hd__a32o_1
X_4808_ _4808_/A VGND VGND VPWR VPWR _4808_/Y sky130_fd_sc_hd__inv_2
X_4739_ _4739_/A VGND VGND VPWR VPWR _6134_/A sky130_fd_sc_hd__buf_6
X_7527_ _8771_/A _7445_/X _8769_/A _7447_/X VGND VGND VPWR VPWR _7527_/X sky130_fd_sc_hd__o22a_1
X_7458_ _4804_/Y _7455_/X _4769_/Y _7457_/X VGND VGND VPWR VPWR _7458_/X sky130_fd_sc_hd__o22a_1
X_6409_ _9415_/Q VGND VGND VPWR VPWR _6409_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_135_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7389_ _6434_/Y _7040_/D _6363_/Y _7110_/X _7388_/X VGND VGND VPWR VPWR _7396_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_135_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9128_ _9379_/CLK _9128_/D _9779_/SET_B VGND VGND VPWR VPWR _9128_/Q sky130_fd_sc_hd__dfrtp_1
X_9059_ _4450_/A1 _9059_/D _6146_/A VGND VGND VPWR VPWR _9059_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_50_csclk _9329_/CLK VGND VGND VPWR VPWR _9770_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6760_ _9504_/Q VGND VGND VPWR VPWR _6760_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_90_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5711_ _9053_/Q _9055_/Q VGND VGND VPWR VPWR _5713_/A sky130_fd_sc_hd__or2_1
X_6691_ _6691_/A _6691_/B _6691_/C _6691_/D VGND VGND VPWR VPWR _6785_/B sky130_fd_sc_hd__and4_1
X_8430_ _8430_/A _8560_/B VGND VGND VPWR VPWR _8431_/B sky130_fd_sc_hd__or2_1
X_5642_ _9054_/Q VGND VGND VPWR VPWR _6997_/A sky130_fd_sc_hd__inv_2
XFILLER_176_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5573_ _5573_/A VGND VGND VPWR VPWR _5574_/A sky130_fd_sc_hd__clkbuf_4
X_8361_ _8361_/A _8361_/B VGND VGND VPWR VPWR _8730_/C sky130_fd_sc_hd__or2_1
X_7312_ _6848_/Y _7082_/X _6824_/Y _7084_/X _7311_/X VGND VGND VPWR VPWR _7331_/A
+ sky130_fd_sc_hd__o221a_1
X_4524_ _5960_/A _4524_/B VGND VGND VPWR VPWR _4525_/A sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_18_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR _9483_/CLK sky130_fd_sc_hd__clkbuf_16
X_8292_ _8514_/A _8292_/B VGND VGND VPWR VPWR _8294_/A sky130_fd_sc_hd__nor2_1
XFILLER_132_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7243_ _7243_/A _7243_/B _7243_/C VGND VGND VPWR VPWR _7243_/Y sky130_fd_sc_hd__nand3_4
XFILLER_104_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4455_ _8936_/X VGND VGND VPWR VPWR _4661_/C sky130_fd_sc_hd__inv_2
XFILLER_104_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7174_ _6650_/Y _7126_/X _6692_/Y _7128_/X VGND VGND VPWR VPWR _7174_/X sky130_fd_sc_hd__o22a_1
XFILLER_131_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6125_ _6120_/Y _5013_/B _6121_/Y _5797_/B _6124_/X VGND VGND VPWR VPWR _6144_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_105_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6056_ _9046_/Q _6054_/A _8955_/A1 _6054_/Y VGND VGND VPWR VPWR _9046_/D sky130_fd_sc_hd__a22o_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5007_ _4949_/A _9697_/Q _5007_/S VGND VGND VPWR VPWR _5008_/A sky130_fd_sc_hd__mux2_1
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_119 _8816_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_108 input86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9746_ _9777_/CLK _9746_/D _9757_/SET_B VGND VGND VPWR VPWR _9746_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_186_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6958_ _6785_/Y _6952_/A _9030_/Q _6952_/Y VGND VGND VPWR VPWR _9030_/D sky130_fd_sc_hd__o22a_1
XFILLER_157_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6889_ _9152_/Q VGND VGND VPWR VPWR _6889_/Y sky130_fd_sc_hd__clkinv_2
X_5909_ _9131_/Q _5907_/A _8845_/X _5907_/Y VGND VGND VPWR VPWR _9131_/D sky130_fd_sc_hd__a22o_1
XFILLER_14_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9677_ _9681_/CLK _9677_/D _6146_/A VGND VGND VPWR VPWR _9677_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8628_ _8130_/B _8554_/B _8454_/B _8133_/A _8408_/Y VGND VGND VPWR VPWR _8628_/X
+ sky130_fd_sc_hd__o2111a_1
X_8559_ _8559_/A _8709_/A _8631_/B _8688_/B VGND VGND VPWR VPWR _8563_/A sky130_fd_sc_hd__or4_1
XFILLER_108_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput307 _8819_/X VGND VGND VPWR VPWR serial_clock sky130_fd_sc_hd__buf_2
Xoutput329 _9014_/Q VGND VGND VPWR VPWR wb_dat_o[10] sky130_fd_sc_hd__buf_2
XFILLER_126_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput318 _9763_/Q VGND VGND VPWR VPWR sram_ro_addr[1] sky130_fd_sc_hd__buf_2
XFILLER_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7930_ _7848_/A _8305_/A _7929_/Y VGND VGND VPWR VPWR _7931_/B sky130_fd_sc_hd__o21ba_1
XFILLER_67_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7861_ _8305_/A VGND VGND VPWR VPWR _8299_/B sky130_fd_sc_hd__inv_2
XFILLER_63_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9600_ _9601_/CLK _9600_/D _9295_/SET_B VGND VGND VPWR VPWR _9600_/Q sky130_fd_sc_hd__dfrtp_1
X_6812_ _9774_/Q VGND VGND VPWR VPWR _6812_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_168_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7792_ _8525_/A _7792_/B VGND VGND VPWR VPWR _7823_/B sky130_fd_sc_hd__nor2_1
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9531_ _9535_/CLK _9531_/D _9528_/SET_B VGND VGND VPWR VPWR _9531_/Q sky130_fd_sc_hd__dfrtp_4
X_6743_ _9122_/Q VGND VGND VPWR VPWR _6743_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_176_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6674_ _9161_/Q VGND VGND VPWR VPWR _6674_/Y sky130_fd_sc_hd__inv_2
X_9462_ _9532_/CLK _9462_/D _9647_/SET_B VGND VGND VPWR VPWR _9462_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5625_ _9292_/Q _5623_/A _8845_/X _5623_/Y VGND VGND VPWR VPWR _9292_/D sky130_fd_sc_hd__a22o_1
X_8413_ _8614_/B _8575_/A VGND VGND VPWR VPWR _8627_/C sky130_fd_sc_hd__or2_1
X_9393_ _9509_/CLK _9393_/D _9528_/SET_B VGND VGND VPWR VPWR _9393_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_176_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8344_ _8279_/A _8378_/B _8640_/A _8279_/C _8311_/B VGND VGND VPWR VPWR _8352_/A
+ sky130_fd_sc_hd__o32a_2
X_5556_ _5671_/A _5556_/B VGND VGND VPWR VPWR _5557_/A sky130_fd_sc_hd__or2_1
XFILLER_183_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8275_ _8275_/A _8693_/B VGND VGND VPWR VPWR _8275_/X sky130_fd_sc_hd__or2_2
XFILLER_105_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4507_ _9777_/Q _4506_/A _5963_/B1 _4506_/Y VGND VGND VPWR VPWR _9777_/D sky130_fd_sc_hd__a22o_1
X_5487_ _9385_/Q _5482_/A _5967_/B1 _5482_/Y VGND VGND VPWR VPWR _9385_/D sky130_fd_sc_hd__a22o_1
X_7226_ _6298_/Y _7048_/B _6297_/Y _7077_/A _7225_/X VGND VGND VPWR VPWR _7233_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_132_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7157_ _6664_/Y _7077_/C _6693_/Y _7077_/D _7156_/X VGND VGND VPWR VPWR _7157_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_86_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6108_ _6103_/Y _5431_/B _6104_/Y _6027_/B _6107_/X VGND VGND VPWR VPWR _6119_/B
+ sky130_fd_sc_hd__o221a_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7088_ _7088_/A VGND VGND VPWR VPWR _7088_/X sky130_fd_sc_hd__buf_8
XFILLER_132_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9729_ _9774_/CLK _9729_/D _9757_/SET_B VGND VGND VPWR VPWR _9729_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_19 _7644_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6390_ _9472_/Q VGND VGND VPWR VPWR _6390_/Y sky130_fd_sc_hd__clkinv_4
X_5410_ _9438_/Q _5406_/A _5966_/B1 _5406_/Y VGND VGND VPWR VPWR _9438_/D sky130_fd_sc_hd__a22o_1
XFILLER_161_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5341_ _9486_/Q _5338_/A _5965_/B1 _5338_/Y VGND VGND VPWR VPWR _9486_/D sky130_fd_sc_hd__a22o_1
X_8060_ _8060_/A VGND VGND VPWR VPWR _8061_/C sky130_fd_sc_hd__inv_2
X_5272_ _9533_/Q _5269_/A _8844_/X _5269_/Y VGND VGND VPWR VPWR _9533_/D sky130_fd_sc_hd__a22o_1
XFILLER_99_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7011_ _9586_/Q _7011_/B VGND VGND VPWR VPWR _7011_/Y sky130_fd_sc_hd__nor2_1
XFILLER_141_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8962_ _7739_/X _8962_/A1 _8975_/S VGND VGND VPWR VPWR _8962_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7913_ _8077_/A _8246_/B _7864_/X _8316_/A _7912_/X VGND VGND VPWR VPWR _7917_/B
+ sky130_fd_sc_hd__o221ai_1
X_8893_ _8892_/X _9147_/Q _9054_/Q VGND VGND VPWR VPWR _8893_/X sky130_fd_sc_hd__mux2_1
X_7844_ _8394_/A _8379_/B _8394_/C _8195_/A VGND VGND VPWR VPWR _7845_/A sky130_fd_sc_hd__or4_1
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7775_ _8193_/A _7775_/B _7775_/C _7775_/D VGND VGND VPWR VPWR _7966_/C sky130_fd_sc_hd__or4_1
XFILLER_178_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9514_ _9514_/CLK _9514_/D _4628_/A VGND VGND VPWR VPWR _9514_/Q sky130_fd_sc_hd__dfrtp_1
X_6726_ _6726_/A VGND VGND VPWR VPWR _6726_/Y sky130_fd_sc_hd__clkinv_2
X_4987_ _4987_/A VGND VGND VPWR VPWR _4987_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_149_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6657_ _9434_/Q VGND VGND VPWR VPWR _6657_/Y sky130_fd_sc_hd__inv_2
X_9445_ _9791_/CLK _9445_/D _9633_/SET_B VGND VGND VPWR VPWR _9445_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_191_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6588_ _9505_/Q VGND VGND VPWR VPWR _8777_/A sky130_fd_sc_hd__inv_6
XFILLER_164_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5608_ _9303_/Q _5604_/A _5966_/B1 _5604_/Y VGND VGND VPWR VPWR _9303_/D sky130_fd_sc_hd__a22o_1
X_9376_ _9379_/CLK _9376_/D _9779_/SET_B VGND VGND VPWR VPWR _9376_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_145_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5539_ _9351_/Q _5536_/A _8844_/X _5536_/Y VGND VGND VPWR VPWR _9351_/D sky130_fd_sc_hd__a22o_1
XFILLER_105_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8327_ _8327_/A _8599_/C _8506_/C _8693_/C VGND VGND VPWR VPWR _8327_/Y sky130_fd_sc_hd__nor4_2
XFILLER_3_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8258_ _8510_/A _8262_/B VGND VGND VPWR VPWR _8367_/B sky130_fd_sc_hd__nor2_1
X_8189_ _8189_/A _8213_/A VGND VGND VPWR VPWR _8189_/Y sky130_fd_sc_hd__nor2_1
XFILLER_160_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7209_ _6372_/Y _7068_/A _6402_/Y _7105_/X VGND VGND VPWR VPWR _7209_/X sky130_fd_sc_hd__o22a_1
XFILLER_143_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput17 mask_rev_in[21] VGND VGND VPWR VPWR _6262_/A sky130_fd_sc_hd__clkbuf_1
Xinput28 mask_rev_in[31] VGND VGND VPWR VPWR _6106_/A sky130_fd_sc_hd__clkbuf_1
Xinput39 mgmt_gpio_in[12] VGND VGND VPWR VPWR _6455_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_143_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4910_ _9520_/Q VGND VGND VPWR VPWR _4910_/Y sky130_fd_sc_hd__inv_4
XFILLER_92_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5890_ _5849_/A _8883_/X _8924_/X _9143_/Q VGND VGND VPWR VPWR _9143_/D sky130_fd_sc_hd__o22a_1
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4841_ _6111_/A _4900_/B VGND VGND VPWR VPWR _4841_/X sky130_fd_sc_hd__or2_4
XFILLER_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7560_ _6275_/Y _7434_/X _6240_/Y _7436_/X VGND VGND VPWR VPWR _7560_/X sky130_fd_sc_hd__o22a_1
X_4772_ _4787_/A _6086_/B VGND VGND VPWR VPWR _5583_/B sky130_fd_sc_hd__or2_4
XFILLER_20_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7491_ _6855_/Y _7445_/X _6871_/Y _7447_/X VGND VGND VPWR VPWR _7491_/X sky130_fd_sc_hd__o22a_1
X_6511_ _9221_/Q VGND VGND VPWR VPWR _8753_/A sky130_fd_sc_hd__inv_6
XFILLER_9_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6442_ _6440_/Y _5526_/B _6441_/Y _5897_/B VGND VGND VPWR VPWR _6442_/X sky130_fd_sc_hd__o22a_1
X_9230_ _9440_/CLK _9230_/D _9685_/SET_B VGND VGND VPWR VPWR _9230_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_173_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9161_ _9532_/CLK _9161_/D _9528_/SET_B VGND VGND VPWR VPWR _9161_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_161_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8112_ _8640_/B VGND VGND VPWR VPWR _8390_/B sky130_fd_sc_hd__inv_4
Xclkbuf_3_0_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A VGND VGND VPWR VPWR _9203_/CLK sky130_fd_sc_hd__clkbuf_2
X_6373_ _9216_/Q VGND VGND VPWR VPWR _6373_/Y sky130_fd_sc_hd__clkinv_2
X_5324_ _9497_/Q _5319_/A _8929_/A1 _5319_/Y VGND VGND VPWR VPWR _9497_/D sky130_fd_sc_hd__a22o_1
XFILLER_114_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9092_ _8837_/A1 _9092_/D _5980_/X VGND VGND VPWR VPWR _9092_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_114_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8043_ _8097_/B _8552_/A _8042_/X VGND VGND VPWR VPWR _8045_/A sky130_fd_sc_hd__o21ai_1
X_5255_ _9544_/Q _5253_/A _5964_/B1 _5253_/Y VGND VGND VPWR VPWR _9544_/D sky130_fd_sc_hd__a22o_1
X_5186_ _9588_/Q _5180_/A _8916_/A1 _5180_/Y VGND VGND VPWR VPWR _9588_/D sky130_fd_sc_hd__a22o_1
XFILLER_113_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8945_ _9083_/Q _9082_/Q _9051_/Q VGND VGND VPWR VPWR _8945_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8876_ _7177_/Y _9634_/Q _8959_/S VGND VGND VPWR VPWR _8876_/X sky130_fd_sc_hd__mux2_1
X_7827_ _8175_/A VGND VGND VPWR VPWR _8476_/A sky130_fd_sc_hd__inv_2
XFILLER_51_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7758_ _8660_/C VGND VGND VPWR VPWR _8282_/C sky130_fd_sc_hd__clkinv_2
XFILLER_8_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6709_ _6704_/Y _5355_/B _6705_/Y _5336_/B _6708_/X VGND VGND VPWR VPWR _6716_/C
+ sky130_fd_sc_hd__o221a_1
X_7689_ _6409_/Y _7445_/X _6404_/Y _7447_/X VGND VGND VPWR VPWR _7689_/X sky130_fd_sc_hd__o22a_1
XFILLER_11_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9428_ _9508_/CLK _9428_/D _9647_/SET_B VGND VGND VPWR VPWR _9428_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_138_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9359_ _9493_/CLK _9359_/D _4628_/A VGND VGND VPWR VPWR _9359_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_105_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _8973_/X _4551_/B _9679_/Q _5062_/D VGND VGND VPWR VPWR _9679_/D sky130_fd_sc_hd__a22o_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6991_ _9791_/Q VGND VGND VPWR VPWR _6991_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8730_ _8730_/A _8730_/B _8730_/C _8730_/D VGND VGND VPWR VPWR _8731_/B sky130_fd_sc_hd__or4_2
X_5942_ _5942_/A VGND VGND VPWR VPWR _5943_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_65_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8661_ _8660_/C _8341_/A _8660_/B _8660_/X _8556_/Y VGND VGND VPWR VPWR _8661_/X
+ sky130_fd_sc_hd__o311a_1
X_5873_ _5873_/A VGND VGND VPWR VPWR _5874_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_21_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8592_ _8592_/A VGND VGND VPWR VPWR _8641_/A sky130_fd_sc_hd__inv_2
X_7612_ _4712_/Y _7415_/X _4784_/Y _7417_/X _7611_/X VGND VGND VPWR VPWR _7626_/B
+ sky130_fd_sc_hd__o221a_1
X_4824_ _6111_/A _4891_/A VGND VGND VPWR VPWR _5100_/B sky130_fd_sc_hd__or2_4
XFILLER_138_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4755_ _4787_/A _4931_/A VGND VGND VPWR VPWR _4756_/A sky130_fd_sc_hd__or2_1
X_7543_ _6337_/Y _7430_/X _6402_/Y _7432_/X _7542_/X VGND VGND VPWR VPWR _7543_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_146_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4686_ _4921_/A _4780_/B VGND VGND VPWR VPWR _5810_/B sky130_fd_sc_hd__or2_4
X_7474_ _7476_/A _9251_/Q _7474_/C _7474_/D VGND VGND VPWR VPWR _7475_/A sky130_fd_sc_hd__or4_1
X_9213_ _9758_/CLK _9213_/D _9779_/SET_B VGND VGND VPWR VPWR _9213_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6425_ _6423_/Y _5450_/B _6424_/Y _5518_/B VGND VGND VPWR VPWR _6425_/X sky130_fd_sc_hd__o22a_1
X_6356_ _9290_/Q VGND VGND VPWR VPWR _6356_/Y sky130_fd_sc_hd__inv_2
XFILLER_161_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9144_ _9279_/CLK _9144_/D _9633_/SET_B VGND VGND VPWR VPWR _9144_/Q sky130_fd_sc_hd__dfrtp_1
X_5307_ _5307_/A VGND VGND VPWR VPWR _5308_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_161_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9075_ _9358_/CLK _9075_/D _9685_/SET_B VGND VGND VPWR VPWR _9075_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6287_ _9343_/Q VGND VGND VPWR VPWR _6287_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8026_ _8097_/B _8130_/B _8023_/X _8407_/A _8454_/B VGND VGND VPWR VPWR _8026_/X
+ sky130_fd_sc_hd__o2111a_1
X_5238_ _9555_/Q _5234_/A _5966_/B1 _5234_/Y VGND VGND VPWR VPWR _9555_/D sky130_fd_sc_hd__a22o_1
XFILLER_29_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5169_ _5169_/A VGND VGND VPWR VPWR _5169_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8928_ _9615_/Q _8844_/X _8930_/S VGND VGND VPWR VPWR _8928_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8859_ _8858_/X _9168_/Q _9054_/Q VGND VGND VPWR VPWR _8859_/X sky130_fd_sc_hd__mux2_1
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4540_ _5966_/B1 _9760_/Q _4540_/S VGND VGND VPWR VPWR _4541_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4471_ _4471_/A VGND VGND VPWR VPWR _4787_/A sky130_fd_sc_hd__buf_8
XFILLER_171_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7190_ _8763_/A _7112_/X _7699_/A _7077_/B VGND VGND VPWR VPWR _7190_/X sky130_fd_sc_hd__o22a_1
X_6210_ _6205_/Y _5507_/B _6206_/Y _6086_/X _6209_/X VGND VGND VPWR VPWR _6211_/D
+ sky130_fd_sc_hd__o221a_2
XFILLER_131_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6141_ _9327_/Q VGND VGND VPWR VPWR _6141_/Y sky130_fd_sc_hd__inv_2
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6072_ _9449_/Q VGND VGND VPWR VPWR _6072_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5023_ _9688_/Q _5015_/A _8916_/A1 _5015_/Y VGND VGND VPWR VPWR _9688_/D sky130_fd_sc_hd__a22o_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6974_ _6974_/A _6974_/B VGND VGND VPWR VPWR _6975_/A sky130_fd_sc_hd__or2_1
X_9762_ _9770_/CLK _9762_/D _7011_/B VGND VGND VPWR VPWR _9762_/Q sky130_fd_sc_hd__dfrtp_4
X_5925_ _7768_/C _7768_/D _5925_/C input149/X VGND VGND VPWR VPWR _5936_/A sky130_fd_sc_hd__or4b_1
X_8713_ _8713_/A _8713_/B _8713_/C _8713_/D VGND VGND VPWR VPWR _8714_/B sky130_fd_sc_hd__or4_1
XFILLER_110_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9693_ _9695_/CLK _9693_/D _9779_/SET_B VGND VGND VPWR VPWR _9693_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_110_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8644_ _8677_/D _8719_/C _8731_/A _8675_/D VGND VGND VPWR VPWR _8647_/A sky130_fd_sc_hd__or4_4
X_5856_ _5849_/X _8861_/X _8924_/X _9170_/Q VGND VGND VPWR VPWR _9170_/D sky130_fd_sc_hd__o22a_1
XFILLER_21_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4807_ _4807_/A VGND VGND VPWR VPWR _4808_/A sky130_fd_sc_hd__buf_2
X_8575_ _8575_/A _8575_/B _8575_/C VGND VGND VPWR VPWR _8576_/D sky130_fd_sc_hd__or3_1
X_5787_ _5787_/A VGND VGND VPWR VPWR _5787_/Y sky130_fd_sc_hd__inv_2
X_4738_ _4787_/A _4927_/A VGND VGND VPWR VPWR _4739_/A sky130_fd_sc_hd__or2_1
X_7526_ _7703_/A _7425_/X _7523_/X _7525_/X VGND VGND VPWR VPWR _7536_/C sky130_fd_sc_hd__o211a_1
XFILLER_21_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7457_ _7457_/A VGND VGND VPWR VPWR _7457_/X sky130_fd_sc_hd__buf_8
X_4669_ _4669_/A _4729_/D _8946_/X _8944_/X VGND VGND VPWR VPWR _4927_/A sky130_fd_sc_hd__or4_4
XFILLER_162_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6408_ _6408_/A _6408_/B _6408_/C _6408_/D VGND VGND VPWR VPWR _6474_/A sky130_fd_sc_hd__and4_1
XFILLER_122_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7388_ _6361_/Y _7112_/X _6441_/Y _7077_/B VGND VGND VPWR VPWR _7388_/X sky130_fd_sc_hd__o22a_1
X_9127_ _9379_/CLK _9127_/D _9646_/SET_B VGND VGND VPWR VPWR _9127_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6339_ _6334_/Y _5968_/B _6335_/Y _5488_/B _6338_/X VGND VGND VPWR VPWR _6352_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_76_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9058_ _9058_/CLK _9058_/D _6041_/X VGND VGND VPWR VPWR _9058_/Q sky130_fd_sc_hd__dfstp_1
X_8009_ _8009_/A _8060_/A VGND VGND VPWR VPWR _8009_/X sky130_fd_sc_hd__or2_1
XFILLER_130_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5710_ _7472_/A VGND VGND VPWR VPWR _5710_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6690_ _6690_/A _6690_/B _6690_/C _6690_/D VGND VGND VPWR VPWR _6691_/D sky130_fd_sc_hd__and4_1
XFILLER_31_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5641_ _9277_/Q VGND VGND VPWR VPWR _5647_/A sky130_fd_sc_hd__inv_2
XFILLER_31_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5572_ _6052_/A _5572_/B VGND VGND VPWR VPWR _5573_/A sky130_fd_sc_hd__or2_1
X_8360_ _8360_/A _8573_/C _8642_/C _8574_/C VGND VGND VPWR VPWR _8364_/A sky130_fd_sc_hd__or4_1
XFILLER_191_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8291_ _8672_/C _8650_/B _8291_/C VGND VGND VPWR VPWR _8292_/B sky130_fd_sc_hd__or3_1
XFILLER_144_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7311_ _6927_/Y _7077_/C _6904_/Y _7077_/D _7310_/X VGND VGND VPWR VPWR _7311_/X
+ sky130_fd_sc_hd__o221a_1
Xclkbuf_1_0_1_csclk clkbuf_1_0_1_csclk/A VGND VGND VPWR VPWR clkbuf_2_1_0_csclk/A
+ sky130_fd_sc_hd__clkbuf_2
X_4523_ _6111_/A _6111_/B VGND VGND VPWR VPWR _4524_/B sky130_fd_sc_hd__or2_4
X_7242_ _7242_/A _7242_/B _7242_/C _7242_/D VGND VGND VPWR VPWR _7243_/C sky130_fd_sc_hd__and4_1
X_4454_ _6052_/A VGND VGND VPWR VPWR _5960_/A sky130_fd_sc_hd__buf_12
XFILLER_131_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7173_ _6763_/Y _5728_/X _6673_/Y _7040_/A _7172_/X VGND VGND VPWR VPWR _7176_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_98_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6124_ _6122_/Y _5757_/B _6123_/Y _5905_/B VGND VGND VPWR VPWR _6124_/X sky130_fd_sc_hd__o22a_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6055_ _9047_/Q _6054_/A _8929_/A1 _6054_/Y VGND VGND VPWR VPWR _9047_/D sky130_fd_sc_hd__a22o_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5006_ _5006_/A VGND VGND VPWR VPWR _5007_/S sky130_fd_sc_hd__clkbuf_1
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_109 input86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6957_ _6629_/Y _6952_/A _9031_/Q _6952_/Y VGND VGND VPWR VPWR _9031_/D sky130_fd_sc_hd__o22a_1
XFILLER_121_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9745_ _9777_/CLK _9745_/D _9757_/SET_B VGND VGND VPWR VPWR _9745_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_41_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5908_ _9132_/Q _5907_/A _8846_/X _5907_/Y VGND VGND VPWR VPWR _9132_/D sky130_fd_sc_hd__a22o_1
X_6888_ _6883_/Y _5829_/B _6884_/Y _5583_/B _6887_/X VGND VGND VPWR VPWR _6901_/B
+ sky130_fd_sc_hd__o221a_1
X_9676_ _9681_/CLK _9676_/D _6146_/A VGND VGND VPWR VPWR _9676_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_139_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5839_ _5839_/A VGND VGND VPWR VPWR _5839_/Y sky130_fd_sc_hd__inv_2
X_8627_ _8627_/A _8627_/B _8627_/C _8627_/D VGND VGND VPWR VPWR _8686_/D sky130_fd_sc_hd__or4_2
XFILLER_14_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8558_ _8558_/A VGND VGND VPWR VPWR _8688_/B sky130_fd_sc_hd__inv_2
XFILLER_147_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7509_ _6710_/Y _7445_/X _6767_/Y _7447_/X VGND VGND VPWR VPWR _7509_/X sky130_fd_sc_hd__o22a_1
XFILLER_135_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8489_ _8720_/A _8713_/A _8703_/A VGND VGND VPWR VPWR _8603_/A sky130_fd_sc_hd__or3_1
XFILLER_162_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput308 _8822_/X VGND VGND VPWR VPWR serial_data_1 sky130_fd_sc_hd__buf_2
XFILLER_99_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput319 _9764_/Q VGND VGND VPWR VPWR sram_ro_addr[2] sky130_fd_sc_hd__buf_2
XFILLER_141_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7860_ _8515_/B _8262_/B VGND VGND VPWR VPWR _8667_/A sky130_fd_sc_hd__nor2_1
XFILLER_63_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6811_ _9722_/Q VGND VGND VPWR VPWR _6811_/Y sky130_fd_sc_hd__inv_2
X_7791_ _8189_/A _7791_/B VGND VGND VPWR VPWR _7792_/B sky130_fd_sc_hd__nor2_1
XFILLER_50_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9530_ _9532_/CLK _9530_/D _9647_/SET_B VGND VGND VPWR VPWR _9530_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6742_ _9634_/Q VGND VGND VPWR VPWR _6742_/Y sky130_fd_sc_hd__inv_2
X_6673_ _9095_/Q VGND VGND VPWR VPWR _6673_/Y sky130_fd_sc_hd__clkinv_2
X_9461_ _9789_/CLK _9461_/D _9647_/SET_B VGND VGND VPWR VPWR _9461_/Q sky130_fd_sc_hd__dfrtp_1
X_9392_ _9483_/CLK _9392_/D _9528_/SET_B VGND VGND VPWR VPWR _9392_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_176_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5624_ _9293_/Q _5623_/A _8846_/X _5623_/Y VGND VGND VPWR VPWR _9293_/D sky130_fd_sc_hd__a22o_1
X_8412_ _8550_/A _8401_/B _8409_/X _8411_/Y VGND VGND VPWR VPWR _8412_/X sky130_fd_sc_hd__o211a_1
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8343_ _7886_/B _8003_/Y _8110_/C VGND VGND VPWR VPWR _8343_/Y sky130_fd_sc_hd__o21ai_2
X_5555_ _9338_/Q _5547_/A _8839_/X _5547_/Y VGND VGND VPWR VPWR _9338_/D sky130_fd_sc_hd__a22o_1
XFILLER_129_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8274_ _8510_/A _8660_/B _8496_/A VGND VGND VPWR VPWR _8693_/B sky130_fd_sc_hd__nor3_1
X_4506_ _4506_/A VGND VGND VPWR VPWR _4506_/Y sky130_fd_sc_hd__inv_2
X_5486_ _9386_/Q _5482_/A _5966_/B1 _5482_/Y VGND VGND VPWR VPWR _9386_/D sky130_fd_sc_hd__a22o_1
X_7225_ _6282_/Y _7040_/C _6304_/Y _7059_/C VGND VGND VPWR VPWR _7225_/X sky130_fd_sc_hd__o22a_1
X_7156_ _6713_/Y _7086_/X _6710_/Y _7088_/X VGND VGND VPWR VPWR _7156_/X sky130_fd_sc_hd__o22a_1
XFILLER_86_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6107_ _6105_/Y _5110_/B _6106_/Y _4822_/X VGND VGND VPWR VPWR _6107_/X sky130_fd_sc_hd__o22a_4
XFILLER_100_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7087_ _7127_/C _7087_/B VGND VGND VPWR VPWR _7088_/A sky130_fd_sc_hd__or2_1
X_6038_ _9069_/Q _4466_/A _8929_/A1 _4466_/Y VGND VGND VPWR VPWR _9069_/D sky130_fd_sc_hd__a22o_1
XFILLER_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7989_ _8098_/A _8386_/B VGND VGND VPWR VPWR _8050_/B sky130_fd_sc_hd__or2_1
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9728_ _9769_/CLK _9728_/D _7011_/B VGND VGND VPWR VPWR _9728_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9659_ _4450_/A1 _9659_/D _6146_/A VGND VGND VPWR VPWR _9659_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_17_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR _9508_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_32_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5340_ _9487_/Q _5338_/A _5964_/B1 _5338_/Y VGND VGND VPWR VPWR _9487_/D sky130_fd_sc_hd__a22o_1
X_5271_ _9534_/Q _5269_/A _8845_/X _5269_/Y VGND VGND VPWR VPWR _9534_/D sky130_fd_sc_hd__a22o_1
XFILLER_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7010_ _9626_/Q _7011_/B VGND VGND VPWR VPWR _7010_/Y sky130_fd_sc_hd__nor2_1
XFILLER_68_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8961_ _7737_/X _8961_/A1 _8975_/S VGND VGND VPWR VPWR _8961_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7912_ _8238_/A _7864_/X _7909_/X _7910_/X _8454_/A VGND VGND VPWR VPWR _7912_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_83_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8892_ _7353_/Y _9629_/Q _8959_/S VGND VGND VPWR VPWR _8892_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7843_ _8515_/B _7848_/A VGND VGND VPWR VPWR _7931_/A sky130_fd_sc_hd__or2_2
XFILLER_63_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7774_ _7959_/A _8583_/A _7774_/C _7774_/D VGND VGND VPWR VPWR _7775_/D sky130_fd_sc_hd__nand4bb_1
X_4986_ _4994_/A VGND VGND VPWR VPWR _4987_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_51_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9513_ _9514_/CLK _9513_/D _4628_/A VGND VGND VPWR VPWR _9513_/Q sky130_fd_sc_hd__dfrtp_1
X_6725_ _9556_/Q VGND VGND VPWR VPWR _6725_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_164_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6656_ _9764_/Q VGND VGND VPWR VPWR _6656_/Y sky130_fd_sc_hd__inv_2
X_9444_ _9785_/CLK _9444_/D _9779_/SET_B VGND VGND VPWR VPWR _9444_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_191_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5607_ _9304_/Q _5604_/A _5965_/B1 _5604_/Y VGND VGND VPWR VPWR _9304_/D sky130_fd_sc_hd__a22o_1
X_9375_ _9379_/CLK _9375_/D _9779_/SET_B VGND VGND VPWR VPWR _9375_/Q sky130_fd_sc_hd__dfrtp_4
X_6587_ _9388_/Q VGND VGND VPWR VPWR _6587_/Y sky130_fd_sc_hd__inv_2
X_5538_ _9352_/Q _5536_/A _8845_/X _5536_/Y VGND VGND VPWR VPWR _9352_/D sky130_fd_sc_hd__a22o_1
X_8326_ _8468_/A _8715_/B VGND VGND VPWR VPWR _8693_/C sky130_fd_sc_hd__or2_1
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8257_ _8257_/A _8674_/B VGND VGND VPWR VPWR _8259_/A sky130_fd_sc_hd__or2_1
X_5469_ _5545_/A _6081_/B VGND VGND VPWR VPWR _5470_/A sky130_fd_sc_hd__or2_1
X_7208_ _6356_/Y _7059_/B _6392_/Y _7068_/C _7207_/X VGND VGND VPWR VPWR _7211_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_105_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8188_ _8305_/A _8188_/B VGND VGND VPWR VPWR _8606_/B sky130_fd_sc_hd__nor2_2
XFILLER_132_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7139_ _6854_/Y _7097_/X _6832_/Y _7099_/X VGND VGND VPWR VPWR _7139_/X sky130_fd_sc_hd__o22a_1
XFILLER_100_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput18 mask_rev_in[22] VGND VGND VPWR VPWR _6208_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_155_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput29 mask_rev_in[3] VGND VGND VPWR VPWR _6618_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_155_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4840_ _4840_/A VGND VGND VPWR VPWR _4840_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4771_ _9312_/Q VGND VGND VPWR VPWR _4771_/Y sky130_fd_sc_hd__inv_2
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6510_ _9267_/Q VGND VGND VPWR VPWR _6510_/Y sky130_fd_sc_hd__inv_2
XFILLER_146_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7490_ _6919_/Y _7425_/X _7487_/X _7489_/X VGND VGND VPWR VPWR _7500_/C sky130_fd_sc_hd__o211a_1
XFILLER_146_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6441_ _9137_/Q VGND VGND VPWR VPWR _6441_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_173_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9160_ _9358_/CLK _9160_/D _9528_/SET_B VGND VGND VPWR VPWR _9160_/Q sky130_fd_sc_hd__dfrtp_1
X_6372_ _9222_/Q VGND VGND VPWR VPWR _6372_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_161_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5323_ _9498_/Q _5319_/A _8925_/A1 _5319_/Y VGND VGND VPWR VPWR _9498_/D sky130_fd_sc_hd__a22o_1
X_8111_ _8378_/B VGND VGND VPWR VPWR _8544_/B sky130_fd_sc_hd__clkinv_4
XFILLER_114_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9091_ _8837_/A1 _9091_/D _5984_/X VGND VGND VPWR VPWR _9091_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_142_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8042_ _8389_/A _8552_/A _8041_/Y VGND VGND VPWR VPWR _8042_/X sky130_fd_sc_hd__o21a_1
X_5254_ _9545_/Q _5253_/A _5963_/B1 _5253_/Y VGND VGND VPWR VPWR _9545_/D sky130_fd_sc_hd__a22o_1
X_5185_ _9589_/Q _5180_/A _8840_/X _5180_/Y VGND VGND VPWR VPWR _9589_/D sky130_fd_sc_hd__a22o_1
XFILLER_110_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8944_ _8943_/X _9675_/Q _9587_/Q VGND VGND VPWR VPWR _8944_/X sky130_fd_sc_hd__mux2_4
XFILLER_56_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8875_ _8874_/X _9138_/Q _9054_/Q VGND VGND VPWR VPWR _8875_/X sky130_fd_sc_hd__mux2_1
XFILLER_169_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7826_ _8515_/A _8272_/A VGND VGND VPWR VPWR _8175_/A sky130_fd_sc_hd__or2_1
XFILLER_24_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7757_ _7757_/A VGND VGND VPWR VPWR _8660_/C sky130_fd_sc_hd__buf_4
X_4969_ _4969_/A VGND VGND VPWR VPWR _4969_/X sky130_fd_sc_hd__clkbuf_1
X_6708_ _6706_/Y _4870_/X _6707_/Y _5602_/B VGND VGND VPWR VPWR _6708_/X sky130_fd_sc_hd__o22a_1
X_7688_ _6458_/Y _7425_/X _7685_/X _7687_/X VGND VGND VPWR VPWR _7698_/C sky130_fd_sc_hd__o211a_1
X_9427_ _9527_/CLK _9427_/D _9528_/SET_B VGND VGND VPWR VPWR _9427_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_137_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6639_ _9220_/Q VGND VGND VPWR VPWR _6639_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_138_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9358_ _9358_/CLK _9358_/D _9685_/SET_B VGND VGND VPWR VPWR _9358_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9289_ _9596_/CLK _9289_/D _9528_/SET_B VGND VGND VPWR VPWR _9289_/Q sky130_fd_sc_hd__dfrtp_1
X_8309_ _7864_/X _8498_/A _8341_/B _8498_/B VGND VGND VPWR VPWR _8309_/X sky130_fd_sc_hd__o22a_1
XFILLER_105_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6990_ _9709_/Q _6023_/Y _4953_/Y _9049_/Q VGND VGND VPWR VPWR _9049_/D sky130_fd_sc_hd__a31o_1
XFILLER_92_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5941_ _5960_/A _5941_/B VGND VGND VPWR VPWR _5942_/A sky130_fd_sc_hd__or2_1
XFILLER_65_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8660_ _8660_/A _8660_/B _8660_/C VGND VGND VPWR VPWR _8660_/X sky130_fd_sc_hd__or3_1
X_5872_ _6052_/A _5872_/B VGND VGND VPWR VPWR _5873_/A sky130_fd_sc_hd__or2_1
XFILLER_61_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8591_ _8510_/A _8498_/A _7879_/B _8397_/A VGND VGND VPWR VPWR _8591_/Y sky130_fd_sc_hd__o211ai_1
X_4823_ _9641_/Q VGND VGND VPWR VPWR _4823_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7611_ _4677_/Y _7419_/X _4809_/Y _7421_/X VGND VGND VPWR VPWR _7611_/X sky130_fd_sc_hd__o22a_1
XFILLER_193_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4754_ _4754_/A VGND VGND VPWR VPWR _4754_/Y sky130_fd_sc_hd__inv_2
X_7542_ _6346_/Y _7434_/X _6329_/Y _7436_/X VGND VGND VPWR VPWR _7542_/X sky130_fd_sc_hd__o22a_1
XFILLER_146_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7473_ _7473_/A VGND VGND VPWR VPWR _7473_/X sky130_fd_sc_hd__buf_8
XFILLER_174_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4685_ _9198_/Q VGND VGND VPWR VPWR _4685_/Y sky130_fd_sc_hd__inv_2
X_9212_ _9655_/CLK _9212_/D _9779_/SET_B VGND VGND VPWR VPWR _9212_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_161_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6424_ _9363_/Q VGND VGND VPWR VPWR _6424_/Y sky130_fd_sc_hd__inv_2
X_9143_ _9203_/CLK _9143_/D _9633_/SET_B VGND VGND VPWR VPWR _9143_/Q sky130_fd_sc_hd__dfrtp_1
X_6355_ _6354_/Y _5121_/B _4844_/X _6158_/X VGND VGND VPWR VPWR _6355_/X sky130_fd_sc_hd__o211a_1
X_9074_ _9687_/CLK _9074_/D _9685_/SET_B VGND VGND VPWR VPWR _9074_/Q sky130_fd_sc_hd__dfrtp_1
X_5306_ _5545_/A _5306_/B VGND VGND VPWR VPWR _5307_/A sky130_fd_sc_hd__or2_1
X_6286_ _6281_/Y _6165_/A _6282_/Y _5045_/B _6285_/X VGND VGND VPWR VPWR _6307_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_130_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8025_ _8624_/B _8137_/B VGND VGND VPWR VPWR _8454_/B sky130_fd_sc_hd__or2_1
XFILLER_0_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5237_ _9556_/Q _5234_/A _5965_/B1 _5234_/Y VGND VGND VPWR VPWR _9556_/D sky130_fd_sc_hd__a22o_1
XFILLER_102_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5168_ _5168_/A VGND VGND VPWR VPWR _5169_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_68_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5099_ _9646_/Q _5091_/A _8916_/A1 _5091_/Y VGND VGND VPWR VPWR _9646_/D sky130_fd_sc_hd__a22o_1
XFILLER_44_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8927_ _9616_/Q _8845_/X _8930_/S VGND VGND VPWR VPWR _8927_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8858_ _7572_/Y _9637_/Q _8978_/S VGND VGND VPWR VPWR _8858_/X sky130_fd_sc_hd__mux2_1
X_8789_ _8789_/A VGND VGND VPWR VPWR _8790_/A sky130_fd_sc_hd__clkbuf_1
X_7809_ _7903_/C _8528_/A _8525_/A _8189_/A VGND VGND VPWR VPWR _7878_/A sky130_fd_sc_hd__or4_1
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4470_ _8936_/X _4665_/B _4801_/C VGND VGND VPWR VPWR _4471_/A sky130_fd_sc_hd__or3_1
XFILLER_143_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6140_ _9197_/Q VGND VGND VPWR VPWR _6140_/Y sky130_fd_sc_hd__inv_2
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6071_ _6071_/A _6071_/B VGND VGND VPWR VPWR _6071_/Y sky130_fd_sc_hd__nand2_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5022_ _9689_/Q _5015_/A _8930_/A1 _5015_/Y VGND VGND VPWR VPWR _9689_/D sky130_fd_sc_hd__a22o_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6973_ _9061_/Q VGND VGND VPWR VPWR _6974_/A sky130_fd_sc_hd__inv_2
X_9761_ _9770_/CLK _9761_/D _7011_/B VGND VGND VPWR VPWR _9761_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_53_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5924_ _9065_/D VGND VGND VPWR VPWR _6147_/B sky130_fd_sc_hd__inv_2
X_8712_ _8738_/A _8712_/B VGND VGND VPWR VPWR _8712_/Y sky130_fd_sc_hd__nor2_1
X_9692_ _9695_/CLK _9692_/D _9779_/SET_B VGND VGND VPWR VPWR _9692_/Q sky130_fd_sc_hd__dfrtp_1
X_8643_ _7987_/Y _8390_/B _8317_/B _8364_/D _8576_/D VGND VGND VPWR VPWR _8675_/D
+ sky130_fd_sc_hd__a2111o_2
X_5855_ _5849_/X _8863_/X _8924_/X _9171_/Q VGND VGND VPWR VPWR _9171_/D sky130_fd_sc_hd__o22a_1
X_4806_ _9770_/Q _9708_/Q _9626_/Q VGND VGND VPWR VPWR _4807_/A sky130_fd_sc_hd__or3_1
XFILLER_119_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5786_ _9218_/Q _5778_/A _8916_/A1 _5778_/Y VGND VGND VPWR VPWR _9218_/D sky130_fd_sc_hd__a22o_1
X_8574_ _8574_/A _8574_/B _8574_/C VGND VGND VPWR VPWR _8730_/D sky130_fd_sc_hd__or3_1
X_4737_ _4737_/A VGND VGND VPWR VPWR _4737_/Y sky130_fd_sc_hd__clkinv_2
X_7525_ _7701_/A _7430_/X _8785_/A _7432_/X _7524_/X VGND VGND VPWR VPWR _7525_/X
+ sky130_fd_sc_hd__o221a_1
X_4668_ _9151_/Q VGND VGND VPWR VPWR _4668_/Y sky130_fd_sc_hd__inv_2
X_7456_ _7456_/A _7466_/A _9255_/Q VGND VGND VPWR VPWR _7457_/A sky130_fd_sc_hd__or3_1
XFILLER_162_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6407_ _6402_/Y _5240_/B _6403_/Y _4491_/B _6406_/X VGND VGND VPWR VPWR _6408_/D
+ sky130_fd_sc_hd__o221a_1
X_7387_ _7387_/A _7387_/B _7387_/C _7387_/D VGND VGND VPWR VPWR _7397_/B sky130_fd_sc_hd__and4_1
X_9126_ _9129_/CLK _9126_/D _9779_/SET_B VGND VGND VPWR VPWR _9126_/Q sky130_fd_sc_hd__dfstp_1
X_4599_ _9733_/Q _4592_/A _5966_/B1 _4592_/Y VGND VGND VPWR VPWR _9733_/D sky130_fd_sc_hd__a22o_1
X_6338_ _6336_/Y _4893_/X _6337_/Y _5905_/B VGND VGND VPWR VPWR _6338_/X sky130_fd_sc_hd__o22a_1
XFILLER_135_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9057_ _9280_/CLK _9057_/D _9757_/SET_B VGND VGND VPWR VPWR _9057_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6269_ _9403_/Q VGND VGND VPWR VPWR _6269_/Y sky130_fd_sc_hd__clkinv_4
X_8008_ _8218_/A _8218_/B _8008_/C VGND VGND VPWR VPWR _8060_/A sky130_fd_sc_hd__or3_4
Xclkbuf_2_3_0_csclk clkbuf_2_3_0_csclk/A VGND VGND VPWR VPWR clkbuf_2_3_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_91_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5640_ _9279_/Q VGND VGND VPWR VPWR _5649_/B sky130_fd_sc_hd__inv_2
XFILLER_129_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5571_ _9328_/Q _5566_/A _5967_/B1 _5566_/Y VGND VGND VPWR VPWR _9328_/D sky130_fd_sc_hd__a22o_1
XFILLER_184_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8290_ _8606_/B _8290_/B VGND VGND VPWR VPWR _8291_/C sky130_fd_sc_hd__or2_1
XFILLER_129_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7310_ _6873_/Y _7086_/X _6867_/Y _7088_/X VGND VGND VPWR VPWR _7310_/X sky130_fd_sc_hd__o22a_1
X_4522_ _8946_/X _4729_/B _8934_/X _4729_/D VGND VGND VPWR VPWR _6111_/B sky130_fd_sc_hd__or4_4
XFILLER_156_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7241_ _6269_/Y _7124_/X _6311_/Y _7068_/B _7240_/X VGND VGND VPWR VPWR _7242_/D
+ sky130_fd_sc_hd__o221a_1
X_4453_ _5133_/A VGND VGND VPWR VPWR _6052_/A sky130_fd_sc_hd__buf_12
XFILLER_7_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7172_ _7172_/A _7392_/B VGND VGND VPWR VPWR _7172_/X sky130_fd_sc_hd__or2_1
X_6123_ _9132_/Q VGND VGND VPWR VPWR _6123_/Y sky130_fd_sc_hd__inv_2
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6054_ _6054_/A VGND VGND VPWR VPWR _6054_/Y sky130_fd_sc_hd__inv_2
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5005_ _9091_/Q _6022_/C _9092_/Q _6022_/B VGND VGND VPWR VPWR _5006_/A sky130_fd_sc_hd__or4_1
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6956_ _6475_/Y _6952_/A _9032_/Q _6952_/Y VGND VGND VPWR VPWR _9032_/D sky130_fd_sc_hd__o22a_2
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9744_ _9777_/CLK _9744_/D _9757_/SET_B VGND VGND VPWR VPWR _9744_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_53_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5907_ _5907_/A VGND VGND VPWR VPWR _5907_/Y sky130_fd_sc_hd__inv_2
XFILLER_179_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9675_ _9681_/CLK _9675_/D _6146_/A VGND VGND VPWR VPWR _9675_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6887_ _6885_/Y _5564_/B _6886_/Y _6052_/C VGND VGND VPWR VPWR _6887_/X sky130_fd_sc_hd__o22a_1
X_5838_ _5838_/A VGND VGND VPWR VPWR _5839_/A sky130_fd_sc_hd__clkbuf_4
X_8626_ _8401_/A _8624_/X _8117_/A _8625_/Y VGND VGND VPWR VPWR _8629_/B sky130_fd_sc_hd__o22ai_2
XFILLER_14_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8557_ _8386_/A _7971_/A _8389_/A _7829_/A _8556_/Y VGND VGND VPWR VPWR _8558_/A
+ sky130_fd_sc_hd__o311a_1
XFILLER_139_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5769_ _5769_/A VGND VGND VPWR VPWR _5770_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_108_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7508_ _6775_/Y _7425_/X _7505_/X _7507_/X VGND VGND VPWR VPWR _7518_/C sky130_fd_sc_hd__o211a_1
XFILLER_147_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8488_ _8488_/A VGND VGND VPWR VPWR _8488_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7439_ _4687_/Y _7425_/X _7428_/X _7438_/X VGND VGND VPWR VPWR _7481_/C sky130_fd_sc_hd__o211a_1
XFILLER_150_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9109_ _9379_/CLK _9109_/D _9779_/SET_B VGND VGND VPWR VPWR _9109_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput309 _8823_/X VGND VGND VPWR VPWR serial_data_2 sky130_fd_sc_hd__buf_2
XFILLER_141_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6810_ _6805_/Y _5232_/B _6806_/Y _4841_/X _6809_/X VGND VGND VPWR VPWR _6829_/A
+ sky130_fd_sc_hd__o221a_1
X_7790_ _8528_/B _7900_/A VGND VGND VPWR VPWR _8538_/C sky130_fd_sc_hd__nand2_1
XFILLER_149_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6741_ _6741_/A _6741_/B _6741_/C _6741_/D VGND VGND VPWR VPWR _6784_/B sky130_fd_sc_hd__and4_1
XFILLER_50_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9460_ _9532_/CLK _9460_/D _9647_/SET_B VGND VGND VPWR VPWR _9460_/Q sky130_fd_sc_hd__dfstp_1
X_6672_ _6667_/Y _5045_/B _6668_/Y _5488_/B _6671_/X VGND VGND VPWR VPWR _6690_/A
+ sky130_fd_sc_hd__o221a_1
X_9391_ _9483_/CLK _9391_/D _9528_/SET_B VGND VGND VPWR VPWR _9391_/Q sky130_fd_sc_hd__dfstp_1
X_5623_ _5623_/A VGND VGND VPWR VPWR _5623_/Y sky130_fd_sc_hd__inv_2
X_8411_ _8734_/B _8574_/A VGND VGND VPWR VPWR _8411_/Y sky130_fd_sc_hd__nor2_1
XFILLER_117_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8342_ _8114_/Y _8115_/Y _8594_/B VGND VGND VPWR VPWR _8356_/A sky130_fd_sc_hd__a21o_1
X_5554_ _9339_/Q _5547_/A _8930_/A1 _5547_/Y VGND VGND VPWR VPWR _9339_/D sky130_fd_sc_hd__a22o_1
XFILLER_129_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8273_ _8273_/A _8715_/B VGND VGND VPWR VPWR _8275_/A sky130_fd_sc_hd__or2_1
XFILLER_105_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4505_ _4505_/A VGND VGND VPWR VPWR _4506_/A sky130_fd_sc_hd__clkbuf_2
X_5485_ _9387_/Q _5482_/A _5965_/B1 _5482_/Y VGND VGND VPWR VPWR _9387_/D sky130_fd_sc_hd__a22o_1
X_7224_ _6244_/Y _7082_/X _6256_/Y _7084_/X _7223_/X VGND VGND VPWR VPWR _7243_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_116_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7155_ _7155_/A _7155_/B _7155_/C VGND VGND VPWR VPWR _7155_/Y sky130_fd_sc_hd__nand3_4
X_6106_ _6106_/A VGND VGND VPWR VPWR _6106_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_112_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7086_ _7086_/A VGND VGND VPWR VPWR _7086_/X sky130_fd_sc_hd__buf_8
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6037_ _9070_/Q _6029_/A _8839_/X _6029_/Y VGND VGND VPWR VPWR _9070_/D sky130_fd_sc_hd__a22o_1
XFILLER_86_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7988_ _7988_/A _8091_/B VGND VGND VPWR VPWR _8386_/B sky130_fd_sc_hd__or2b_2
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6939_ _9232_/Q VGND VGND VPWR VPWR _6939_/Y sky130_fd_sc_hd__clkinv_2
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9727_ _9769_/CLK _9727_/D _7011_/B VGND VGND VPWR VPWR _9727_/Q sky130_fd_sc_hd__dfstp_1
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9658_ _9779_/CLK _9658_/D _9779_/SET_B VGND VGND VPWR VPWR _9658_/Q sky130_fd_sc_hd__dfrtp_1
X_8609_ _8609_/A VGND VGND VPWR VPWR _8666_/C sky130_fd_sc_hd__inv_2
X_9589_ _9617_/CLK _9589_/D _9295_/SET_B VGND VGND VPWR VPWR _9589_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_0_csclk _8847_/X VGND VGND VPWR VPWR clkbuf_0_csclk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_135_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_1_0_1_csclk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5270_ _9535_/Q _5269_/A _8846_/X _5269_/Y VGND VGND VPWR VPWR _9535_/D sky130_fd_sc_hd__a22o_1
XFILLER_141_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8960_ _7735_/X _5060_/X _8960_/S VGND VGND VPWR VPWR _8960_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7911_ _8521_/B _8239_/B VGND VGND VPWR VPWR _8454_/A sky130_fd_sc_hd__or2_1
XFILLER_83_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8891_ _8890_/X _9146_/Q _9054_/Q VGND VGND VPWR VPWR _8891_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7842_ _8660_/B _8496_/A VGND VGND VPWR VPWR _7848_/A sky130_fd_sc_hd__or2_2
X_7773_ _8525_/A VGND VGND VPWR VPWR _8583_/A sky130_fd_sc_hd__inv_6
X_4985_ _9701_/Q _4966_/A _4949_/A _4966_/Y VGND VGND VPWR VPWR _9701_/D sky130_fd_sc_hd__a22o_1
XFILLER_23_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6724_ _9374_/Q VGND VGND VPWR VPWR _6724_/Y sky130_fd_sc_hd__clkinv_2
X_9512_ _9514_/CLK _9512_/D _4628_/A VGND VGND VPWR VPWR _9512_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_23_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9443_ _9791_/CLK _9443_/D _9779_/SET_B VGND VGND VPWR VPWR _9443_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_192_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6655_ _6650_/Y _6027_/B _6651_/Y _4602_/B _6654_/X VGND VGND VPWR VPWR _6691_/A
+ sky130_fd_sc_hd__o221a_1
X_5606_ _9305_/Q _5604_/A _5964_/B1 _5604_/Y VGND VGND VPWR VPWR _9305_/D sky130_fd_sc_hd__a22o_1
X_9374_ _9379_/CLK _9374_/D _9646_/SET_B VGND VGND VPWR VPWR _9374_/Q sky130_fd_sc_hd__dfrtp_1
X_6586_ _6586_/A _6586_/B _6586_/C VGND VGND VPWR VPWR _6628_/B sky130_fd_sc_hd__and3_1
X_5537_ _9353_/Q _5536_/A _8846_/X _5536_/Y VGND VGND VPWR VPWR _9353_/D sky130_fd_sc_hd__a22o_1
X_8325_ _8325_/A VGND VGND VPWR VPWR _8468_/A sky130_fd_sc_hd__inv_2
XFILLER_117_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8256_ _8260_/A _8264_/B VGND VGND VPWR VPWR _8674_/B sky130_fd_sc_hd__nor2_1
XFILLER_11_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7207_ _6428_/Y _7079_/B _6377_/Y _7059_/A VGND VGND VPWR VPWR _7207_/X sky130_fd_sc_hd__o22a_1
XFILLER_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5468_ _9398_/Q _5460_/A _5967_/B1 _5460_/Y VGND VGND VPWR VPWR _9398_/D sky130_fd_sc_hd__a22o_1
X_8187_ _8187_/A VGND VGND VPWR VPWR _8650_/B sky130_fd_sc_hd__inv_2
X_5399_ _9446_/Q _5395_/A _5963_/B1 _5395_/Y VGND VGND VPWR VPWR _9446_/D sky130_fd_sc_hd__a22o_1
XFILLER_59_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7138_ _6933_/Y _7048_/B _6921_/Y _7077_/A _7137_/X VGND VGND VPWR VPWR _7145_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7069_ _7073_/C _7085_/B VGND VGND VPWR VPWR _7070_/A sky130_fd_sc_hd__or2_1
XFILLER_59_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput19 mask_rev_in[23] VGND VGND VPWR VPWR _6093_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_136_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4770_ _4805_/A _4843_/B VGND VGND VPWR VPWR _5089_/B sky130_fd_sc_hd__or2_4
XFILLER_186_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6440_ _9358_/Q VGND VGND VPWR VPWR _6440_/Y sky130_fd_sc_hd__inv_2
X_6371_ _9260_/Q VGND VGND VPWR VPWR _6371_/Y sky130_fd_sc_hd__inv_4
XFILLER_173_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8110_ _8625_/A _8282_/B _8110_/C VGND VGND VPWR VPWR _8708_/B sky130_fd_sc_hd__and3_2
X_5322_ _9499_/Q _5319_/A _8844_/X _5319_/Y VGND VGND VPWR VPWR _9499_/D sky130_fd_sc_hd__a22o_1
XFILLER_142_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9090_ _9709_/CLK _9090_/D _5988_/X VGND VGND VPWR VPWR _9090_/Q sky130_fd_sc_hd__dfrtp_2
X_8041_ _8041_/A _8685_/A VGND VGND VPWR VPWR _8041_/Y sky130_fd_sc_hd__nor2_1
X_5253_ _5253_/A VGND VGND VPWR VPWR _5253_/Y sky130_fd_sc_hd__inv_2
X_5184_ _9590_/Q _5180_/A _8841_/X _5180_/Y VGND VGND VPWR VPWR _9590_/D sky130_fd_sc_hd__a22o_1
XFILLER_87_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8943_ _9082_/Q _4949_/A _9051_/Q VGND VGND VPWR VPWR _8943_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8874_ _7155_/Y _9633_/Q _8959_/S VGND VGND VPWR VPWR _8874_/X sky130_fd_sc_hd__mux2_1
X_7825_ _7825_/A VGND VGND VPWR VPWR _8515_/A sky130_fd_sc_hd__buf_2
X_7756_ _7832_/A _7756_/B _7837_/C VGND VGND VPWR VPWR _7757_/A sky130_fd_sc_hd__or3_1
XFILLER_184_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4968_ _4994_/A VGND VGND VPWR VPWR _4969_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_137_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6707_ _9304_/Q VGND VGND VPWR VPWR _6707_/Y sky130_fd_sc_hd__inv_2
X_4899_ _9437_/Q VGND VGND VPWR VPWR _4899_/Y sky130_fd_sc_hd__clkinv_2
X_7687_ _6331_/Y _7430_/X _6412_/Y _7432_/X _7686_/X VGND VGND VPWR VPWR _7687_/X
+ sky130_fd_sc_hd__o221a_1
X_9426_ _9527_/CLK _9426_/D _9528_/SET_B VGND VGND VPWR VPWR _9426_/Q sky130_fd_sc_hd__dfrtp_1
X_6638_ _9228_/Q VGND VGND VPWR VPWR _6638_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_192_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9357_ _9358_/CLK _9357_/D _9685_/SET_B VGND VGND VPWR VPWR _9357_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_138_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8308_ _7836_/A _8299_/A _7836_/B _7879_/Y VGND VGND VPWR VPWR _8497_/A sky130_fd_sc_hd__a31o_1
X_6569_ _9735_/Q VGND VGND VPWR VPWR _6569_/Y sky130_fd_sc_hd__inv_2
X_9288_ _9483_/CLK _9288_/D _9528_/SET_B VGND VGND VPWR VPWR _9288_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_16_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR _9344_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_133_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8239_ _8341_/A _8239_/B VGND VGND VPWR VPWR _8361_/B sky130_fd_sc_hd__nor2_1
XFILLER_59_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5940_ _9059_/Q _7731_/A _9119_/Q _5938_/Y _5939_/X VGND VGND VPWR VPWR _9119_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_92_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5871_ _9159_/Q _5866_/A _8839_/X _5866_/Y VGND VGND VPWR VPWR _9159_/D sky130_fd_sc_hd__a22o_1
X_7610_ _4920_/Y _7400_/X _4731_/A _7405_/X _7609_/X VGND VGND VPWR VPWR _7626_/A
+ sky130_fd_sc_hd__o221a_1
X_8590_ _8605_/B _8543_/Y _8564_/X _8589_/X VGND VGND VPWR VPWR _8590_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_61_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4822_ _6158_/A _4929_/A VGND VGND VPWR VPWR _4822_/X sky130_fd_sc_hd__or2_4
XFILLER_193_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4753_ _9789_/Q VGND VGND VPWR VPWR _4753_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7541_ _6422_/Y _7427_/X _6360_/Y _5699_/X VGND VGND VPWR VPWR _7541_/X sky130_fd_sc_hd__o22a_1
X_7472_ _7472_/A _7476_/C _9255_/Q VGND VGND VPWR VPWR _7473_/A sky130_fd_sc_hd__or3_1
X_9211_ _9613_/CLK _9211_/D _9646_/SET_B VGND VGND VPWR VPWR _9211_/Q sky130_fd_sc_hd__dfrtp_1
X_4684_ _4675_/Y _5507_/B _4677_/Y _5080_/B _4683_/X VGND VGND VPWR VPWR _4705_/B
+ sky130_fd_sc_hd__o221a_1
X_6423_ _9410_/Q VGND VGND VPWR VPWR _6423_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_174_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9142_ _9280_/CLK _9142_/D _9757_/SET_B VGND VGND VPWR VPWR _9142_/Q sky130_fd_sc_hd__dfrtp_1
X_6354_ _9631_/Q VGND VGND VPWR VPWR _6354_/Y sky130_fd_sc_hd__inv_2
X_9073_ _9687_/CLK _9073_/D _9685_/SET_B VGND VGND VPWR VPWR _9073_/Q sky130_fd_sc_hd__dfrtp_2
X_6285_ _7238_/A _5610_/B _6284_/Y _5837_/B VGND VGND VPWR VPWR _6285_/X sky130_fd_sc_hd__o22a_1
X_5305_ _9510_/Q _5300_/A _5967_/B1 _5300_/Y VGND VGND VPWR VPWR _9510_/D sky130_fd_sc_hd__a22o_1
XFILLER_142_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8024_ _8521_/A _8137_/B VGND VGND VPWR VPWR _8407_/A sky130_fd_sc_hd__or2_1
X_5236_ _9557_/Q _5234_/A _5964_/B1 _5234_/Y VGND VGND VPWR VPWR _9557_/D sky130_fd_sc_hd__a22o_1
XFILLER_124_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5167_ _5545_/A _6322_/A VGND VGND VPWR VPWR _5168_/A sky130_fd_sc_hd__or2_1
XFILLER_130_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5098_ _9647_/Q _5091_/A _8930_/A1 _5091_/Y VGND VGND VPWR VPWR _9647_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8926_ _9605_/Q _8842_/X _8926_/S VGND VGND VPWR VPWR _8926_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8857_ _8856_/X _9167_/Q _9054_/Q VGND VGND VPWR VPWR _8857_/X sky130_fd_sc_hd__mux2_1
X_8788_ _8788_/A VGND VGND VPWR VPWR _8788_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_169_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7808_ _8660_/C _8119_/A VGND VGND VPWR VPWR _8587_/A sky130_fd_sc_hd__nor2_2
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7739_ _9068_/Q _7739_/A2 _9067_/Q _7739_/B2 _7738_/X VGND VGND VPWR VPWR _7739_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_137_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9409_ _9493_/CLK _9409_/D _4628_/A VGND VGND VPWR VPWR _9409_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_165_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6070_ _6065_/Y _5837_/B _6066_/Y _5660_/B _6069_/X VGND VGND VPWR VPWR _6071_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_112_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5021_ _9690_/Q _5015_/A _8955_/A1 _5015_/Y VGND VGND VPWR VPWR _9690_/D sky130_fd_sc_hd__a22o_1
XFILLER_66_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9760_ _9770_/CLK _9760_/D _7011_/B VGND VGND VPWR VPWR _9760_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_38_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8711_ _8117_/A _8624_/X _8117_/B _8625_/Y _8710_/Y VGND VGND VPWR VPWR _8712_/B
+ sky130_fd_sc_hd__o221ai_4
X_6972_ _4936_/Y _6964_/A _9020_/Q _6964_/Y VGND VGND VPWR VPWR _9020_/D sky130_fd_sc_hd__o22a_1
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9691_ _9695_/CLK _9691_/D _9779_/SET_B VGND VGND VPWR VPWR _9691_/Q sky130_fd_sc_hd__dfrtp_1
X_5923_ _9120_/Q _5918_/A _5967_/B1 _5918_/Y VGND VGND VPWR VPWR _9120_/D sky130_fd_sc_hd__a22o_1
X_8642_ _8642_/A _8642_/B _8642_/C _8642_/D VGND VGND VPWR VPWR _8731_/A sky130_fd_sc_hd__or4_2
X_5854_ _5849_/X _8865_/X _8924_/X _9172_/Q VGND VGND VPWR VPWR _9172_/D sky130_fd_sc_hd__o22a_1
X_8573_ _8573_/A _8573_/B _8573_/C VGND VGND VPWR VPWR _8642_/D sky130_fd_sc_hd__or3_1
X_4805_ _4805_/A _4931_/B VGND VGND VPWR VPWR _5534_/B sky130_fd_sc_hd__or2_4
XFILLER_119_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5785_ _9219_/Q _5778_/A _8930_/A1 _5778_/Y VGND VGND VPWR VPWR _9219_/D sky130_fd_sc_hd__a22o_1
X_7524_ _8779_/A _7434_/X _8777_/A _7436_/X VGND VGND VPWR VPWR _7524_/X sky130_fd_sc_hd__o22a_1
X_4736_ _4732_/Y _5621_/B _4734_/Y _5797_/B VGND VGND VPWR VPWR _4736_/X sky130_fd_sc_hd__o22a_1
XFILLER_9_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4667_ _4898_/A _4843_/B VGND VGND VPWR VPWR _5905_/B sky130_fd_sc_hd__or2_4
X_7455_ _7455_/A VGND VGND VPWR VPWR _7455_/X sky130_fd_sc_hd__buf_8
XFILLER_162_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7386_ _6369_/Y _7048_/D _6445_/Y _7040_/B _7385_/X VGND VGND VPWR VPWR _7387_/D
+ sky130_fd_sc_hd__o221a_1
X_6406_ _6404_/Y _5480_/B _6405_/Y _4577_/B VGND VGND VPWR VPWR _6406_/X sky130_fd_sc_hd__o22a_1
XFILLER_122_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9125_ _9379_/CLK _9125_/D _9646_/SET_B VGND VGND VPWR VPWR _9125_/Q sky130_fd_sc_hd__dfstp_1
X_6337_ _9129_/Q VGND VGND VPWR VPWR _6337_/Y sky130_fd_sc_hd__clkinv_2
X_4598_ _9734_/Q _4592_/A _5965_/B1 _4592_/Y VGND VGND VPWR VPWR _9734_/D sky130_fd_sc_hd__a22o_1
XFILLER_88_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6268_ _9767_/Q VGND VGND VPWR VPWR _6268_/Y sky130_fd_sc_hd__clkinv_2
X_9056_ _9203_/CLK _9056_/D _9633_/SET_B VGND VGND VPWR VPWR _9056_/Q sky130_fd_sc_hd__dfrtp_4
X_5219_ _9568_/Q _5218_/Y _8917_/X _5218_/A VGND VGND VPWR VPWR _9568_/D sky130_fd_sc_hd__o22a_1
X_8007_ _8003_/Y _8566_/B _8064_/C VGND VGND VPWR VPWR _8016_/A sky130_fd_sc_hd__o21a_1
X_6199_ _9552_/Q VGND VGND VPWR VPWR _6199_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8909_ _7730_/Y _9699_/Q _9048_/Q VGND VGND VPWR VPWR _8909_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5570_ _9329_/Q _5566_/A _5966_/B1 _5566_/Y VGND VGND VPWR VPWR _9329_/D sky130_fd_sc_hd__a22o_1
XFILLER_144_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4521_ _4521_/A VGND VGND VPWR VPWR _9770_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7240_ _6291_/Y _7126_/X _6241_/Y _7128_/X VGND VGND VPWR VPWR _7240_/X sky130_fd_sc_hd__o22a_1
X_4452_ _8939_/X VGND VGND VPWR VPWR _5133_/A sky130_fd_sc_hd__clkinv_2
XFILLER_144_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7171_ _6775_/Y _7059_/D _6724_/Y _7116_/X _7170_/X VGND VGND VPWR VPWR _7176_/B
+ sky130_fd_sc_hd__o221a_1
X_6122_ _9238_/Q VGND VGND VPWR VPWR _6122_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6053_ _6053_/A VGND VGND VPWR VPWR _6054_/A sky130_fd_sc_hd__clkbuf_2
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5004_ _5004_/A VGND VGND VPWR VPWR _5004_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_66_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6955_ _6326_/Y _6952_/A _9033_/Q _6952_/Y VGND VGND VPWR VPWR _9033_/D sky130_fd_sc_hd__o22a_1
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9743_ _9777_/CLK _9743_/D _9757_/SET_B VGND VGND VPWR VPWR _9743_/Q sky130_fd_sc_hd__dfstp_1
X_5906_ _5906_/A VGND VGND VPWR VPWR _5907_/A sky130_fd_sc_hd__clkbuf_4
X_9674_ _9674_/CLK _9674_/D _9633_/SET_B VGND VGND VPWR VPWR _9674_/Q sky130_fd_sc_hd__dfrtp_1
X_8625_ _8625_/A _8625_/B VGND VGND VPWR VPWR _8625_/Y sky130_fd_sc_hd__nor2_1
X_6886_ _9045_/Q VGND VGND VPWR VPWR _6886_/Y sky130_fd_sc_hd__inv_2
XFILLER_179_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5837_ _6052_/A _5837_/B VGND VGND VPWR VPWR _5838_/A sky130_fd_sc_hd__or2_1
XFILLER_22_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8556_ _8601_/D VGND VGND VPWR VPWR _8556_/Y sky130_fd_sc_hd__inv_2
X_5768_ _5960_/A _5768_/B VGND VGND VPWR VPWR _5769_/A sky130_fd_sc_hd__or2_1
X_8487_ _8487_/A _8486_/X VGND VGND VPWR VPWR _8488_/A sky130_fd_sc_hd__or2b_1
X_7507_ _6754_/Y _7430_/X _6761_/Y _7432_/X _7506_/X VGND VGND VPWR VPWR _7507_/X
+ sky130_fd_sc_hd__o221a_1
X_4719_ _4903_/B _4780_/B VGND VGND VPWR VPWR _5594_/B sky130_fd_sc_hd__or2_4
X_7438_ _4664_/Y _7430_/X _4793_/Y _7432_/X _7437_/X VGND VGND VPWR VPWR _7438_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_30_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5699_ _5699_/A VGND VGND VPWR VPWR _5699_/X sky130_fd_sc_hd__buf_8
XFILLER_162_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7369_ _6516_/Y _7059_/D _6555_/Y _7116_/X _7368_/X VGND VGND VPWR VPWR _7374_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_89_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9108_ _9379_/CLK _9108_/D _9779_/SET_B VGND VGND VPWR VPWR _9108_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9039_ _9039_/CLK _9039_/D VGND VGND VPWR VPWR _9039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6740_ _6735_/Y _5278_/B _6736_/Y _5344_/B _6739_/X VGND VGND VPWR VPWR _6741_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_35_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6671_ _6669_/Y _4832_/X _6670_/Y _4590_/B VGND VGND VPWR VPWR _6671_/X sky130_fd_sc_hd__o22a_1
X_9390_ _9483_/CLK _9390_/D _9528_/SET_B VGND VGND VPWR VPWR _9390_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_188_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5622_ _5622_/A VGND VGND VPWR VPWR _5623_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_149_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8410_ _8410_/A VGND VGND VPWR VPWR _8734_/B sky130_fd_sc_hd__inv_2
X_5553_ _9340_/Q _5547_/A _8841_/X _5547_/Y VGND VGND VPWR VPWR _9340_/D sky130_fd_sc_hd__a22o_1
XFILLER_136_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8341_ _8341_/A _8341_/B _8496_/A VGND VGND VPWR VPWR _8594_/B sky130_fd_sc_hd__nor3_1
XFILLER_117_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4504_ _5259_/A _4504_/B VGND VGND VPWR VPWR _4505_/A sky130_fd_sc_hd__or2_1
XFILLER_144_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8272_ _8272_/A _8660_/B _8496_/A VGND VGND VPWR VPWR _8715_/B sky130_fd_sc_hd__nor3_1
X_5484_ _9388_/Q _5482_/A _5964_/B1 _5482_/Y VGND VGND VPWR VPWR _9388_/D sky130_fd_sc_hd__a22o_1
X_7223_ _6309_/Y _7077_/C _6287_/Y _7077_/D _7222_/X VGND VGND VPWR VPWR _7223_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7154_ _7154_/A _7154_/B _7154_/C _7154_/D VGND VGND VPWR VPWR _7155_/C sky130_fd_sc_hd__and4_1
XFILLER_104_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6105_ _9639_/Q VGND VGND VPWR VPWR _6105_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7085_ _7127_/C _7085_/B VGND VGND VPWR VPWR _7086_/A sky130_fd_sc_hd__or2_1
XFILLER_58_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6036_ _9071_/Q _6029_/A _8840_/X _6029_/Y VGND VGND VPWR VPWR _9071_/D sky130_fd_sc_hd__a22o_1
XFILLER_100_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7987_ _8551_/A VGND VGND VPWR VPWR _7987_/Y sky130_fd_sc_hd__inv_2
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6938_ _9308_/Q VGND VGND VPWR VPWR _6938_/Y sky130_fd_sc_hd__clkinv_2
X_9726_ _9769_/CLK _9726_/D _7011_/B VGND VGND VPWR VPWR _9726_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6869_ _6867_/Y _5442_/B _6868_/Y _5251_/B VGND VGND VPWR VPWR _6869_/X sky130_fd_sc_hd__o22a_1
X_9657_ _9779_/CLK _9657_/D _9779_/SET_B VGND VGND VPWR VPWR _9657_/Q sky130_fd_sc_hd__dfrtp_1
X_9588_ _9601_/CLK _9588_/D _9295_/SET_B VGND VGND VPWR VPWR _9588_/Q sky130_fd_sc_hd__dfrtp_1
X_8608_ _8496_/A _8515_/B _8305_/B _8019_/C _8447_/X VGND VGND VPWR VPWR _8609_/A
+ sky130_fd_sc_hd__o311a_1
XFILLER_22_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8539_ _8539_/A _8721_/C _8538_/X VGND VGND VPWR VPWR _8705_/D sky130_fd_sc_hd__or3b_2
XFILLER_182_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7910_ _8515_/B _8239_/B VGND VGND VPWR VPWR _7910_/X sky130_fd_sc_hd__or2_1
X_8890_ _7331_/Y _9628_/Q _8959_/S VGND VGND VPWR VPWR _8890_/X sky130_fd_sc_hd__mux2_1
X_7841_ _7841_/A VGND VGND VPWR VPWR _8515_/B sky130_fd_sc_hd__buf_12
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7772_ _7903_/C VGND VGND VPWR VPWR _7959_/A sky130_fd_sc_hd__inv_2
X_4984_ _4984_/A VGND VGND VPWR VPWR _4984_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_23_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6723_ _9439_/Q VGND VGND VPWR VPWR _6723_/Y sky130_fd_sc_hd__inv_2
X_9511_ _9514_/CLK _9511_/D _4628_/A VGND VGND VPWR VPWR _9511_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_51_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6654_ _6652_/Y _4504_/B _6653_/Y _5178_/B VGND VGND VPWR VPWR _6654_/X sky130_fd_sc_hd__o22a_1
X_9442_ _9791_/CLK _9442_/D _9633_/SET_B VGND VGND VPWR VPWR _9442_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_164_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5605_ _9306_/Q _5604_/A _8843_/X _5604_/Y VGND VGND VPWR VPWR _9306_/D sky130_fd_sc_hd__a22o_1
XFILLER_31_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9373_ _9379_/CLK _9373_/D _9779_/SET_B VGND VGND VPWR VPWR _9373_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6585_ _8745_/A _5013_/B _6581_/Y _5789_/B _6584_/X VGND VGND VPWR VPWR _6586_/C
+ sky130_fd_sc_hd__o221a_1
X_5536_ _5536_/A VGND VGND VPWR VPWR _5536_/Y sky130_fd_sc_hd__inv_2
X_8324_ _8324_/A _8498_/B VGND VGND VPWR VPWR _8506_/C sky130_fd_sc_hd__nor2_1
XFILLER_132_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5467_ _9399_/Q _5460_/A _5966_/B1 _5460_/Y VGND VGND VPWR VPWR _9399_/D sky130_fd_sc_hd__a22o_1
X_8255_ _8255_/A _8493_/B VGND VGND VPWR VPWR _8257_/A sky130_fd_sc_hd__or2_1
X_7206_ _6396_/Y _7095_/X _6368_/Y _7068_/D _7205_/X VGND VGND VPWR VPWR _7211_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_87_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8186_ _8186_/A VGND VGND VPWR VPWR _8672_/C sky130_fd_sc_hd__clkinv_2
X_5398_ _9447_/Q _5395_/A _8844_/X _5395_/Y VGND VGND VPWR VPWR _9447_/D sky130_fd_sc_hd__a22o_1
XFILLER_113_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7137_ _6910_/Y _7040_/C _6799_/Y _7059_/C VGND VGND VPWR VPWR _7137_/X sky130_fd_sc_hd__o22a_1
XFILLER_59_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7068_ _7068_/A _7068_/B _7068_/C _7068_/D VGND VGND VPWR VPWR _7078_/C sky130_fd_sc_hd__and4_1
X_6019_ _6019_/A VGND VGND VPWR VPWR _9081_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9709_ _9709_/CLK _9709_/D _4948_/X VGND VGND VPWR VPWR _9709_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6370_ _6368_/Y _5757_/B _6369_/Y _5810_/B VGND VGND VPWR VPWR _6370_/X sky130_fd_sc_hd__o22a_1
XFILLER_9_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5321_ _9500_/Q _5319_/A _8845_/X _5319_/Y VGND VGND VPWR VPWR _9500_/D sky130_fd_sc_hd__a22o_1
XFILLER_127_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8040_ _8624_/B _8552_/A VGND VGND VPWR VPWR _8685_/A sky130_fd_sc_hd__nor2_1
X_5252_ _5252_/A VGND VGND VPWR VPWR _5253_/A sky130_fd_sc_hd__clkbuf_2
X_5183_ _9591_/Q _5180_/A _8842_/X _5180_/Y VGND VGND VPWR VPWR _9591_/D sky130_fd_sc_hd__a22o_1
XFILLER_3_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8942_ _9089_/Q _9088_/Q _9051_/Q VGND VGND VPWR VPWR _8942_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8873_ _8872_/X _9175_/Q _9054_/Q VGND VGND VPWR VPWR _8873_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7824_ _8538_/C _7899_/A _8084_/A VGND VGND VPWR VPWR _7825_/A sky130_fd_sc_hd__or3_1
XFILLER_24_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4967_ _9707_/Q _4966_/A _9706_/Q _4966_/Y VGND VGND VPWR VPWR _9707_/D sky130_fd_sc_hd__a22o_1
X_7755_ _8660_/A VGND VGND VPWR VPWR _8299_/A sky130_fd_sc_hd__inv_2
X_7686_ _6330_/Y _7434_/X _6347_/Y _7436_/X VGND VGND VPWR VPWR _7686_/X sky130_fd_sc_hd__o22a_1
X_6706_ _6706_/A VGND VGND VPWR VPWR _6706_/Y sky130_fd_sc_hd__clkinv_4
X_4898_ _4898_/A _4931_/B VGND VGND VPWR VPWR _5344_/B sky130_fd_sc_hd__or2_4
XFILLER_192_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9425_ _9527_/CLK _9425_/D _9647_/SET_B VGND VGND VPWR VPWR _9425_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_149_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6637_ _9206_/Q VGND VGND VPWR VPWR _6637_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9356_ _9358_/CLK _9356_/D _9685_/SET_B VGND VGND VPWR VPWR _9356_/Q sky130_fd_sc_hd__dfstp_1
X_6568_ _9497_/Q VGND VGND VPWR VPWR _8789_/A sky130_fd_sc_hd__clkinv_8
XFILLER_164_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8307_ _8305_/B _8264_/B _8441_/A VGND VGND VPWR VPWR _8310_/B sky130_fd_sc_hd__o21ai_1
X_5519_ _5519_/A VGND VGND VPWR VPWR _5520_/A sky130_fd_sc_hd__clkbuf_2
X_9287_ _9483_/CLK _9287_/D _9528_/SET_B VGND VGND VPWR VPWR _9287_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_133_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6499_ _6497_/Y _5742_/B _6498_/Y _5810_/B VGND VGND VPWR VPWR _6499_/X sky130_fd_sc_hd__o22a_1
XFILLER_154_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8238_ _8238_/A _8260_/B VGND VGND VPWR VPWR _8574_/B sky130_fd_sc_hd__nor2_1
X_8169_ _8169_/A VGND VGND VPWR VPWR _8373_/A sky130_fd_sc_hd__inv_2
XFILLER_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5870_ _9160_/Q _5866_/A _5966_/B1 _5866_/Y VGND VGND VPWR VPWR _9160_/D sky130_fd_sc_hd__a22o_1
X_4821_ _4821_/A VGND VGND VPWR VPWR _4821_/Y sky130_fd_sc_hd__inv_2
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4752_ _4787_/A _4929_/A VGND VGND VPWR VPWR _5545_/B sky130_fd_sc_hd__or2_4
X_7540_ _6372_/Y _7415_/X _6462_/Y _7417_/X _7539_/X VGND VGND VPWR VPWR _7554_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4683_ input61/X _4680_/Y _4681_/Y _6052_/C VGND VGND VPWR VPWR _4683_/X sky130_fd_sc_hd__o2bb2a_1
X_7471_ _7471_/A VGND VGND VPWR VPWR _7471_/X sky130_fd_sc_hd__buf_8
X_9210_ _9652_/CLK _9210_/D _9647_/SET_B VGND VGND VPWR VPWR _9210_/Q sky130_fd_sc_hd__dfrtp_1
X_6422_ _9446_/Q VGND VGND VPWR VPWR _6422_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_146_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9141_ _9279_/CLK _9141_/D _9757_/SET_B VGND VGND VPWR VPWR _9141_/Q sky130_fd_sc_hd__dfrtp_1
X_6353_ _9194_/Q VGND VGND VPWR VPWR _6353_/Y sky130_fd_sc_hd__clkinv_2
X_9072_ _9358_/CLK _9072_/D _9685_/SET_B VGND VGND VPWR VPWR _9072_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_161_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6284_ _9182_/Q VGND VGND VPWR VPWR _6284_/Y sky130_fd_sc_hd__inv_2
X_5304_ _9511_/Q _5300_/A _5966_/B1 _5300_/Y VGND VGND VPWR VPWR _9511_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8023_ _8389_/A _8130_/B _8020_/X _8403_/A _8450_/A VGND VGND VPWR VPWR _8023_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_88_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5235_ _9558_/Q _5234_/A _5963_/B1 _5234_/Y VGND VGND VPWR VPWR _9558_/D sky130_fd_sc_hd__a22o_1
XFILLER_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5166_ _9602_/Q _5158_/A _8916_/A1 _5158_/Y VGND VGND VPWR VPWR _9602_/D sky130_fd_sc_hd__a22o_1
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5097_ _9648_/Q _5091_/A _8955_/A1 _5091_/Y VGND VGND VPWR VPWR _9648_/D sky130_fd_sc_hd__a22o_1
XFILLER_110_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8925_ _9606_/Q _8925_/A1 _8926_/S VGND VGND VPWR VPWR _8925_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8856_ _7554_/Y _9636_/Q _8978_/S VGND VGND VPWR VPWR _8856_/X sky130_fd_sc_hd__mux2_1
X_8787_ _8787_/A VGND VGND VPWR VPWR _8788_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_169_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7807_ _8394_/D _8521_/A VGND VGND VPWR VPWR _8119_/A sky130_fd_sc_hd__or2_2
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5999_ _9088_/Q _5995_/A _8913_/X _5995_/Y VGND VGND VPWR VPWR _9088_/D sky130_fd_sc_hd__a22o_1
X_7738_ _9066_/Q _7738_/B VGND VGND VPWR VPWR _7738_/X sky130_fd_sc_hd__and2_1
XFILLER_33_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9408_ _9493_/CLK _9408_/D _4628_/A VGND VGND VPWR VPWR _9408_/Q sky130_fd_sc_hd__dfstp_1
X_7669_ _6479_/Y _7430_/X _6597_/Y _7432_/X _7668_/X VGND VGND VPWR VPWR _7669_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_137_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9339_ _9508_/CLK _9339_/D _9647_/SET_B VGND VGND VPWR VPWR _9339_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_121_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput290 _9755_/Q VGND VGND VPWR VPWR pll_trim[23] sky130_fd_sc_hd__buf_2
XFILLER_75_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5020_ _9691_/Q _5015_/A _8929_/A1 _5015_/Y VGND VGND VPWR VPWR _9691_/D sky130_fd_sc_hd__a22o_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8710_ _8710_/A VGND VGND VPWR VPWR _8710_/Y sky130_fd_sc_hd__inv_2
X_6971_ _6946_/Y _6964_/A _9021_/Q _6964_/Y VGND VGND VPWR VPWR _9021_/D sky130_fd_sc_hd__o22a_1
XFILLER_80_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9690_ _9695_/CLK _9690_/D _9779_/SET_B VGND VGND VPWR VPWR _9690_/Q sky130_fd_sc_hd__dfrtp_1
X_5922_ _9121_/Q _5918_/A _8930_/A1 _5918_/Y VGND VGND VPWR VPWR _9121_/D sky130_fd_sc_hd__a22o_1
XFILLER_53_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_15_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR _9501_/CLK sky130_fd_sc_hd__clkbuf_16
X_8641_ _8641_/A _8641_/B _8641_/C _8343_/Y VGND VGND VPWR VPWR _8719_/C sky130_fd_sc_hd__or4b_2
XFILLER_80_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5853_ _5849_/X _8867_/X _8924_/X _9173_/Q VGND VGND VPWR VPWR _9173_/D sky130_fd_sc_hd__o22a_1
X_4804_ _9346_/Q VGND VGND VPWR VPWR _4804_/Y sky130_fd_sc_hd__clkinv_4
X_8572_ _8641_/B _8719_/A _8572_/C _8677_/C VGND VGND VPWR VPWR _8576_/A sky130_fd_sc_hd__or4_1
X_5784_ _9220_/Q _5778_/A _8955_/A1 _5778_/Y VGND VGND VPWR VPWR _9220_/D sky130_fd_sc_hd__a22o_1
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4735_ _6158_/B _4780_/B VGND VGND VPWR VPWR _5797_/B sky130_fd_sc_hd__or2_4
X_7523_ _8793_/A _7427_/X _8763_/A _5699_/X VGND VGND VPWR VPWR _7523_/X sky130_fd_sc_hd__o22a_1
XFILLER_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7454_ _7456_/A _7466_/A _7474_/D VGND VGND VPWR VPWR _7455_/A sky130_fd_sc_hd__or3_1
X_4666_ _4666_/A VGND VGND VPWR VPWR _4843_/B sky130_fd_sc_hd__buf_8
XFILLER_134_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7385_ _6373_/Y _7068_/A _6412_/Y _7105_/X VGND VGND VPWR VPWR _7385_/X sky130_fd_sc_hd__o22a_1
X_6405_ _9744_/Q VGND VGND VPWR VPWR _6405_/Y sky130_fd_sc_hd__inv_2
X_4597_ _9735_/Q _4592_/A _5964_/B1 _4592_/Y VGND VGND VPWR VPWR _9735_/D sky130_fd_sc_hd__a22o_1
XFILLER_162_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9124_ _9655_/CLK _9124_/D _7011_/B VGND VGND VPWR VPWR _9124_/Q sky130_fd_sc_hd__dfrtp_1
X_6336_ _6336_/A VGND VGND VPWR VPWR _6336_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9055_ _9203_/CLK _9055_/D _9633_/SET_B VGND VGND VPWR VPWR _9055_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_170_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6267_ _6262_/Y _4907_/X _6263_/Y _5240_/B _6266_/X VGND VGND VPWR VPWR _6280_/B
+ sky130_fd_sc_hd__o221a_1
X_5218_ _5218_/A VGND VGND VPWR VPWR _5218_/Y sky130_fd_sc_hd__inv_2
X_8006_ _8525_/C VGND VGND VPWR VPWR _8064_/C sky130_fd_sc_hd__clkinv_2
X_6198_ _6193_/Y _6322_/A _6194_/Y _5837_/B _6197_/X VGND VGND VPWR VPWR _6211_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_130_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5149_ _9616_/Q _5147_/A _8845_/X _5147_/Y VGND VGND VPWR VPWR _9616_/D sky130_fd_sc_hd__a22o_1
XFILLER_151_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8908_ _7726_/Y _4949_/A _9048_/Q VGND VGND VPWR VPWR _8908_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8839_ _4949_/A _9659_/Q _9587_/Q VGND VGND VPWR VPWR _8839_/X sky130_fd_sc_hd__mux2_8
XFILLER_25_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4520_ _5967_/B1 _9770_/Q _4520_/S VGND VGND VPWR VPWR _4521_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4451_ _9575_/Q _4901_/A _9081_/Q VGND VGND VPWR VPWR _8990_/A sky130_fd_sc_hd__mux2_1
X_7170_ _6694_/Y _7118_/X _6686_/Y _7048_/C VGND VGND VPWR VPWR _7170_/X sky130_fd_sc_hd__o22a_1
X_6121_ _9211_/Q VGND VGND VPWR VPWR _6121_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_98_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6052_ _6052_/A _6052_/B _6052_/C VGND VGND VPWR VPWR _6053_/A sky130_fd_sc_hd__or3_2
XFILLER_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5003_ _6040_/A VGND VGND VPWR VPWR _5004_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_38_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6954_ _6237_/Y _6952_/A _9034_/Q _6952_/Y VGND VGND VPWR VPWR _9034_/D sky130_fd_sc_hd__o22a_1
X_9742_ _9777_/CLK _9742_/D _9757_/SET_B VGND VGND VPWR VPWR _9742_/Q sky130_fd_sc_hd__dfstp_1
X_5905_ _6052_/A _5905_/B VGND VGND VPWR VPWR _5906_/A sky130_fd_sc_hd__or2_1
X_9673_ _9674_/CLK _9673_/D _9633_/SET_B VGND VGND VPWR VPWR _9673_/Q sky130_fd_sc_hd__dfrtp_1
X_8624_ _8632_/A _8624_/B VGND VGND VPWR VPWR _8624_/X sky130_fd_sc_hd__and2_1
XFILLER_22_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6885_ _9329_/Q VGND VGND VPWR VPWR _6885_/Y sky130_fd_sc_hd__inv_2
X_5836_ _9185_/Q _5831_/A _5967_/B1 _5831_/Y VGND VGND VPWR VPWR _9185_/D sky130_fd_sc_hd__a22o_1
X_5767_ _9231_/Q _5759_/A _8839_/X _5759_/Y VGND VGND VPWR VPWR _9231_/D sky130_fd_sc_hd__a22o_1
X_8555_ _8119_/A _8397_/B _8168_/A _8401_/B _8169_/A VGND VGND VPWR VPWR _8631_/B
+ sky130_fd_sc_hd__o221ai_1
X_8486_ _8514_/B _8485_/X VGND VGND VPWR VPWR _8486_/X sky130_fd_sc_hd__or2b_1
X_4718_ _9307_/Q VGND VGND VPWR VPWR _4718_/Y sky130_fd_sc_hd__inv_2
X_7506_ _6694_/Y _7434_/X _6760_/Y _7436_/X VGND VGND VPWR VPWR _7506_/X sky130_fd_sc_hd__o22a_1
X_5698_ _7456_/A _7462_/A _7474_/D VGND VGND VPWR VPWR _5699_/A sky130_fd_sc_hd__or3_1
XFILLER_162_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7437_ _4846_/Y _7434_/X _4926_/Y _7436_/X VGND VGND VPWR VPWR _7437_/X sky130_fd_sc_hd__o22a_1
X_4649_ _9714_/Q _4636_/A _8949_/X _4636_/Y VGND VGND VPWR VPWR _9714_/D sky130_fd_sc_hd__a22o_1
XFILLER_162_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7368_ _6606_/Y _7118_/X _6503_/Y _7048_/C VGND VGND VPWR VPWR _7368_/X sky130_fd_sc_hd__o22a_1
X_6319_ _6314_/Y _5089_/B _6315_/Y _5949_/B _6318_/X VGND VGND VPWR VPWR _6325_/B
+ sky130_fd_sc_hd__o221a_1
X_9107_ _9378_/CLK _9107_/D _9646_/SET_B VGND VGND VPWR VPWR _9107_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_89_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7299_ _7299_/A _7299_/B _7299_/C _7299_/D VGND VGND VPWR VPWR _7309_/B sky130_fd_sc_hd__and4_1
XFILLER_39_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9038_ _9664_/CLK _9038_/D VGND VGND VPWR VPWR _9038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6670_ _9734_/Q VGND VGND VPWR VPWR _6670_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_176_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5621_ _6052_/A _5621_/B VGND VGND VPWR VPWR _5622_/A sky130_fd_sc_hd__or2_1
X_8340_ _8079_/C _8340_/B _8340_/C _8394_/A VGND VGND VPWR VPWR _8722_/A sky130_fd_sc_hd__and4b_1
X_5552_ _9341_/Q _5547_/A _8929_/A1 _5547_/Y VGND VGND VPWR VPWR _9341_/D sky130_fd_sc_hd__a22o_1
X_8271_ _8271_/A _8506_/B VGND VGND VPWR VPWR _8273_/A sky130_fd_sc_hd__or2_1
X_4503_ _4911_/A _4921_/A VGND VGND VPWR VPWR _4504_/B sky130_fd_sc_hd__or2_4
XFILLER_117_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5483_ _9389_/Q _5482_/A _5963_/B1 _5482_/Y VGND VGND VPWR VPWR _9389_/D sky130_fd_sc_hd__a22o_1
XFILLER_144_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7222_ _6274_/Y _7086_/X _6239_/Y _7088_/X VGND VGND VPWR VPWR _7222_/X sky130_fd_sc_hd__o22a_1
X_7153_ _6871_/Y _7124_/X _6884_/Y _7068_/B _7152_/X VGND VGND VPWR VPWR _7154_/D
+ sky130_fd_sc_hd__o221a_1
X_6104_ _9077_/Q VGND VGND VPWR VPWR _6104_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_98_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7084_ _7084_/A VGND VGND VPWR VPWR _7084_/X sky130_fd_sc_hd__buf_8
X_6035_ _9072_/Q _6029_/A _8841_/X _6029_/Y VGND VGND VPWR VPWR _9072_/D sky130_fd_sc_hd__a22o_1
XFILLER_112_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7986_ _7986_/A VGND VGND VPWR VPWR _8551_/A sky130_fd_sc_hd__buf_2
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9725_ _9769_/CLK _9725_/D _9757_/SET_B VGND VGND VPWR VPWR _9725_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6937_ _6932_/Y _5789_/B _6933_/Y _5818_/B _6936_/X VGND VGND VPWR VPWR _6944_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_25_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6868_ _9542_/Q VGND VGND VPWR VPWR _6868_/Y sky130_fd_sc_hd__inv_2
X_9656_ _9779_/CLK _9656_/D _9779_/SET_B VGND VGND VPWR VPWR _9656_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_167_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9587_ _4450_/A1 _9587_/D _6146_/A VGND VGND VPWR VPWR _9587_/Q sky130_fd_sc_hd__dfrtp_4
X_5819_ _5819_/A VGND VGND VPWR VPWR _5820_/A sky130_fd_sc_hd__clkbuf_4
X_8607_ _8607_/A _8607_/B _8607_/C _7910_/X VGND VGND VPWR VPWR _8735_/A sky130_fd_sc_hd__or4b_2
X_8538_ _8583_/A _8538_/B _8538_/C _8538_/D VGND VGND VPWR VPWR _8538_/X sky130_fd_sc_hd__or4_1
XFILLER_155_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6799_ _9126_/Q VGND VGND VPWR VPWR _6799_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8469_ _7848_/A _8305_/A _8097_/B _8554_/A VGND VGND VPWR VPWR _8698_/A sky130_fd_sc_hd__o22ai_1
XFILLER_123_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput190 wb_dat_i[3] VGND VGND VPWR VPWR _8964_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_83_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7840_ _8379_/D _8394_/B _8394_/C _8195_/A VGND VGND VPWR VPWR _7841_/A sky130_fd_sc_hd__or4_1
XFILLER_36_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7771_ _7771_/A _7771_/B _7771_/C _7771_/D VGND VGND VPWR VPWR _7775_/C sky130_fd_sc_hd__nand4_1
X_4983_ _4994_/A VGND VGND VPWR VPWR _4984_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6722_ _6717_/Y _5317_/B _6718_/Y _5518_/B _6721_/X VGND VGND VPWR VPWR _6741_/A
+ sky130_fd_sc_hd__o221a_1
X_9510_ _9514_/CLK _9510_/D _4628_/A VGND VGND VPWR VPWR _9510_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6653_ _8803_/A VGND VGND VPWR VPWR _6653_/Y sky130_fd_sc_hd__inv_2
X_9441_ _9514_/CLK _9441_/D _9685_/SET_B VGND VGND VPWR VPWR _9441_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_149_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5604_ _5604_/A VGND VGND VPWR VPWR _5604_/Y sky130_fd_sc_hd__inv_2
XFILLER_191_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6584_ _6582_/Y _5621_/B _6583_/Y _5526_/B VGND VGND VPWR VPWR _6584_/X sky130_fd_sc_hd__o22a_2
X_9372_ _9379_/CLK _9372_/D _9779_/SET_B VGND VGND VPWR VPWR _9372_/Q sky130_fd_sc_hd__dfstp_1
X_5535_ _5535_/A VGND VGND VPWR VPWR _5536_/A sky130_fd_sc_hd__clkbuf_4
X_8323_ _8463_/A _8645_/B VGND VGND VPWR VPWR _8599_/C sky130_fd_sc_hd__or2_1
XFILLER_11_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5466_ _9400_/Q _5460_/A _5965_/B1 _5460_/Y VGND VGND VPWR VPWR _9400_/D sky130_fd_sc_hd__a22o_1
X_8254_ _8341_/A _8254_/B VGND VGND VPWR VPWR _8493_/B sky130_fd_sc_hd__nor2_1
XFILLER_160_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7205_ _6329_/Y _7097_/X _6349_/Y _7099_/X VGND VGND VPWR VPWR _7205_/X sky130_fd_sc_hd__o22a_1
XFILLER_160_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8185_ _8185_/A VGND VGND VPWR VPWR _8514_/A sky130_fd_sc_hd__inv_2
X_5397_ _9448_/Q _5395_/A _8845_/X _5395_/Y VGND VGND VPWR VPWR _9448_/D sky130_fd_sc_hd__a22o_1
X_7136_ _6825_/Y _7082_/X _6787_/Y _7084_/X _7135_/X VGND VGND VPWR VPWR _7155_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_101_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7067_ _7067_/A VGND VGND VPWR VPWR _7068_/D sky130_fd_sc_hd__clkbuf_16
X_6018_ _8916_/A1 _9081_/Q _6018_/S VGND VGND VPWR VPWR _6019_/A sky130_fd_sc_hd__mux2_1
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7969_ _7969_/A _8120_/B VGND VGND VPWR VPWR _7970_/A sky130_fd_sc_hd__or2_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9708_ _9709_/CLK _9708_/D _4957_/X VGND VGND VPWR VPWR _9708_/Q sky130_fd_sc_hd__dfrtp_2
X_9639_ _9639_/CLK _9639_/D _9633_/SET_B VGND VGND VPWR VPWR _9639_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5320_ _9501_/Q _5319_/A _8846_/X _5319_/Y VGND VGND VPWR VPWR _9501_/D sky130_fd_sc_hd__a22o_1
XFILLER_142_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5251_ _5259_/A _5251_/B VGND VGND VPWR VPWR _5252_/A sky130_fd_sc_hd__or2_1
XFILLER_142_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5182_ _9592_/Q _5180_/A _8925_/A1 _5180_/Y VGND VGND VPWR VPWR _9592_/D sky130_fd_sc_hd__a22o_1
XFILLER_87_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8941_ _8940_/X _9681_/Q _9587_/Q VGND VGND VPWR VPWR _8941_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8872_ _7698_/Y _9631_/Q _8978_/S VGND VGND VPWR VPWR _8872_/X sky130_fd_sc_hd__mux2_1
X_7823_ _7823_/A _7823_/B _8538_/B VGND VGND VPWR VPWR _7899_/A sky130_fd_sc_hd__or3b_1
XFILLER_24_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7754_ _8379_/D _8394_/B _7838_/B VGND VGND VPWR VPWR _8660_/A sky130_fd_sc_hd__or3_4
XFILLER_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4966_ _4966_/A VGND VGND VPWR VPWR _4966_/Y sky130_fd_sc_hd__clkinv_2
X_6705_ _9486_/Q VGND VGND VPWR VPWR _6705_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_51_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4897_ _9476_/Q VGND VGND VPWR VPWR _4897_/Y sky130_fd_sc_hd__clkinv_4
X_7685_ _6391_/Y _7427_/X _6361_/Y _5699_/X VGND VGND VPWR VPWR _7685_/X sky130_fd_sc_hd__o22a_1
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9424_ _9535_/CLK _9424_/D _9528_/SET_B VGND VGND VPWR VPWR _9424_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_137_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6636_ _7172_/A _5610_/B _6632_/Y _5594_/B _6635_/X VGND VGND VPWR VPWR _6649_/A
+ sky130_fd_sc_hd__o221a_1
X_9355_ _9358_/CLK _9355_/D _9685_/SET_B VGND VGND VPWR VPWR _9355_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_138_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6567_ _6567_/A _6567_/B _6567_/C _6567_/D VGND VGND VPWR VPWR _6628_/A sky130_fd_sc_hd__and4_1
XFILLER_192_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8306_ _8521_/B _7885_/B _8447_/B _8215_/X _8397_/A VGND VGND VPWR VPWR _8306_/X
+ sky130_fd_sc_hd__o2111a_1
X_5518_ _5671_/A _5518_/B VGND VGND VPWR VPWR _5519_/A sky130_fd_sc_hd__or2_1
X_9286_ _9483_/CLK _9286_/D _9528_/SET_B VGND VGND VPWR VPWR _9286_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_145_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6498_ _9201_/Q VGND VGND VPWR VPWR _6498_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_160_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5449_ _9411_/Q _5444_/A _5967_/B1 _5444_/Y VGND VGND VPWR VPWR _9411_/D sky130_fd_sc_hd__a22o_1
X_8237_ _8237_/A _8358_/B _8642_/B _8359_/B VGND VGND VPWR VPWR _8241_/A sky130_fd_sc_hd__or4_1
XFILLER_154_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8168_ _8168_/A _8378_/B VGND VGND VPWR VPWR _8169_/A sky130_fd_sc_hd__or2_1
X_7119_ _4846_/Y _7118_/X _4675_/Y _7048_/C VGND VGND VPWR VPWR _7119_/X sky130_fd_sc_hd__o22a_1
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8099_ _8195_/A _8099_/B VGND VGND VPWR VPWR _8100_/A sky130_fd_sc_hd__or2_1
XFILLER_170_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4820_ _4813_/Y _4537_/B _4814_/Y _6027_/B _4819_/X VGND VGND VPWR VPWR _4830_/C
+ sky130_fd_sc_hd__o221a_1
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4751_ _9338_/Q VGND VGND VPWR VPWR _4751_/Y sky130_fd_sc_hd__inv_2
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7470_ _7472_/A _7470_/B _9255_/Q VGND VGND VPWR VPWR _7471_/A sky130_fd_sc_hd__or3_1
X_4682_ _4787_/A _4876_/B VGND VGND VPWR VPWR _6052_/C sky130_fd_sc_hd__or2_4
X_6421_ _9376_/Q VGND VGND VPWR VPWR _6421_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9140_ _9279_/CLK _9140_/D _9757_/SET_B VGND VGND VPWR VPWR _9140_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_161_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6352_ _6352_/A _6352_/B _6352_/C _6352_/D VGND VGND VPWR VPWR _6475_/A sky130_fd_sc_hd__and4_1
X_9071_ _9358_/CLK _9071_/D _9685_/SET_B VGND VGND VPWR VPWR _9071_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_154_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6283_ _9299_/Q VGND VGND VPWR VPWR _7238_/A sky130_fd_sc_hd__clkinv_2
X_5303_ _9512_/Q _5300_/A _5965_/B1 _5300_/Y VGND VGND VPWR VPWR _9512_/D sky130_fd_sc_hd__a22o_1
XFILLER_142_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8022_ _8624_/B _8130_/B VGND VGND VPWR VPWR _8450_/A sky130_fd_sc_hd__or2_1
X_5234_ _5234_/A VGND VGND VPWR VPWR _5234_/Y sky130_fd_sc_hd__inv_2
X_5165_ _9603_/Q _5158_/A _8840_/X _5158_/Y VGND VGND VPWR VPWR _9603_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5096_ _9649_/Q _5091_/A _8929_/A1 _5091_/Y VGND VGND VPWR VPWR _9649_/D sky130_fd_sc_hd__a22o_1
XFILLER_83_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8924_ _9055_/Q _8819_/X _9054_/Q VGND VGND VPWR VPWR _8924_/X sky130_fd_sc_hd__mux2_8
XFILLER_37_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8855_ _8854_/X _9166_/Q _9054_/Q VGND VGND VPWR VPWR _8855_/X sky130_fd_sc_hd__mux2_1
X_7806_ _7806_/A VGND VGND VPWR VPWR _8521_/A sky130_fd_sc_hd__buf_8
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8786_ _8786_/A VGND VGND VPWR VPWR _8786_/X sky130_fd_sc_hd__clkbuf_1
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5998_ _5998_/A VGND VGND VPWR VPWR _5998_/X sky130_fd_sc_hd__clkbuf_1
X_7737_ _9068_/Q _7737_/A2 _9067_/Q _7737_/B2 _7736_/X VGND VGND VPWR VPWR _7737_/X
+ sky130_fd_sc_hd__a221o_1
X_4949_ _4949_/A VGND VGND VPWR VPWR _4949_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_137_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7668_ _6606_/Y _7434_/X _6604_/Y _7436_/X VGND VGND VPWR VPWR _7668_/X sky130_fd_sc_hd__o22a_1
XFILLER_177_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6619_ _6617_/Y _5121_/B _6618_/Y _4870_/X VGND VGND VPWR VPWR _6619_/X sky130_fd_sc_hd__o22a_1
XFILLER_20_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9407_ _9493_/CLK _9407_/D _4628_/A VGND VGND VPWR VPWR _9407_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_153_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7599_ _6074_/Y _7445_/X _6090_/Y _7447_/X VGND VGND VPWR VPWR _7599_/X sky130_fd_sc_hd__o22a_1
XFILLER_165_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9338_ _9535_/CLK _9338_/D _9528_/SET_B VGND VGND VPWR VPWR _9338_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_106_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9269_ _9535_/CLK _9269_/D _9528_/SET_B VGND VGND VPWR VPWR _9269_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_160_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput280 _9746_/Q VGND VGND VPWR VPWR pll_trim[14] sky130_fd_sc_hd__buf_2
XFILLER_121_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput291 _9756_/Q VGND VGND VPWR VPWR pll_trim[24] sky130_fd_sc_hd__buf_2
XFILLER_87_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6970_ _6785_/Y _6964_/A _9022_/Q _6964_/Y VGND VGND VPWR VPWR _9022_/D sky130_fd_sc_hd__o22a_1
XFILLER_81_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5921_ _9122_/Q _5918_/A _5965_/B1 _5918_/Y VGND VGND VPWR VPWR _9122_/D sky130_fd_sc_hd__a22o_1
XFILLER_34_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8640_ _8640_/A _8640_/B _8640_/C VGND VGND VPWR VPWR _8641_/C sky130_fd_sc_hd__nor3_1
X_5852_ _5849_/X _8869_/X _8924_/X _9174_/Q VGND VGND VPWR VPWR _9174_/D sky130_fd_sc_hd__o22a_1
X_8571_ _8571_/A _8571_/B _8571_/C VGND VGND VPWR VPWR _8677_/C sky130_fd_sc_hd__or3_1
X_5783_ _9221_/Q _5778_/A _8929_/A1 _5778_/Y VGND VGND VPWR VPWR _9221_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4803_ _4903_/B _4931_/B VGND VGND VPWR VPWR _5290_/B sky130_fd_sc_hd__or2_4
X_4734_ _9204_/Q VGND VGND VPWR VPWR _4734_/Y sky130_fd_sc_hd__inv_2
X_7522_ _8753_/A _7415_/X _8745_/A _7417_/X _7521_/X VGND VGND VPWR VPWR _7536_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_9_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7453_ _7453_/A VGND VGND VPWR VPWR _7453_/X sky130_fd_sc_hd__buf_8
X_4665_ _8936_/X _4665_/B _4665_/C VGND VGND VPWR VPWR _4666_/A sky130_fd_sc_hd__or3_1
X_7384_ _6393_/Y _7059_/B _6423_/Y _7068_/C _7383_/X VGND VGND VPWR VPWR _7387_/C
+ sky130_fd_sc_hd__o221a_1
X_4596_ _9736_/Q _4592_/A _5963_/B1 _4592_/Y VGND VGND VPWR VPWR _9736_/D sky130_fd_sc_hd__a22o_1
X_6404_ _9389_/Q VGND VGND VPWR VPWR _6404_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_127_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6335_ _9384_/Q VGND VGND VPWR VPWR _6335_/Y sky130_fd_sc_hd__inv_2
X_9123_ _9655_/CLK _9123_/D _9779_/SET_B VGND VGND VPWR VPWR _9123_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_142_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9054_ _9279_/CLK _9054_/D _9633_/SET_B VGND VGND VPWR VPWR _9054_/Q sky130_fd_sc_hd__dfrtp_4
X_8005_ _8005_/A VGND VGND VPWR VPWR _8566_/B sky130_fd_sc_hd__inv_2
XFILLER_103_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6266_ _6264_/Y _5431_/B _6265_/Y _4602_/B VGND VGND VPWR VPWR _6266_/X sky130_fd_sc_hd__o22a_1
X_5217_ _6135_/A _6322_/A _5259_/A _8976_/X VGND VGND VPWR VPWR _5218_/A sky130_fd_sc_hd__a211o_4
X_6197_ _6195_/Y _5355_/B _6196_/Y _5344_/B VGND VGND VPWR VPWR _6197_/X sky130_fd_sc_hd__o22a_1
XFILLER_57_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5148_ _9617_/Q _5147_/A _8846_/X _5147_/Y VGND VGND VPWR VPWR _9617_/D sky130_fd_sc_hd__a22o_1
X_5079_ _5079_/A VGND VGND VPWR VPWR _9659_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8907_ _7725_/X _9088_/Q _9051_/Q VGND VGND VPWR VPWR _8907_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8838_ input85/X _4949_/A _9626_/Q VGND VGND VPWR VPWR _8838_/X sky130_fd_sc_hd__mux2_2
X_8769_ _8769_/A VGND VGND VPWR VPWR _8770_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_25_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4450_ _9576_/Q _4450_/A1 _9788_/Q VGND VGND VPWR VPWR _8991_/A sky130_fd_sc_hd__mux2_1
X_6120_ _9695_/Q VGND VGND VPWR VPWR _6120_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_152_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6051_ _6051_/A VGND VGND VPWR VPWR _6051_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _5002_/A VGND VGND VPWR VPWR _9698_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6953_ _6145_/Y _6952_/A _9035_/Q _6952_/Y VGND VGND VPWR VPWR _9035_/D sky130_fd_sc_hd__o22a_1
X_9741_ _9777_/CLK _9741_/D _9757_/SET_B VGND VGND VPWR VPWR _9741_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6884_ _9313_/Q VGND VGND VPWR VPWR _6884_/Y sky130_fd_sc_hd__clkinv_2
X_5904_ _9133_/Q _5899_/A _8839_/X _5899_/Y VGND VGND VPWR VPWR _9133_/D sky130_fd_sc_hd__a22o_1
X_9672_ _9695_/CLK _9672_/D _9779_/SET_B VGND VGND VPWR VPWR _9672_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_179_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8623_ _8098_/A _8622_/X _8547_/X VGND VGND VPWR VPWR _8710_/A sky130_fd_sc_hd__o21ai_2
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5835_ _9186_/Q _5831_/A _5966_/B1 _5831_/Y VGND VGND VPWR VPWR _9186_/D sky130_fd_sc_hd__a22o_1
XFILLER_139_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5766_ _9232_/Q _5759_/A _8840_/X _5759_/Y VGND VGND VPWR VPWR _9232_/D sky130_fd_sc_hd__a22o_1
X_8554_ _8554_/A _8554_/B VGND VGND VPWR VPWR _8709_/A sky130_fd_sc_hd__nor2_1
XFILLER_22_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8485_ _8485_/A _8514_/C VGND VGND VPWR VPWR _8485_/X sky130_fd_sc_hd__or2_1
X_7505_ _6763_/Y _7427_/X _6661_/Y _5699_/X VGND VGND VPWR VPWR _7505_/X sky130_fd_sc_hd__o22a_1
X_4717_ _4876_/B _4843_/B VGND VGND VPWR VPWR _5837_/B sky130_fd_sc_hd__or2_4
X_5697_ _9255_/Q VGND VGND VPWR VPWR _7474_/D sky130_fd_sc_hd__inv_2
X_4648_ _4648_/A VGND VGND VPWR VPWR _4648_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_30_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7436_ _7436_/A VGND VGND VPWR VPWR _7436_/X sky130_fd_sc_hd__buf_6
XFILLER_162_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9106_ _9379_/CLK _9106_/D _9646_/SET_B VGND VGND VPWR VPWR _9106_/Q sky130_fd_sc_hd__dfstp_1
X_7367_ _6486_/Y _7040_/D _6508_/Y _7110_/X _7366_/X VGND VGND VPWR VPWR _7374_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_89_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4579_ _4579_/A VGND VGND VPWR VPWR _4579_/Y sky130_fd_sc_hd__clkinv_2
X_6318_ _6316_/Y _5660_/B _6317_/Y _6134_/A VGND VGND VPWR VPWR _6318_/X sky130_fd_sc_hd__o22a_1
XFILLER_115_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7298_ _4685_/Y _7048_/D _4823_/Y _7040_/B _7297_/X VGND VGND VPWR VPWR _7299_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9037_ _9664_/CLK _9037_/D VGND VGND VPWR VPWR _9037_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6249_ _6249_/A VGND VGND VPWR VPWR _6249_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_14_csclk clkbuf_2_2_0_csclk/X VGND VGND VPWR VPWR _9534_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_96_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_29_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR _9653_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_63_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5620_ _9294_/Q _5612_/A _8916_/A1 _5612_/Y VGND VGND VPWR VPWR _9294_/D sky130_fd_sc_hd__a22o_1
XFILLER_149_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5551_ _9342_/Q _5547_/A _8925_/A1 _5547_/Y VGND VGND VPWR VPWR _9342_/D sky130_fd_sc_hd__a22o_1
X_8270_ _8341_/A _8270_/B VGND VGND VPWR VPWR _8506_/B sky130_fd_sc_hd__nor2_1
X_4502_ _8934_/X _8932_/X _8946_/X _4729_/B VGND VGND VPWR VPWR _4921_/A sky130_fd_sc_hd__or4_4
XFILLER_172_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7221_ _7221_/A _7221_/B _7221_/C VGND VGND VPWR VPWR _7221_/Y sky130_fd_sc_hd__nand3_4
X_5482_ _5482_/A VGND VGND VPWR VPWR _5482_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7152_ _6823_/Y _7126_/X _6844_/Y _7128_/X VGND VGND VPWR VPWR _7152_/X sky130_fd_sc_hd__o22a_1
X_6103_ _9423_/Q VGND VGND VPWR VPWR _6103_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7083_ _7098_/C _7125_/A _7127_/C VGND VGND VPWR VPWR _7084_/A sky130_fd_sc_hd__or3_1
X_6034_ _9073_/Q _6029_/A _8842_/X _6029_/Y VGND VGND VPWR VPWR _9073_/D sky130_fd_sc_hd__a22o_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7985_ _7997_/B _7992_/B VGND VGND VPWR VPWR _7986_/A sky130_fd_sc_hd__or2_1
XFILLER_54_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6936_ _7326_/A _5632_/B _6935_/Y _5768_/B VGND VGND VPWR VPWR _6936_/X sky130_fd_sc_hd__o22a_1
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9724_ _9769_/CLK _9724_/D _9757_/SET_B VGND VGND VPWR VPWR _9724_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6867_ _9412_/Q VGND VGND VPWR VPWR _6867_/Y sky130_fd_sc_hd__clkinv_2
X_9655_ _9655_/CLK _9655_/D _9779_/SET_B VGND VGND VPWR VPWR _9655_/Q sky130_fd_sc_hd__dfrtp_1
X_8606_ _8672_/B _8606_/B VGND VGND VPWR VPWR _8705_/B sky130_fd_sc_hd__or2_1
X_5818_ _6052_/A _5818_/B VGND VGND VPWR VPWR _5819_/A sky130_fd_sc_hd__or2_1
X_9586_ _8837_/A1 _9586_/D _5190_/X VGND VGND VPWR VPWR _9586_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6798_ _6793_/Y _5534_/B _6794_/Y _4907_/X _6797_/X VGND VGND VPWR VPWR _6830_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_148_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5749_ _9240_/Q _5744_/A _8839_/X _5744_/Y VGND VGND VPWR VPWR _9240_/D sky130_fd_sc_hd__a22o_1
X_8537_ _7836_/A _8299_/B _8061_/C _8536_/Y _8474_/B VGND VGND VPWR VPWR _8617_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_182_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8468_ _8468_/A _8630_/A VGND VGND VPWR VPWR _8470_/B sky130_fd_sc_hd__or2_1
XFILLER_135_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8399_ _8213_/A _8117_/B _8395_/X _8398_/Y VGND VGND VPWR VPWR _8399_/X sky130_fd_sc_hd__o211a_1
X_7419_ _7419_/A VGND VGND VPWR VPWR _7419_/X sky130_fd_sc_hd__buf_6
XFILLER_150_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput180 wb_dat_i[23] VGND VGND VPWR VPWR _7750_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_95_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput191 wb_dat_i[4] VGND VGND VPWR VPWR _8965_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7770_ _7770_/A _7770_/B VGND VGND VPWR VPWR _7775_/B sky130_fd_sc_hd__nand2_1
X_4982_ _9702_/Q _4966_/A _9701_/Q _4966_/Y VGND VGND VPWR VPWR _9702_/D sky130_fd_sc_hd__a22o_1
XFILLER_189_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6721_ _6719_/Y _5450_/B _6720_/Y _5431_/B VGND VGND VPWR VPWR _6721_/X sky130_fd_sc_hd__o22a_1
XFILLER_189_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9440_ _9440_/CLK _9440_/D _4628_/A VGND VGND VPWR VPWR _9440_/Q sky130_fd_sc_hd__dfrtp_1
X_6652_ _9775_/Q VGND VGND VPWR VPWR _6652_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_31_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9371_ _9371_/CLK _9371_/D _9295_/SET_B VGND VGND VPWR VPWR _9371_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_149_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5603_ _5603_/A VGND VGND VPWR VPWR _5604_/A sky130_fd_sc_hd__clkbuf_2
X_6583_ _9357_/Q VGND VGND VPWR VPWR _6583_/Y sky130_fd_sc_hd__clkinv_4
X_8322_ _7862_/Y _8302_/Y _8318_/X _8493_/C _8657_/A VGND VGND VPWR VPWR _8327_/A
+ sky130_fd_sc_hd__a2111o_2
X_5534_ _5545_/A _5534_/B VGND VGND VPWR VPWR _5535_/A sky130_fd_sc_hd__or2_1
XFILLER_145_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5465_ _9401_/Q _5460_/A _5964_/B1 _5460_/Y VGND VGND VPWR VPWR _9401_/D sky130_fd_sc_hd__a22o_1
X_8253_ _8253_/A _8577_/B VGND VGND VPWR VPWR _8255_/A sky130_fd_sc_hd__or2_1
XFILLER_160_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8184_ _8184_/A _8636_/B VGND VGND VPWR VPWR _8295_/A sky130_fd_sc_hd__or2_1
XFILLER_132_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7204_ _6353_/Y _7048_/B _6462_/Y _7077_/A _7203_/X VGND VGND VPWR VPWR _7211_/A
+ sky130_fd_sc_hd__o221a_1
X_7135_ _6891_/Y _7077_/C _6916_/Y _7077_/D _7134_/X VGND VGND VPWR VPWR _7135_/X
+ sky130_fd_sc_hd__o221a_1
X_5396_ _9449_/Q _5395_/A _8846_/X _5395_/Y VGND VGND VPWR VPWR _9449_/D sky130_fd_sc_hd__a22o_1
XFILLER_160_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7066_ _9246_/Q _9245_/Q _7098_/C _7073_/C VGND VGND VPWR VPWR _7067_/A sky130_fd_sc_hd__or4_1
XFILLER_59_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6017_ _9082_/Q _5995_/A _8902_/X _5995_/Y VGND VGND VPWR VPWR _9082_/D sky130_fd_sc_hd__a22o_1
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7968_ _7968_/A _8218_/A VGND VGND VPWR VPWR _8120_/B sky130_fd_sc_hd__or2_1
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9707_ _4446_/A1 _9707_/D _4963_/X VGND VGND VPWR VPWR _9707_/Q sky130_fd_sc_hd__dfrtp_1
X_7899_ _7899_/A _8525_/C VGND VGND VPWR VPWR _8472_/A sky130_fd_sc_hd__or2_2
X_6919_ _9107_/Q VGND VGND VPWR VPWR _6919_/Y sky130_fd_sc_hd__clkinv_2
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9638_ _9639_/CLK _9638_/D _9633_/SET_B VGND VGND VPWR VPWR _9638_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_183_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9569_ _8837_/A1 _9569_/D _5213_/X VGND VGND VPWR VPWR _9569_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_136_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5250_ _9546_/Q _5242_/A _5967_/B1 _5242_/Y VGND VGND VPWR VPWR _9546_/D sky130_fd_sc_hd__a22o_1
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5181_ _9593_/Q _5180_/A _8844_/X _5180_/Y VGND VGND VPWR VPWR _9593_/D sky130_fd_sc_hd__a22o_1
XFILLER_142_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8940_ _9088_/Q _9087_/Q _9051_/Q VGND VGND VPWR VPWR _8940_/X sky130_fd_sc_hd__mux2_1
X_8871_ _8870_/X _9174_/Q _9054_/Q VGND VGND VPWR VPWR _8871_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7822_ _8202_/A _8272_/A VGND VGND VPWR VPWR _8703_/A sky130_fd_sc_hd__nor2_4
XFILLER_36_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7753_ _8394_/C _7839_/A VGND VGND VPWR VPWR _7838_/B sky130_fd_sc_hd__or2_2
X_4965_ _4965_/A VGND VGND VPWR VPWR _4966_/A sky130_fd_sc_hd__buf_8
XFILLER_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6704_ _9470_/Q VGND VGND VPWR VPWR _6704_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9423_ _9684_/CLK _9423_/D _9685_/SET_B VGND VGND VPWR VPWR _9423_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_177_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7684_ _6373_/Y _7415_/X _6416_/Y _7417_/X _7683_/X VGND VGND VPWR VPWR _7698_/B
+ sky130_fd_sc_hd__o221a_1
X_4896_ _4896_/A _4896_/B _4896_/C _4896_/D VGND VGND VPWR VPWR _4935_/C sky130_fd_sc_hd__and4_1
XFILLER_165_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6635_ _6633_/Y _5660_/B _6634_/Y _5671_/B VGND VGND VPWR VPWR _6635_/X sky130_fd_sc_hd__o22a_1
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9354_ _9354_/CLK _9354_/D _9685_/SET_B VGND VGND VPWR VPWR _9354_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6566_ _6561_/Y _4832_/X _8791_/A _5355_/B _6565_/X VGND VGND VPWR VPWR _6567_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_192_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9285_ _9687_/CLK _9285_/D _9528_/SET_B VGND VGND VPWR VPWR _9285_/Q sky130_fd_sc_hd__dfrtp_1
X_5517_ _9364_/Q _5509_/A _8839_/X _5509_/Y VGND VGND VPWR VPWR _9364_/D sky130_fd_sc_hd__a22o_1
XFILLER_152_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8305_ _8305_/A _8305_/B VGND VGND VPWR VPWR _8447_/B sky130_fd_sc_hd__or2_1
X_6497_ _9243_/Q VGND VGND VPWR VPWR _6497_/Y sky130_fd_sc_hd__clkinv_2
X_8236_ _8236_/A VGND VGND VPWR VPWR _8359_/B sky130_fd_sc_hd__inv_2
XFILLER_172_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5448_ _9412_/Q _5444_/A _5966_/B1 _5444_/Y VGND VGND VPWR VPWR _9412_/D sky130_fd_sc_hd__a22o_1
X_5379_ _9460_/Q _5376_/A _8841_/X _5376_/Y VGND VGND VPWR VPWR _9460_/D sky130_fd_sc_hd__a22o_1
X_8167_ _8167_/A _8715_/A VGND VGND VPWR VPWR _8172_/A sky130_fd_sc_hd__or2_1
XFILLER_87_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8098_ _8098_/A _8098_/B VGND VGND VPWR VPWR _8688_/A sky130_fd_sc_hd__nor2_1
XFILLER_99_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7118_ _7118_/A VGND VGND VPWR VPWR _7118_/X sky130_fd_sc_hd__buf_8
XFILLER_86_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7049_ _7098_/C _7125_/A _7073_/C VGND VGND VPWR VPWR _7050_/A sky130_fd_sc_hd__or3_1
XFILLER_47_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4750_ _4787_/A _4900_/B VGND VGND VPWR VPWR _5602_/B sky130_fd_sc_hd__or2_4
XFILLER_186_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4681_ _9044_/Q VGND VGND VPWR VPWR _4681_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_146_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6420_ _6415_/Y _5382_/B _6416_/Y _5941_/B _6419_/X VGND VGND VPWR VPWR _6433_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_174_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6351_ _6346_/Y _5267_/B _6347_/Y _5328_/B _6350_/X VGND VGND VPWR VPWR _6352_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_161_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5302_ _9513_/Q _5300_/A _5964_/B1 _5300_/Y VGND VGND VPWR VPWR _9513_/D sky130_fd_sc_hd__a22o_1
X_9070_ _9687_/CLK _9070_/D _9685_/SET_B VGND VGND VPWR VPWR _9070_/Q sky130_fd_sc_hd__dfstp_1
X_6282_ _9672_/Q VGND VGND VPWR VPWR _6282_/Y sky130_fd_sc_hd__clkinv_2
X_8021_ _8521_/A _8130_/B VGND VGND VPWR VPWR _8403_/A sky130_fd_sc_hd__or2_1
X_5233_ _5233_/A VGND VGND VPWR VPWR _5234_/A sky130_fd_sc_hd__clkbuf_2
X_5164_ _9604_/Q _5158_/A _8841_/X _5158_/Y VGND VGND VPWR VPWR _9604_/D sky130_fd_sc_hd__a22o_1
XFILLER_124_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_opt_3_0_csclk clkbuf_2_1_0_csclk/X VGND VGND VPWR VPWR clkbuf_opt_3_0_csclk/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_96_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5095_ _9650_/Q _5091_/A _8925_/A1 _5091_/Y VGND VGND VPWR VPWR _9650_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8923_ _9621_/Q _8929_/A1 _8955_/S VGND VGND VPWR VPWR _8923_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8854_ _7536_/Y _9635_/Q _8978_/S VGND VGND VPWR VPWR _8854_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7805_ _7839_/A _8632_/A VGND VGND VPWR VPWR _7806_/A sky130_fd_sc_hd__or2_1
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8785_ _8785_/A VGND VGND VPWR VPWR _8786_/A sky130_fd_sc_hd__clkbuf_1
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5997_ _6040_/A VGND VGND VPWR VPWR _5998_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_52_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7736_ _9066_/Q _7736_/B VGND VGND VPWR VPWR _7736_/X sky130_fd_sc_hd__and2_1
X_4948_ _4948_/A VGND VGND VPWR VPWR _4948_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_177_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7667_ _6543_/Y _7427_/X _6484_/Y _5699_/X VGND VGND VPWR VPWR _7667_/X sky130_fd_sc_hd__o22a_1
X_4879_ _9771_/Q VGND VGND VPWR VPWR _4879_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6618_ _6618_/A VGND VGND VPWR VPWR _6618_/Y sky130_fd_sc_hd__inv_2
X_9406_ _9493_/CLK _9406_/D _4628_/A VGND VGND VPWR VPWR _9406_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7598_ _6127_/Y _7425_/X _7595_/X _7597_/X VGND VGND VPWR VPWR _7608_/C sky130_fd_sc_hd__o211a_1
X_9337_ _9532_/CLK _9337_/D _9528_/SET_B VGND VGND VPWR VPWR _9337_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_152_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6549_ _9776_/Q VGND VGND VPWR VPWR _6549_/Y sky130_fd_sc_hd__inv_2
X_9268_ _9354_/CLK _9268_/D _9685_/SET_B VGND VGND VPWR VPWR _9268_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8219_ _8279_/C _8311_/B VGND VGND VPWR VPWR _8219_/Y sky130_fd_sc_hd__nor2_1
XFILLER_160_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9199_ _9789_/CLK _9199_/D _4628_/A VGND VGND VPWR VPWR _9199_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput270 _9725_/Q VGND VGND VPWR VPWR pll_div[4] sky130_fd_sc_hd__buf_2
Xoutput281 _9747_/Q VGND VGND VPWR VPWR pll_trim[15] sky130_fd_sc_hd__buf_2
Xoutput292 _9757_/Q VGND VGND VPWR VPWR pll_trim[25] sky130_fd_sc_hd__buf_2
XFILLER_58_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5920_ _9123_/Q _5918_/A _5964_/B1 _5918_/Y VGND VGND VPWR VPWR _9123_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5851_ _5849_/X _8871_/X _8924_/X _9175_/Q VGND VGND VPWR VPWR _9175_/D sky130_fd_sc_hd__o22a_1
X_8570_ _8213_/A _8117_/A _8341_/B _8260_/B _8352_/B VGND VGND VPWR VPWR _8572_/C
+ sky130_fd_sc_hd__o221ai_4
X_5782_ _9222_/Q _5778_/A _8925_/A1 _5778_/Y VGND VGND VPWR VPWR _9222_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4802_ _4802_/A VGND VGND VPWR VPWR _4931_/B sky130_fd_sc_hd__buf_6
XFILLER_166_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4733_ _4787_/A _4917_/A VGND VGND VPWR VPWR _5621_/B sky130_fd_sc_hd__or2_4
X_7521_ _8743_/A _7419_/X _8781_/A _7421_/X VGND VGND VPWR VPWR _7521_/X sky130_fd_sc_hd__o22a_1
X_7452_ _7466_/A _7470_/B _7474_/D VGND VGND VPWR VPWR _7453_/A sky130_fd_sc_hd__or3_1
XFILLER_9_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4664_ _9125_/Q VGND VGND VPWR VPWR _4664_/Y sky130_fd_sc_hd__clkinv_2
X_6403_ _9782_/Q VGND VGND VPWR VPWR _6403_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7383_ _6417_/Y _7079_/B _6379_/Y _7059_/A VGND VGND VPWR VPWR _7383_/X sky130_fd_sc_hd__o22a_1
X_4595_ _9737_/Q _4592_/A _8844_/X _4592_/Y VGND VGND VPWR VPWR _9737_/D sky130_fd_sc_hd__a22o_1
X_6334_ _9097_/Q VGND VGND VPWR VPWR _6334_/Y sky130_fd_sc_hd__inv_2
X_9122_ _9785_/CLK _9122_/D _7011_/B VGND VGND VPWR VPWR _9122_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_130_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6265_ _9731_/Q VGND VGND VPWR VPWR _6265_/Y sky130_fd_sc_hd__inv_2
X_9053_ _9279_/CLK _9053_/D _9633_/SET_B VGND VGND VPWR VPWR _9053_/Q sky130_fd_sc_hd__dfstp_1
X_8004_ _8394_/D _8164_/A VGND VGND VPWR VPWR _8005_/A sky130_fd_sc_hd__or2_1
XFILLER_135_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5216_ _9569_/Q _5214_/Y _5985_/B _5215_/Y VGND VGND VPWR VPWR _9569_/D sky130_fd_sc_hd__o22a_1
X_6196_ _9482_/Q VGND VGND VPWR VPWR _6196_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5147_ _5147_/A VGND VGND VPWR VPWR _5147_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5078_ _8961_/X _9659_/Q _5078_/S VGND VGND VPWR VPWR _5079_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8906_ _9614_/Q _8925_/A1 _8930_/S VGND VGND VPWR VPWR _8906_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8837_ input83/X _8837_/A1 _9586_/Q VGND VGND VPWR VPWR _8837_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8768_ _8768_/A VGND VGND VPWR VPWR _8768_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_178_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7719_ _9087_/Q _7719_/B VGND VGND VPWR VPWR _7721_/A sky130_fd_sc_hd__nand2_1
XFILLER_138_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8699_ _8699_/A _8699_/B _8699_/C _8699_/D VGND VGND VPWR VPWR _8732_/A sky130_fd_sc_hd__or4_1
XFILLER_180_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6050_ _6050_/A VGND VGND VPWR VPWR _6051_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_112_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5001_ _8908_/X _9698_/Q _5001_/S VGND VGND VPWR VPWR _5002_/A sky130_fd_sc_hd__mux2_1
X_6952_ _6952_/A VGND VGND VPWR VPWR _6952_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_81_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9740_ _9777_/CLK _9740_/D _9757_/SET_B VGND VGND VPWR VPWR _9740_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_38_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5903_ _9134_/Q _5899_/A _5966_/B1 _5899_/Y VGND VGND VPWR VPWR _9134_/D sky130_fd_sc_hd__a22o_1
X_6883_ _9186_/Q VGND VGND VPWR VPWR _6883_/Y sky130_fd_sc_hd__inv_2
X_9671_ _9674_/CLK _9671_/D _9633_/SET_B VGND VGND VPWR VPWR _9671_/Q sky130_fd_sc_hd__dfrtp_1
X_8622_ _7971_/A _8116_/B _8624_/B _8397_/A _8395_/B VGND VGND VPWR VPWR _8622_/X
+ sky130_fd_sc_hd__o311a_1
X_5834_ _9187_/Q _5831_/A _5965_/B1 _5831_/Y VGND VGND VPWR VPWR _9187_/D sky130_fd_sc_hd__a22o_1
XFILLER_22_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5765_ _9233_/Q _5759_/A _8841_/X _5759_/Y VGND VGND VPWR VPWR _9233_/D sky130_fd_sc_hd__a22o_1
X_8553_ _8553_/A _8627_/D _8686_/C _8630_/D VGND VGND VPWR VPWR _8559_/A sky130_fd_sc_hd__or4_2
XFILLER_22_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8484_ _8188_/B _8389_/A _8086_/B VGND VGND VPWR VPWR _8514_/C sky130_fd_sc_hd__o21ai_1
XFILLER_147_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4716_ _9177_/Q VGND VGND VPWR VPWR _4716_/Y sky130_fd_sc_hd__clkinv_2
X_7504_ _6639_/Y _7415_/X _6681_/Y _7417_/X _7503_/X VGND VGND VPWR VPWR _7518_/B
+ sky130_fd_sc_hd__o221a_1
X_5696_ _5724_/B _7462_/A _7456_/A VGND VGND VPWR VPWR _5696_/Y sky130_fd_sc_hd__nor3_1
X_4647_ _4994_/A VGND VGND VPWR VPWR _4648_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_30_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7435_ _7472_/A _7470_/B _7474_/D VGND VGND VPWR VPWR _7436_/A sky130_fd_sc_hd__or3_1
XFILLER_162_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7366_ _6484_/Y _7112_/X _6528_/Y _7077_/B VGND VGND VPWR VPWR _7366_/X sky130_fd_sc_hd__o22a_1
XFILLER_162_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6317_ _6317_/A VGND VGND VPWR VPWR _6317_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4578_ _4578_/A VGND VGND VPWR VPWR _4579_/A sky130_fd_sc_hd__clkbuf_4
X_9105_ _9777_/CLK _9105_/D _7011_/B VGND VGND VPWR VPWR _9105_/Q sky130_fd_sc_hd__dfrtp_1
X_7297_ _4712_/Y _7068_/A _4836_/Y _7105_/X VGND VGND VPWR VPWR _7297_/X sky130_fd_sc_hd__o22a_1
X_9036_ _9664_/CLK _9036_/D VGND VGND VPWR VPWR _9036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6248_ _6243_/Y _4577_/B _6244_/Y _5317_/B _6247_/X VGND VGND VPWR VPWR _6248_/X
+ sky130_fd_sc_hd__o221a_2
X_6179_ _9275_/Q VGND VGND VPWR VPWR _6179_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_103_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5550_ _9343_/Q _5547_/A _8844_/X _5547_/Y VGND VGND VPWR VPWR _9343_/D sky130_fd_sc_hd__a22o_1
XFILLER_157_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5481_ _5481_/A VGND VGND VPWR VPWR _5482_/A sky130_fd_sc_hd__clkbuf_2
X_4501_ _9778_/Q _4493_/A _5967_/B1 _4493_/Y VGND VGND VPWR VPWR _9778_/D sky130_fd_sc_hd__a22o_1
XANTENNA_0 wb_clk_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7220_ _7220_/A _7220_/B _7220_/C _7220_/D VGND VGND VPWR VPWR _7221_/C sky130_fd_sc_hd__and4_1
XFILLER_6_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7151_ _6818_/Y _5728_/X _6913_/Y _7040_/A _7150_/X VGND VGND VPWR VPWR _7154_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6102_ _6097_/Y _4832_/X _6098_/Y _5534_/B _6101_/X VGND VGND VPWR VPWR _6119_/A
+ sky130_fd_sc_hd__o221a_2
X_7082_ _7082_/A VGND VGND VPWR VPWR _7082_/X sky130_fd_sc_hd__buf_8
X_6033_ _9074_/Q _6029_/A _8843_/X _6029_/Y VGND VGND VPWR VPWR _9074_/D sky130_fd_sc_hd__a22o_1
XFILLER_140_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7984_ _8525_/A _8091_/B _8098_/A VGND VGND VPWR VPWR _7997_/B sky130_fd_sc_hd__or3_2
XFILLER_94_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6935_ _9227_/Q VGND VGND VPWR VPWR _6935_/Y sky130_fd_sc_hd__inv_2
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9723_ _9769_/CLK _9723_/D _9757_/SET_B VGND VGND VPWR VPWR _9723_/Q sky130_fd_sc_hd__dfstp_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6866_ _9464_/Q VGND VGND VPWR VPWR _6866_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_22_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9654_ _9779_/CLK _9654_/D _9779_/SET_B VGND VGND VPWR VPWR _9654_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_179_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8605_ _8605_/A _8605_/B VGND VGND VPWR VPWR _8707_/B sky130_fd_sc_hd__or2_1
X_5817_ _9198_/Q _5812_/A _8839_/X _5812_/Y VGND VGND VPWR VPWR _9198_/D sky130_fd_sc_hd__a22o_1
X_6797_ _6795_/Y _4537_/B _6796_/Y _4564_/B VGND VGND VPWR VPWR _6797_/X sky130_fd_sc_hd__o22a_2
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9585_ _9674_/CLK _9585_/D _9633_/SET_B VGND VGND VPWR VPWR _9585_/Q sky130_fd_sc_hd__dfrtp_2
X_5748_ _9241_/Q _5744_/A _8930_/A1 _5744_/Y VGND VGND VPWR VPWR _9241_/D sky130_fd_sc_hd__a22o_1
X_8536_ _8536_/A VGND VGND VPWR VPWR _8536_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5679_ _6052_/A _5679_/B VGND VGND VPWR VPWR _5680_/A sky130_fd_sc_hd__or2_1
XFILLER_135_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8467_ _8467_/A VGND VGND VPWR VPWR _8630_/A sky130_fd_sc_hd__inv_2
X_8398_ _8396_/Y _8397_/Y _8121_/Y VGND VGND VPWR VPWR _8398_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_123_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7418_ _7476_/A _9251_/Q _7456_/A _9255_/Q VGND VGND VPWR VPWR _7419_/A sky130_fd_sc_hd__or4_1
XFILLER_116_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7349_ _6712_/Y _5728_/X _6685_/Y _7040_/A _7348_/X VGND VGND VPWR VPWR _7352_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_173_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9019_ _9039_/CLK _9019_/D VGND VGND VPWR VPWR _9019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput181 wb_dat_i[24] VGND VGND VPWR VPWR _7737_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput170 wb_dat_i[14] VGND VGND VPWR VPWR _7749_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_95_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput192 wb_dat_i[5] VGND VGND VPWR VPWR _8966_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4981_ _4981_/A VGND VGND VPWR VPWR _4981_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_91_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6720_ _9418_/Q VGND VGND VPWR VPWR _6720_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6651_ _9728_/Q VGND VGND VPWR VPWR _6651_/Y sky130_fd_sc_hd__inv_2
X_6582_ _9289_/Q VGND VGND VPWR VPWR _6582_/Y sky130_fd_sc_hd__inv_2
X_9370_ _9371_/CLK _9370_/D _9295_/SET_B VGND VGND VPWR VPWR _9370_/Q sky130_fd_sc_hd__dfrtp_1
X_5602_ _5671_/A _5602_/B VGND VGND VPWR VPWR _5603_/A sky130_fd_sc_hd__or2_1
XFILLER_31_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5533_ _9354_/Q _5528_/A _8839_/X _5528_/Y VGND VGND VPWR VPWR _9354_/D sky130_fd_sc_hd__a22o_1
X_8321_ _8461_/A _8674_/B VGND VGND VPWR VPWR _8657_/A sky130_fd_sc_hd__or2_1
X_8252_ _8319_/A _8260_/B VGND VGND VPWR VPWR _8577_/B sky130_fd_sc_hd__nor2_1
X_5464_ _9402_/Q _5460_/A _5963_/B1 _5460_/Y VGND VGND VPWR VPWR _9402_/D sky130_fd_sc_hd__a22o_1
X_8183_ _8096_/A _8386_/A _8097_/B _9066_/Q VGND VGND VPWR VPWR _8636_/B sky130_fd_sc_hd__o31ai_4
XFILLER_132_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7203_ _6463_/Y _7040_/C _6337_/Y _7059_/C VGND VGND VPWR VPWR _7203_/X sky130_fd_sc_hd__o22a_1
X_5395_ _5395_/A VGND VGND VPWR VPWR _5395_/Y sky130_fd_sc_hd__inv_2
XFILLER_160_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7134_ _6853_/Y _7086_/X _6855_/Y _7088_/X VGND VGND VPWR VPWR _7134_/X sky130_fd_sc_hd__o22a_1
XFILLER_86_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7065_ _7065_/A VGND VGND VPWR VPWR _7068_/C sky130_fd_sc_hd__buf_8
X_6016_ _6016_/A VGND VGND VPWR VPWR _6016_/X sky130_fd_sc_hd__clkbuf_1
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7967_ _7756_/B _8102_/B _7756_/B _8102_/B VGND VGND VPWR VPWR _7968_/A sky130_fd_sc_hd__o2bb2a_1
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9706_ _4446_/A1 _9706_/D _4969_/X VGND VGND VPWR VPWR _9706_/Q sky130_fd_sc_hd__dfrtp_1
X_7898_ _8008_/C _7898_/B VGND VGND VPWR VPWR _8525_/C sky130_fd_sc_hd__or2_4
XFILLER_168_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6918_ _6913_/Y _5968_/B _6914_/Y _5621_/B _6917_/X VGND VGND VPWR VPWR _6925_/C
+ sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_13_csclk clkbuf_2_2_0_csclk/X VGND VGND VPWR VPWR _9532_/CLK sky130_fd_sc_hd__clkbuf_16
X_6849_ _6849_/A VGND VGND VPWR VPWR _6849_/Y sky130_fd_sc_hd__inv_2
X_9637_ _9791_/CLK _9637_/D _9633_/SET_B VGND VGND VPWR VPWR _9637_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_52_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9568_ _9617_/CLK _9568_/D _9295_/SET_B VGND VGND VPWR VPWR _9568_/Q sky130_fd_sc_hd__dfrtp_2
X_9499_ _9501_/CLK _9499_/D _9647_/SET_B VGND VGND VPWR VPWR _9499_/Q sky130_fd_sc_hd__dfrtp_1
X_8519_ _8516_/Y _8517_/Y _8518_/X _8453_/C VGND VGND VPWR VPWR _8607_/A sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_28_csclk clkbuf_opt_6_0_csclk/X VGND VGND VPWR VPWR _9378_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_190_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5180_ _5180_/A VGND VGND VPWR VPWR _5180_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_96_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8870_ _7680_/Y _9630_/Q _8978_/S VGND VGND VPWR VPWR _8870_/X sky130_fd_sc_hd__mux2_1
X_7821_ _8394_/A _8394_/B _7838_/B VGND VGND VPWR VPWR _8272_/A sky130_fd_sc_hd__or3_4
X_7752_ _8379_/B VGND VGND VPWR VPWR _8394_/B sky130_fd_sc_hd__inv_2
X_4964_ _9048_/Q _4964_/B _9051_/Q VGND VGND VPWR VPWR _4965_/A sky130_fd_sc_hd__or3_1
XFILLER_36_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6703_ _6698_/Y _6251_/A _6699_/Y _4577_/B _6702_/X VGND VGND VPWR VPWR _6716_/B
+ sky130_fd_sc_hd__o221a_4
XFILLER_51_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9422_ _9684_/CLK _9422_/D _9685_/SET_B VGND VGND VPWR VPWR _9422_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_177_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4895_ _4887_/Y _4590_/B _4888_/Y _5298_/B _4894_/X VGND VGND VPWR VPWR _4896_/D
+ sky130_fd_sc_hd__o221a_1
X_7683_ _6464_/Y _7419_/X _6341_/Y _7421_/X VGND VGND VPWR VPWR _7683_/X sky130_fd_sc_hd__o22a_1
XFILLER_149_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6634_ _9266_/Q VGND VGND VPWR VPWR _6634_/Y sky130_fd_sc_hd__clkinv_2
X_9353_ _9378_/CLK _9353_/D _9646_/SET_B VGND VGND VPWR VPWR _9353_/Q sky130_fd_sc_hd__dfrtp_1
X_6565_ _8783_/A _6027_/B _6564_/Y _4861_/X VGND VGND VPWR VPWR _6565_/X sky130_fd_sc_hd__o22a_1
X_9284_ _9358_/CLK _9284_/D _9528_/SET_B VGND VGND VPWR VPWR _9284_/Q sky130_fd_sc_hd__dfrtp_1
X_5516_ _9365_/Q _5509_/A _8930_/A1 _5509_/Y VGND VGND VPWR VPWR _9365_/D sky130_fd_sc_hd__a22o_1
X_6496_ _9128_/Q VGND VGND VPWR VPWR _7701_/A sky130_fd_sc_hd__clkinv_4
X_8304_ _8451_/A _8642_/B VGND VGND VPWR VPWR _8304_/Y sky130_fd_sc_hd__nor2_1
XFILLER_160_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5447_ _9413_/Q _5444_/A _5965_/B1 _5444_/Y VGND VGND VPWR VPWR _9413_/D sky130_fd_sc_hd__a22o_1
X_8235_ _8510_/A _8239_/B VGND VGND VPWR VPWR _8236_/A sky130_fd_sc_hd__or2_1
XFILLER_154_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5378_ _9461_/Q _5376_/A _8842_/X _5376_/Y VGND VGND VPWR VPWR _9461_/D sky130_fd_sc_hd__a22o_1
XFILLER_120_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8166_ _8168_/A _8640_/B VGND VGND VPWR VPWR _8715_/A sky130_fd_sc_hd__nor2_1
X_8097_ _8170_/A _8097_/B VGND VGND VPWR VPWR _8098_/B sky130_fd_sc_hd__or2_1
X_7117_ _9246_/Q _9245_/Q _7127_/B _7127_/C VGND VGND VPWR VPWR _7118_/A sky130_fd_sc_hd__or4_1
X_7048_ _7392_/B _7048_/B _7048_/C _7048_/D VGND VGND VPWR VPWR _7078_/A sky130_fd_sc_hd__and4_1
XFILLER_47_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8999_ _9567_/Q _8775_/A VGND VGND VPWR VPWR mgmt_gpio_out[22] sky130_fd_sc_hd__ebufn_8
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4680_ _5178_/B VGND VGND VPWR VPWR _4680_/Y sky130_fd_sc_hd__inv_4
XFILLER_186_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6350_ _6348_/Y _5404_/B _6349_/Y _5278_/B VGND VGND VPWR VPWR _6350_/X sky130_fd_sc_hd__o22a_1
XFILLER_154_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5301_ _9514_/Q _5300_/A _5963_/B1 _5300_/Y VGND VGND VPWR VPWR _9514_/D sky130_fd_sc_hd__a22o_1
XFILLER_142_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6281_ _8801_/A VGND VGND VPWR VPWR _6281_/Y sky130_fd_sc_hd__inv_2
X_8020_ _8401_/A _8389_/A _8097_/B _8401_/A _8019_/X VGND VGND VPWR VPWR _8020_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_69_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5232_ _5259_/A _5232_/B VGND VGND VPWR VPWR _5233_/A sky130_fd_sc_hd__or2_1
X_5163_ _9605_/Q _5158_/A _8842_/X _5158_/Y VGND VGND VPWR VPWR _9605_/D sky130_fd_sc_hd__a22o_1
XFILLER_124_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5094_ _9651_/Q _5091_/A _8844_/X _5091_/Y VGND VGND VPWR VPWR _9651_/D sky130_fd_sc_hd__a22o_1
XFILLER_96_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8922_ _9604_/Q _8841_/X _8926_/S VGND VGND VPWR VPWR _8922_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8853_ _8852_/X _9165_/Q _9054_/Q VGND VGND VPWR VPWR _8853_/X sky130_fd_sc_hd__mux2_1
X_7804_ _8379_/C _8394_/A _8379_/B VGND VGND VPWR VPWR _8632_/A sky130_fd_sc_hd__or3_4
XFILLER_64_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8784_ _8784_/A VGND VGND VPWR VPWR _8784_/X sky130_fd_sc_hd__clkbuf_1
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5996_ _9089_/Q _5995_/A _8907_/X _5995_/Y VGND VGND VPWR VPWR _9089_/D sky130_fd_sc_hd__a22o_1
XFILLER_52_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7735_ _9067_/Q _5058_/X _7733_/X _7734_/X VGND VGND VPWR VPWR _7735_/X sky130_fd_sc_hd__a211o_1
X_4947_ _4994_/A VGND VGND VPWR VPWR _4948_/A sky130_fd_sc_hd__clkbuf_1
X_4878_ _6158_/B _4931_/B VGND VGND VPWR VPWR _5496_/B sky130_fd_sc_hd__or2_4
X_7666_ _6581_/Y _7415_/X _6539_/Y _7417_/X _7665_/X VGND VGND VPWR VPWR _7680_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_177_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6617_ _9630_/Q VGND VGND VPWR VPWR _6617_/Y sky130_fd_sc_hd__inv_2
X_9405_ _9758_/CLK _9405_/D _7011_/B VGND VGND VPWR VPWR _9405_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9336_ _9532_/CLK _9336_/D _9647_/SET_B VGND VGND VPWR VPWR _9336_/Q sky130_fd_sc_hd__dfrtp_1
X_7597_ _6123_/Y _7430_/X _6083_/Y _7432_/X _7596_/X VGND VGND VPWR VPWR _7597_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_118_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6548_ _6543_/Y _5374_/B _6544_/Y _5110_/B _6547_/X VGND VGND VPWR VPWR _6567_/A
+ sky130_fd_sc_hd__o221a_1
X_9267_ _9354_/CLK _9267_/D _9685_/SET_B VGND VGND VPWR VPWR _9267_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6479_ _9123_/Q VGND VGND VPWR VPWR _6479_/Y sky130_fd_sc_hd__inv_2
X_8218_ _8218_/A _8218_/B _8218_/C VGND VGND VPWR VPWR _8279_/C sky130_fd_sc_hd__or3_2
X_9198_ _9440_/CLK _9198_/D _4628_/A VGND VGND VPWR VPWR _9198_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput271 _9719_/Q VGND VGND VPWR VPWR pll_ena sky130_fd_sc_hd__buf_2
Xoutput260 _7017_/A VGND VGND VPWR VPWR pad_flash_io1_oeb sky130_fd_sc_hd__buf_2
XFILLER_160_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8149_ _8164_/A _8552_/A VGND VGND VPWR VPWR _8685_/B sky130_fd_sc_hd__nor2_1
Xoutput293 _9734_/Q VGND VGND VPWR VPWR pll_trim[2] sky130_fd_sc_hd__buf_2
Xoutput282 _9748_/Q VGND VGND VPWR VPWR pll_trim[16] sky130_fd_sc_hd__buf_2
XFILLER_58_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5850_ _9176_/Q _8924_/X _8873_/X _5849_/X VGND VGND VPWR VPWR _9176_/D sky130_fd_sc_hd__o22a_1
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5781_ _9223_/Q _5778_/A _8844_/X _5778_/Y VGND VGND VPWR VPWR _9223_/D sky130_fd_sc_hd__a22o_1
X_4801_ _8936_/X _8938_/X _4801_/C VGND VGND VPWR VPWR _4802_/A sky130_fd_sc_hd__or3_1
X_4732_ _9286_/Q VGND VGND VPWR VPWR _4732_/Y sky130_fd_sc_hd__inv_2
X_7520_ _8775_/A _7408_/X _7705_/A _7410_/X _7519_/X VGND VGND VPWR VPWR _7536_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4663_ _4891_/A _4780_/B VGND VGND VPWR VPWR _5556_/B sky130_fd_sc_hd__or2_4
X_7451_ _7451_/A VGND VGND VPWR VPWR _7451_/X sky130_fd_sc_hd__buf_8
XFILLER_147_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6402_ _9550_/Q VGND VGND VPWR VPWR _6402_/Y sky130_fd_sc_hd__inv_2
X_7382_ _6399_/Y _7095_/X _6374_/Y _7068_/D _7381_/X VGND VGND VPWR VPWR _7387_/B
+ sky130_fd_sc_hd__o221a_1
X_4594_ _9738_/Q _4592_/A _8845_/X _4592_/Y VGND VGND VPWR VPWR _9738_/D sky130_fd_sc_hd__a22o_1
X_6333_ _6328_/Y _5458_/B _6329_/Y _5306_/B _6332_/X VGND VGND VPWR VPWR _6352_/A
+ sky130_fd_sc_hd__o221a_1
X_9121_ _9655_/CLK _9121_/D _9779_/SET_B VGND VGND VPWR VPWR _9121_/Q sky130_fd_sc_hd__dfrtp_1
X_6264_ _9421_/Q VGND VGND VPWR VPWR _6264_/Y sky130_fd_sc_hd__inv_6
XFILLER_115_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9052_ _9709_/CLK _9052_/D _6043_/X VGND VGND VPWR VPWR _9052_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8003_ _8009_/A VGND VGND VPWR VPWR _8003_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5215_ _9048_/Q _7008_/A VGND VGND VPWR VPWR _5215_/Y sky130_fd_sc_hd__nor2_1
X_6195_ _9474_/Q VGND VGND VPWR VPWR _6195_/Y sky130_fd_sc_hd__clkinv_2
X_5146_ _5146_/A VGND VGND VPWR VPWR _5147_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_28_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5077_ _5077_/A VGND VGND VPWR VPWR _9660_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8905_ _9612_/Q _8955_/A1 _8930_/S VGND VGND VPWR VPWR _8905_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8836_ input84/X _4629_/C _9626_/Q VGND VGND VPWR VPWR _8836_/X sky130_fd_sc_hd__mux2_2
XFILLER_44_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8767_ _8767_/A VGND VGND VPWR VPWR _8768_/A sky130_fd_sc_hd__clkbuf_1
X_5979_ _6040_/A VGND VGND VPWR VPWR _5980_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_8_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7718_ _7718_/A VGND VGND VPWR VPWR _7719_/B sky130_fd_sc_hd__inv_2
XFILLER_178_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8698_ _8698_/A _8708_/A _7931_/A VGND VGND VPWR VPWR _8699_/B sky130_fd_sc_hd__or3b_1
XFILLER_138_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7649_ _6712_/Y _7427_/X _6632_/Y _5699_/X VGND VGND VPWR VPWR _7649_/X sky130_fd_sc_hd__o22a_2
XFILLER_60_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9319_ _9344_/CLK _9319_/D _9295_/SET_B VGND VGND VPWR VPWR _9319_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_109_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _5000_/A VGND VGND VPWR VPWR _5000_/X sky130_fd_sc_hd__clkbuf_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6951_ _6951_/A VGND VGND VPWR VPWR _6952_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5902_ _9135_/Q _5899_/A _8841_/X _5899_/Y VGND VGND VPWR VPWR _9135_/D sky130_fd_sc_hd__a22o_1
X_6882_ _6879_/Y _5797_/B _7150_/A _5610_/B _6881_/Y VGND VGND VPWR VPWR _6901_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_34_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9670_ _9674_/CLK _9670_/D _9633_/SET_B VGND VGND VPWR VPWR _9670_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_179_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8621_ _8713_/D VGND VGND VPWR VPWR _8621_/Y sky130_fd_sc_hd__inv_2
X_5833_ _9188_/Q _5831_/A _5964_/B1 _5831_/Y VGND VGND VPWR VPWR _9188_/D sky130_fd_sc_hd__a22o_1
XFILLER_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8552_ _8552_/A _8554_/B VGND VGND VPWR VPWR _8630_/D sky130_fd_sc_hd__nor2_1
XFILLER_61_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5764_ _9234_/Q _5759_/A _8929_/A1 _5759_/Y VGND VGND VPWR VPWR _9234_/D sky130_fd_sc_hd__a22o_1
X_7503_ _6667_/Y _7419_/X _6692_/Y _7421_/X VGND VGND VPWR VPWR _7503_/X sky130_fd_sc_hd__o22a_1
X_8483_ _8483_/A _8605_/A VGND VGND VPWR VPWR _8485_/A sky130_fd_sc_hd__or2_1
X_4715_ _4706_/Y _5671_/B _4708_/Y _5776_/B _4714_/X VGND VGND VPWR VPWR _4791_/A
+ sky130_fd_sc_hd__o221a_1
X_5695_ _9254_/Q _9253_/Q VGND VGND VPWR VPWR _7456_/A sky130_fd_sc_hd__or2_4
XFILLER_107_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7434_ _7434_/A VGND VGND VPWR VPWR _7434_/X sky130_fd_sc_hd__buf_6
X_4646_ _9715_/Q _4636_/A _8950_/X _4636_/Y VGND VGND VPWR VPWR _9715_/D sky130_fd_sc_hd__a22o_2
XFILLER_190_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7365_ _7365_/A _7365_/B _7365_/C _7365_/D VGND VGND VPWR VPWR _7375_/B sky130_fd_sc_hd__and4_1
X_4577_ _5960_/A _4577_/B VGND VGND VPWR VPWR _4578_/A sky130_fd_sc_hd__or2_1
XFILLER_190_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6316_ _9274_/Q VGND VGND VPWR VPWR _6316_/Y sky130_fd_sc_hd__clkinv_2
X_9104_ _9775_/CLK _9104_/D _7011_/B VGND VGND VPWR VPWR _9104_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_143_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7296_ _4749_/Y _7059_/B _4890_/Y _7068_/C _7295_/X VGND VGND VPWR VPWR _7299_/C
+ sky130_fd_sc_hd__o221a_2
XFILLER_89_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9035_ _9039_/CLK _9035_/D VGND VGND VPWR VPWR _9035_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6247_ _6245_/Y _4822_/X _6246_/Y _5393_/B VGND VGND VPWR VPWR _6247_/X sky130_fd_sc_hd__o22a_1
X_6178_ _9262_/Q VGND VGND VPWR VPWR _6178_/Y sky130_fd_sc_hd__inv_2
XFILLER_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5129_ _6040_/A VGND VGND VPWR VPWR _5130_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8819_ _9239_/Q _9772_/Q _9787_/Q VGND VGND VPWR VPWR _8819_/X sky130_fd_sc_hd__mux2_4
XFILLER_25_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5480_ _5671_/A _5480_/B VGND VGND VPWR VPWR _5481_/A sky130_fd_sc_hd__or2_1
X_4500_ _9779_/Q _4493_/A _8930_/A1 _4493_/Y VGND VGND VPWR VPWR _9779_/D sky130_fd_sc_hd__a22o_1
XFILLER_172_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_1 _7155_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7150_ _7150_/A _7392_/B VGND VGND VPWR VPWR _7150_/X sky130_fd_sc_hd__or2_1
X_7081_ _7098_/C _7127_/A _7127_/C VGND VGND VPWR VPWR _7082_/A sky130_fd_sc_hd__or3_1
X_6101_ _6099_/Y _4893_/X _6100_/Y _4841_/X VGND VGND VPWR VPWR _6101_/X sky130_fd_sc_hd__o22a_1
X_6032_ _9075_/Q _6029_/A _8844_/X _6029_/Y VGND VGND VPWR VPWR _9075_/D sky130_fd_sc_hd__a22o_1
XFILLER_112_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7983_ _8097_/B VGND VGND VPWR VPWR _8544_/A sky130_fd_sc_hd__clkinv_4
XFILLER_39_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6934_ _9282_/Q VGND VGND VPWR VPWR _7326_/A sky130_fd_sc_hd__clkinv_2
XFILLER_81_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9722_ _9769_/CLK _9722_/D _7011_/B VGND VGND VPWR VPWR _9722_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_19_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9653_ _9653_/CLK _9653_/D _9646_/SET_B VGND VGND VPWR VPWR _9653_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6865_ _9477_/Q VGND VGND VPWR VPWR _6865_/Y sky130_fd_sc_hd__inv_4
X_8604_ _8604_/A VGND VGND VPWR VPWR _8604_/X sky130_fd_sc_hd__clkbuf_1
X_5816_ _9199_/Q _5812_/A _5966_/B1 _5812_/Y VGND VGND VPWR VPWR _9199_/D sky130_fd_sc_hd__a22o_1
X_6796_ _9749_/Q VGND VGND VPWR VPWR _6796_/Y sky130_fd_sc_hd__inv_2
X_9584_ _9674_/CLK _9584_/D _9633_/SET_B VGND VGND VPWR VPWR _9584_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5747_ _9242_/Q _5744_/A _8841_/X _5744_/Y VGND VGND VPWR VPWR _9242_/D sky130_fd_sc_hd__a22o_1
X_8535_ _8535_/A _8668_/C _8615_/D _8699_/A VGND VGND VPWR VPWR _8541_/A sky130_fd_sc_hd__or4_2
XFILLER_10_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8466_ _8466_/A _8615_/C VGND VGND VPWR VPWR _8470_/A sky130_fd_sc_hd__or2_1
XFILLER_41_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5678_ _9264_/Q _5673_/A _8839_/X _5673_/Y VGND VGND VPWR VPWR _9264_/D sky130_fd_sc_hd__a22o_1
X_7417_ _7417_/A VGND VGND VPWR VPWR _7417_/X sky130_fd_sc_hd__buf_6
X_8397_ _8397_/A _8397_/B VGND VGND VPWR VPWR _8397_/Y sky130_fd_sc_hd__nor2_1
XFILLER_123_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4629_ _9789_/Q _9096_/Q _4629_/C VGND VGND VPWR VPWR _7022_/B sky130_fd_sc_hd__or3_4
XFILLER_150_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7348_ _7348_/A _7392_/B VGND VGND VPWR VPWR _7348_/X sky130_fd_sc_hd__or2_1
XFILLER_104_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7279_ _6065_/Y _7040_/D _6098_/Y _7110_/X _7278_/X VGND VGND VPWR VPWR _7286_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_103_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9018_ _9039_/CLK _9018_/D VGND VGND VPWR VPWR _9018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput171 wb_dat_i[15] VGND VGND VPWR VPWR _7751_/B2 sky130_fd_sc_hd__clkbuf_1
Xinput160 wb_adr_i[6] VGND VGND VPWR VPWR _7903_/C sky130_fd_sc_hd__buf_4
XFILLER_83_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput182 wb_dat_i[25] VGND VGND VPWR VPWR _7739_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput193 wb_dat_i[6] VGND VGND VPWR VPWR _8967_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4980_ _4994_/A VGND VGND VPWR VPWR _4981_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_91_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6650_ _9072_/Q VGND VGND VPWR VPWR _6650_/Y sky130_fd_sc_hd__inv_4
XFILLER_149_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5601_ _9307_/Q _5596_/A _8839_/X _5596_/Y VGND VGND VPWR VPWR _9307_/D sky130_fd_sc_hd__a22o_1
XFILLER_31_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6581_ _9215_/Q VGND VGND VPWR VPWR _6581_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5532_ _9355_/Q _5528_/A _5966_/B1 _5528_/Y VGND VGND VPWR VPWR _9355_/D sky130_fd_sc_hd__a22o_1
X_8320_ _8320_/A VGND VGND VPWR VPWR _8461_/A sky130_fd_sc_hd__inv_2
XFILLER_117_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_9_csclk clkbuf_2_2_0_csclk/X VGND VGND VPWR VPWR _9687_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_172_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5463_ _9403_/Q _5460_/A _8844_/X _5460_/Y VGND VGND VPWR VPWR _9403_/D sky130_fd_sc_hd__a22o_1
X_8251_ _8251_/A _8597_/B VGND VGND VPWR VPWR _8253_/A sky130_fd_sc_hd__or2_1
X_8182_ _8433_/B _8182_/B VGND VGND VPWR VPWR _8184_/A sky130_fd_sc_hd__nor2_1
XFILLER_132_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7202_ _6427_/Y _7082_/X _6390_/Y _7084_/X _7201_/X VGND VGND VPWR VPWR _7221_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_99_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5394_ _5394_/A VGND VGND VPWR VPWR _5395_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_132_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7133_ _7133_/A VGND VGND VPWR VPWR _7133_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7064_ _7075_/A _7109_/B VGND VGND VPWR VPWR _7065_/A sky130_fd_sc_hd__or2_1
XFILLER_67_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6015_ _6040_/A VGND VGND VPWR VPWR _6016_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_82_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7966_ _7966_/A _7966_/B _7966_/C VGND VGND VPWR VPWR _8102_/B sky130_fd_sc_hd__or3_1
X_9705_ _4446_/A1 _9705_/D _4972_/X VGND VGND VPWR VPWR _9705_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7897_ _7897_/A VGND VGND VPWR VPWR _8008_/C sky130_fd_sc_hd__inv_2
X_6917_ _6915_/Y _5507_/B _6916_/Y _5545_/B VGND VGND VPWR VPWR _6917_/X sky130_fd_sc_hd__o22a_1
XFILLER_168_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6848_ _9511_/Q VGND VGND VPWR VPWR _6848_/Y sky130_fd_sc_hd__clkinv_2
X_9636_ _9639_/CLK _9636_/D _9633_/SET_B VGND VGND VPWR VPWR _9636_/Q sky130_fd_sc_hd__dfrtp_1
X_9567_ _9617_/CLK _9567_/D _9295_/SET_B VGND VGND VPWR VPWR _9567_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_168_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8518_ _8518_/A _8518_/B VGND VGND VPWR VPWR _8518_/X sky130_fd_sc_hd__or2_4
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6779_ _9517_/Q VGND VGND VPWR VPWR _6779_/Y sky130_fd_sc_hd__inv_2
X_9498_ _9534_/CLK _9498_/D _9647_/SET_B VGND VGND VPWR VPWR _9498_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_151_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8449_ _8449_/A _8449_/B VGND VGND VPWR VPWR _8453_/B sky130_fd_sc_hd__or2_1
XFILLER_123_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7820_ _8660_/B VGND VGND VPWR VPWR _8282_/B sky130_fd_sc_hd__inv_2
XFILLER_64_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7751_ _9068_/Q _7751_/A2 _9067_/Q _7751_/B2 _7750_/X VGND VGND VPWR VPWR _7751_/X
+ sky130_fd_sc_hd__a221o_1
X_4963_ _4963_/A VGND VGND VPWR VPWR _4963_/X sky130_fd_sc_hd__clkbuf_1
X_7682_ _6424_/Y _7400_/X _6362_/Y _7405_/X _7681_/X VGND VGND VPWR VPWR _7698_/A
+ sky130_fd_sc_hd__o221a_1
X_6702_ _6700_/Y _5480_/B _6701_/Y _5564_/B VGND VGND VPWR VPWR _6702_/X sky130_fd_sc_hd__o22a_2
XFILLER_51_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9421_ _9684_/CLK _9421_/D _9528_/SET_B VGND VGND VPWR VPWR _9421_/Q sky130_fd_sc_hd__dfrtp_2
X_6633_ _9271_/Q VGND VGND VPWR VPWR _6633_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_149_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4894_ _4890_/Y _5450_/B _4892_/Y _4893_/X VGND VGND VPWR VPWR _4894_/X sky130_fd_sc_hd__o22a_1
XFILLER_192_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9352_ _9352_/CLK _9352_/D _9646_/SET_B VGND VGND VPWR VPWR _9352_/Q sky130_fd_sc_hd__dfrtp_1
X_6564_ _6564_/A VGND VGND VPWR VPWR _6564_/Y sky130_fd_sc_hd__inv_2
X_9283_ _9687_/CLK _9283_/D _9528_/SET_B VGND VGND VPWR VPWR _9283_/Q sky130_fd_sc_hd__dfstp_1
X_5515_ _9366_/Q _5509_/A _8955_/A1 _5509_/Y VGND VGND VPWR VPWR _9366_/D sky130_fd_sc_hd__a22o_1
X_6495_ _9284_/Q VGND VGND VPWR VPWR _7370_/A sky130_fd_sc_hd__inv_2
X_8303_ _8303_/A VGND VGND VPWR VPWR _8451_/A sky130_fd_sc_hd__inv_2
XFILLER_105_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5446_ _9414_/Q _5444_/A _5964_/B1 _5444_/Y VGND VGND VPWR VPWR _9414_/D sky130_fd_sc_hd__a22o_1
X_8234_ _8238_/A _8264_/B VGND VGND VPWR VPWR _8642_/B sky130_fd_sc_hd__nor2_1
XFILLER_160_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5377_ _9462_/Q _5376_/A _8843_/X _5376_/Y VGND VGND VPWR VPWR _9462_/D sky130_fd_sc_hd__a22o_1
XFILLER_120_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8165_ _8165_/A _8708_/D VGND VGND VPWR VPWR _8167_/A sky130_fd_sc_hd__or2_1
XFILLER_99_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8096_ _8096_/A _8096_/B VGND VGND VPWR VPWR _8170_/A sky130_fd_sc_hd__or2_1
X_7116_ _7116_/A VGND VGND VPWR VPWR _7116_/X sky130_fd_sc_hd__buf_8
X_7047_ _7047_/A VGND VGND VPWR VPWR _7048_/D sky130_fd_sc_hd__clkbuf_16
XFILLER_47_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8998_ _9566_/Q _8773_/A VGND VGND VPWR VPWR mgmt_gpio_out[21] sky130_fd_sc_hd__ebufn_8
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7949_ _8188_/B _8378_/B VGND VGND VPWR VPWR _8185_/A sky130_fd_sc_hd__or2_1
XFILLER_70_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9619_ _9674_/CLK _9619_/D _9633_/SET_B VGND VGND VPWR VPWR _9619_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_183_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5300_ _5300_/A VGND VGND VPWR VPWR _5300_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6280_ _6280_/A _6280_/B _6280_/C _6280_/D VGND VGND VPWR VPWR _6326_/B sky130_fd_sc_hd__and4_2
XFILLER_142_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5231_ _5231_/A VGND VGND VPWR VPWR _9559_/D sky130_fd_sc_hd__clkbuf_1
X_5162_ _9606_/Q _5158_/A _8925_/A1 _5158_/Y VGND VGND VPWR VPWR _9606_/D sky130_fd_sc_hd__a22o_1
XFILLER_123_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_12_csclk clkbuf_2_2_0_csclk/X VGND VGND VPWR VPWR _9535_/CLK sky130_fd_sc_hd__clkbuf_16
X_5093_ _9652_/Q _5091_/A _8845_/X _5091_/Y VGND VGND VPWR VPWR _9652_/D sky130_fd_sc_hd__a22o_1
XFILLER_110_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8921_ _9607_/Q _8844_/X _8926_/S VGND VGND VPWR VPWR _8921_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_27_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR _9352_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8852_ _7518_/Y _9634_/Q _8978_/S VGND VGND VPWR VPWR _8852_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8783_ _8783_/A VGND VGND VPWR VPWR _8784_/A sky130_fd_sc_hd__clkbuf_1
X_7803_ _8188_/B _8624_/B VGND VGND VPWR VPWR _8562_/A sky130_fd_sc_hd__nor2_1
X_7734_ _7734_/A _7734_/B _9068_/Q VGND VGND VPWR VPWR _7734_/X sky130_fd_sc_hd__and3_1
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5995_ _5995_/A VGND VGND VPWR VPWR _5995_/Y sky130_fd_sc_hd__inv_2
X_4946_ _9710_/Q _9696_/Q _9050_/Q _5993_/B VGND VGND VPWR VPWR _9710_/D sky130_fd_sc_hd__o211a_1
XFILLER_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4877_ _9372_/Q VGND VGND VPWR VPWR _4877_/Y sky130_fd_sc_hd__inv_2
X_7665_ _6533_/Y _7419_/X _6609_/Y _7421_/X VGND VGND VPWR VPWR _7665_/X sky130_fd_sc_hd__o22a_1
XFILLER_192_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7596_ _6109_/Y _7434_/X _6110_/Y _7436_/X VGND VGND VPWR VPWR _7596_/X sky130_fd_sc_hd__o22a_1
X_6616_ _9445_/Q VGND VGND VPWR VPWR _8793_/A sky130_fd_sc_hd__clkinv_8
X_9404_ _9758_/CLK _9404_/D _7011_/B VGND VGND VPWR VPWR _9404_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_153_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9335_ _9535_/CLK _9335_/D _9528_/SET_B VGND VGND VPWR VPWR _9335_/Q sky130_fd_sc_hd__dfstp_1
X_6547_ _6545_/Y _4613_/B _6546_/Y _4577_/B VGND VGND VPWR VPWR _6547_/X sky130_fd_sc_hd__o22a_2
XFILLER_192_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6478_ _9259_/Q VGND VGND VPWR VPWR _8757_/A sky130_fd_sc_hd__inv_6
X_9266_ _9354_/CLK _9266_/D _9685_/SET_B VGND VGND VPWR VPWR _9266_/Q sky130_fd_sc_hd__dfstp_1
Xoutput250 _8830_/X VGND VGND VPWR VPWR mgmt_gpio_out[37] sky130_fd_sc_hd__buf_2
XFILLER_160_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5429_ _9425_/Q _5422_/A _8930_/A1 _5422_/Y VGND VGND VPWR VPWR _9425_/D sky130_fd_sc_hd__a22o_1
X_8217_ _8341_/A _8341_/B _8009_/A _8215_/X _8216_/X VGND VGND VPWR VPWR _8217_/Y
+ sky130_fd_sc_hd__o2111ai_1
X_9197_ _9653_/CLK _9197_/D _9646_/SET_B VGND VGND VPWR VPWR _9197_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput261 _9729_/Q VGND VGND VPWR VPWR pll90_sel[0] sky130_fd_sc_hd__buf_2
X_8148_ _8148_/A _8577_/A VGND VGND VPWR VPWR _8150_/A sky130_fd_sc_hd__or2_1
Xoutput294 _9735_/Q VGND VGND VPWR VPWR pll_trim[3] sky130_fd_sc_hd__buf_2
Xoutput272 _9726_/Q VGND VGND VPWR VPWR pll_sel[0] sky130_fd_sc_hd__buf_2
Xoutput283 _9749_/Q VGND VGND VPWR VPWR pll_trim[17] sky130_fd_sc_hd__buf_2
XFILLER_181_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8079_ _8379_/D _8394_/B _8079_/C VGND VGND VPWR VPWR _8080_/A sky130_fd_sc_hd__or3_1
XFILLER_75_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_1_wb_clk_i clkbuf_1_1_1_wb_clk_i/A VGND VGND VPWR VPWR clkbuf_2_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_151_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4800_ _9515_/Q VGND VGND VPWR VPWR _4800_/Y sky130_fd_sc_hd__clkinv_2
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5780_ _9224_/Q _5778_/A _8845_/X _5778_/Y VGND VGND VPWR VPWR _9224_/D sky130_fd_sc_hd__a22o_1
XFILLER_34_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4731_ _4731_/A _5742_/B VGND VGND VPWR VPWR _4731_/X sky130_fd_sc_hd__or2_1
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7450_ _7474_/C _7466_/A _9255_/Q VGND VGND VPWR VPWR _7451_/A sky130_fd_sc_hd__or3_1
X_4662_ _4662_/A VGND VGND VPWR VPWR _4780_/B sky130_fd_sc_hd__buf_8
XFILLER_174_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6401_ _6396_/Y _5344_/B _6397_/Y _5298_/B _6400_/X VGND VGND VPWR VPWR _6408_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_174_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7381_ _6347_/Y _7097_/X _6340_/Y _7099_/X VGND VGND VPWR VPWR _7381_/X sky130_fd_sc_hd__o22a_1
X_4593_ _9739_/Q _4592_/A _8846_/X _4592_/Y VGND VGND VPWR VPWR _9739_/D sky130_fd_sc_hd__a22o_1
X_9120_ _9655_/CLK _9120_/D _7011_/B VGND VGND VPWR VPWR _9120_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_127_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6332_ _6330_/Y _5290_/B _6331_/Y _5916_/B VGND VGND VPWR VPWR _6332_/X sky130_fd_sc_hd__o22a_1
XFILLER_142_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6263_ _9551_/Q VGND VGND VPWR VPWR _6263_/Y sky130_fd_sc_hd__clkinv_4
X_9051_ _8837_/A1 _9051_/D _6045_/X VGND VGND VPWR VPWR _9051_/Q sky130_fd_sc_hd__dfrtp_4
X_8002_ _8394_/D _8077_/A VGND VGND VPWR VPWR _8009_/A sky130_fd_sc_hd__or2_1
XFILLER_88_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5214_ _5214_/A _5985_/B VGND VGND VPWR VPWR _5214_/Y sky130_fd_sc_hd__nor2_1
X_6194_ _9183_/Q VGND VGND VPWR VPWR _6194_/Y sky130_fd_sc_hd__clkinv_2
X_5145_ _6134_/A _5156_/B VGND VGND VPWR VPWR _5146_/A sky130_fd_sc_hd__or2_1
XFILLER_111_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5076_ _8962_/X _9660_/Q _5078_/S VGND VGND VPWR VPWR _5077_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8904_ _9624_/Q _8845_/X _8955_/S VGND VGND VPWR VPWR _8904_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8835_ _6582_/Y input92/X _8835_/S VGND VGND VPWR VPWR _8835_/X sky130_fd_sc_hd__mux2_1
X_8766_ _8766_/A VGND VGND VPWR VPWR _8766_/X sky130_fd_sc_hd__clkbuf_1
X_5978_ _9093_/Q _5970_/A _8839_/X _5970_/Y VGND VGND VPWR VPWR _9093_/D sky130_fd_sc_hd__a22o_1
X_8697_ _8697_/A VGND VGND VPWR VPWR _8697_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7717_ _9086_/Q _7716_/B _7718_/A VGND VGND VPWR VPWR _7717_/X sky130_fd_sc_hd__o21a_1
X_4929_ _4929_/A _4931_/B VGND VGND VPWR VPWR _5458_/B sky130_fd_sc_hd__or2_4
X_7648_ _6640_/Y _7415_/X _6772_/Y _7417_/X _7647_/X VGND VGND VPWR VPWR _7662_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_193_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7579_ _6224_/Y _7430_/X _6199_/Y _7432_/X _7578_/X VGND VGND VPWR VPWR _7579_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_153_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9318_ _9508_/CLK _9318_/D _9295_/SET_B VGND VGND VPWR VPWR _9318_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9249_ _9279_/CLK _9249_/D _9633_/SET_B VGND VGND VPWR VPWR _9249_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_106_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6950_ _6974_/B _6950_/B VGND VGND VPWR VPWR _6951_/A sky130_fd_sc_hd__or2_1
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5901_ _9136_/Q _5899_/A _8842_/X _5899_/Y VGND VGND VPWR VPWR _9136_/D sky130_fd_sc_hd__a22o_1
XFILLER_81_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6881_ input47/X _8955_/S input53/X _6322_/Y VGND VGND VPWR VPWR _6881_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_34_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8620_ _8706_/A _8705_/B _8703_/B _8620_/D VGND VGND VPWR VPWR _8620_/Y sky130_fd_sc_hd__nor4_1
X_5832_ _9189_/Q _5831_/A _5963_/B1 _5831_/Y VGND VGND VPWR VPWR _9189_/D sky130_fd_sc_hd__a22o_1
XFILLER_61_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5763_ _9235_/Q _5759_/A _8925_/A1 _5759_/Y VGND VGND VPWR VPWR _9235_/D sky130_fd_sc_hd__a22o_1
X_8551_ _8551_/A _8554_/B VGND VGND VPWR VPWR _8686_/C sky130_fd_sc_hd__nor2_1
XFILLER_14_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4714_ _7304_/A _5632_/B _4712_/Y _5789_/B VGND VGND VPWR VPWR _4714_/X sky130_fd_sc_hd__o22a_1
X_7502_ _6724_/Y _7400_/X _6664_/Y _7405_/X _7501_/X VGND VGND VPWR VPWR _7518_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_187_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8482_ _8562_/A _8650_/B VGND VGND VPWR VPWR _8605_/A sky130_fd_sc_hd__or2_1
XFILLER_108_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5694_ _5694_/A VGND VGND VPWR VPWR _7462_/A sky130_fd_sc_hd__buf_4
XFILLER_147_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4645_ _4645_/A VGND VGND VPWR VPWR _4645_/X sky130_fd_sc_hd__clkbuf_1
X_7433_ _7462_/A _7474_/C _7474_/D VGND VGND VPWR VPWR _7434_/A sky130_fd_sc_hd__or3_1
XFILLER_162_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7364_ _6498_/Y _7048_/D _6551_/Y _7040_/B _7363_/X VGND VGND VPWR VPWR _7365_/D
+ sky130_fd_sc_hd__o221a_1
X_4576_ _6158_/A _4876_/B VGND VGND VPWR VPWR _4577_/B sky130_fd_sc_hd__or2_4
XFILLER_190_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6315_ _9111_/Q VGND VGND VPWR VPWR _6315_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_1_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9103_ _9777_/CLK _9103_/D _9633_/SET_B VGND VGND VPWR VPWR _9103_/Q sky130_fd_sc_hd__dfstp_1
X_9034_ _9664_/CLK _9034_/D VGND VGND VPWR VPWR _9034_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7295_ _4902_/Y _7079_/B _4706_/Y _7059_/A VGND VGND VPWR VPWR _7295_/X sky130_fd_sc_hd__o22a_1
XFILLER_130_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6246_ _9447_/Q VGND VGND VPWR VPWR _6246_/Y sky130_fd_sc_hd__inv_2
X_6177_ _6175_/Y _5818_/B _6176_/Y _5572_/B VGND VGND VPWR VPWR _6187_/A sky130_fd_sc_hd__o22a_1
X_5128_ _9627_/Q _5123_/A _5967_/B1 _5123_/Y VGND VGND VPWR VPWR _9627_/D sky130_fd_sc_hd__a22o_1
XFILLER_29_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5059_ _7734_/A _5059_/B VGND VGND VPWR VPWR _5060_/A sky130_fd_sc_hd__and2_1
XFILLER_44_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8818_ _8818_/A VGND VGND VPWR VPWR _8818_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_158_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8749_ _8749_/A VGND VGND VPWR VPWR _8750_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_166_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_2 _7155_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6100_ _6100_/A VGND VGND VPWR VPWR _6100_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7080_ _7080_/A VGND VGND VPWR VPWR _8959_/S sky130_fd_sc_hd__buf_6
X_6031_ _9076_/Q _6029_/A _8845_/X _6029_/Y VGND VGND VPWR VPWR _9076_/D sky130_fd_sc_hd__a22o_1
XFILLER_140_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7982_ _7982_/A VGND VGND VPWR VPWR _8552_/A sky130_fd_sc_hd__clkbuf_4
X_6933_ _9191_/Q VGND VGND VPWR VPWR _6933_/Y sky130_fd_sc_hd__inv_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9721_ _9769_/CLK _9721_/D _9757_/SET_B VGND VGND VPWR VPWR _9721_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9652_ _9652_/CLK _9652_/D _9647_/SET_B VGND VGND VPWR VPWR _9652_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_81_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6864_ _6859_/Y _5496_/B _6860_/Y _5240_/B _6863_/X VGND VGND VPWR VPWR _6877_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_22_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8603_ _8603_/A _8603_/B _8603_/C _8603_/D VGND VGND VPWR VPWR _8604_/A sky130_fd_sc_hd__or4_1
X_5815_ _9200_/Q _5812_/A _8841_/X _5812_/Y VGND VGND VPWR VPWR _9200_/D sky130_fd_sc_hd__a22o_1
X_6795_ _9760_/Q VGND VGND VPWR VPWR _6795_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9583_ _9674_/CLK _9583_/D _9633_/SET_B VGND VGND VPWR VPWR _9583_/Q sky130_fd_sc_hd__dfrtp_1
X_5746_ _9243_/Q _5744_/A _8842_/X _5744_/Y VGND VGND VPWR VPWR _9243_/D sky130_fd_sc_hd__a22o_1
X_8534_ _8471_/Y _8523_/Y _8518_/X _8470_/B VGND VGND VPWR VPWR _8699_/A sky130_fd_sc_hd__a31o_1
XFILLER_182_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5677_ _9265_/Q _5673_/A _5966_/B1 _5673_/Y VGND VGND VPWR VPWR _9265_/D sky130_fd_sc_hd__a22o_1
X_8465_ _8305_/A _8270_/B _8097_/B _8552_/A VGND VGND VPWR VPWR _8615_/C sky130_fd_sc_hd__o22ai_1
XFILLER_135_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7416_ _7466_/A _7470_/B _9255_/Q VGND VGND VPWR VPWR _7417_/A sky130_fd_sc_hd__or3_1
X_4628_ _4628_/A VGND VGND VPWR VPWR _6052_/B sky130_fd_sc_hd__inv_2
XFILLER_163_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8396_ _8396_/A VGND VGND VPWR VPWR _8396_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7347_ _6731_/Y _7059_/D _6718_/Y _7116_/X _7346_/X VGND VGND VPWR VPWR _7352_/B
+ sky130_fd_sc_hd__o221a_1
X_4559_ _5966_/B1 _9757_/Q _4561_/S VGND VGND VPWR VPWR _4560_/A sky130_fd_sc_hd__mux2_1
XFILLER_131_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7278_ _6141_/Y _7112_/X _6128_/Y _7077_/B VGND VGND VPWR VPWR _7278_/X sky130_fd_sc_hd__o22a_1
X_9017_ _9664_/CLK _9017_/D VGND VGND VPWR VPWR _9017_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6229_ _6224_/Y _5905_/B _6225_/Y _5420_/B _6228_/X VGND VGND VPWR VPWR _6236_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_66_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput172 wb_dat_i[16] VGND VGND VPWR VPWR _7736_/B sky130_fd_sc_hd__clkbuf_1
Xinput150 wb_adr_i[26] VGND VGND VPWR VPWR input150/X sky130_fd_sc_hd__clkbuf_1
Xinput161 wb_adr_i[7] VGND VGND VPWR VPWR _8528_/A sky130_fd_sc_hd__buf_6
XFILLER_48_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput183 wb_dat_i[26] VGND VGND VPWR VPWR _7741_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput194 wb_dat_i[7] VGND VGND VPWR VPWR _8968_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_189_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5600_ _9308_/Q _5596_/A _8930_/A1 _5596_/Y VGND VGND VPWR VPWR _9308_/D sky130_fd_sc_hd__a22o_1
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6580_ _9691_/Q VGND VGND VPWR VPWR _8745_/A sky130_fd_sc_hd__clkinv_4
XFILLER_192_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5531_ _9356_/Q _5528_/A _8841_/X _5528_/Y VGND VGND VPWR VPWR _9356_/D sky130_fd_sc_hd__a22o_1
XFILLER_31_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8250_ _8250_/A VGND VGND VPWR VPWR _8597_/B sky130_fd_sc_hd__inv_2
X_7201_ _6371_/Y _7077_/C _6461_/Y _7077_/D _7200_/X VGND VGND VPWR VPWR _7201_/X
+ sky130_fd_sc_hd__o221a_1
X_5462_ _9404_/Q _5460_/A _8845_/X _5460_/Y VGND VGND VPWR VPWR _9404_/D sky130_fd_sc_hd__a22o_1
X_8181_ _8651_/A _8562_/A _8636_/A _8180_/Y VGND VGND VPWR VPWR _8182_/B sky130_fd_sc_hd__or4b_1
XFILLER_132_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5393_ _5545_/A _5393_/B VGND VGND VPWR VPWR _5394_/A sky130_fd_sc_hd__or2_1
X_7132_ _7132_/A _7132_/B _7132_/C VGND VGND VPWR VPWR _7133_/A sky130_fd_sc_hd__and3_4
XFILLER_113_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7063_ _7063_/A VGND VGND VPWR VPWR _7068_/B sky130_fd_sc_hd__buf_8
XFILLER_143_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6014_ _9083_/Q _5995_/A _8900_/X _5995_/Y VGND VGND VPWR VPWR _9083_/D sky130_fd_sc_hd__a22o_1
XFILLER_39_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9704_ _4446_/A1 _9704_/D _4975_/X VGND VGND VPWR VPWR _9704_/Q sky130_fd_sc_hd__dfrtp_1
X_7965_ _8583_/A _8091_/B VGND VGND VPWR VPWR _7971_/A sky130_fd_sc_hd__or2_2
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6916_ _9339_/Q VGND VGND VPWR VPWR _6916_/Y sky130_fd_sc_hd__inv_2
X_7896_ _7896_/A _8341_/B VGND VGND VPWR VPWR _7896_/X sky130_fd_sc_hd__or2_1
XFILLER_35_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6847_ _6847_/A VGND VGND VPWR VPWR _6847_/Y sky130_fd_sc_hd__inv_4
X_9635_ _9791_/CLK _9635_/D _9633_/SET_B VGND VGND VPWR VPWR _9635_/Q sky130_fd_sc_hd__dfrtp_1
X_9566_ _9617_/CLK _9566_/D _9295_/SET_B VGND VGND VPWR VPWR _9566_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_139_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6778_ _6778_/A VGND VGND VPWR VPWR _6778_/Y sky130_fd_sc_hd__inv_2
XFILLER_167_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8517_ _8517_/A VGND VGND VPWR VPWR _8517_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5729_ _6994_/A _5692_/Y _5724_/Y _5724_/B _5728_/X VGND VGND VPWR VPWR _5730_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_182_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9497_ _9501_/CLK _9497_/D _9647_/SET_B VGND VGND VPWR VPWR _9497_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_163_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8448_ _8612_/A _8448_/B _8448_/C _8447_/X VGND VGND VPWR VPWR _8449_/B sky130_fd_sc_hd__or4b_1
XFILLER_190_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8379_ _8202_/A _8379_/B _8379_/C _8379_/D VGND VGND VPWR VPWR _8585_/A sky130_fd_sc_hd__and4b_1
XFILLER_136_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7750_ _9066_/Q _7750_/B VGND VGND VPWR VPWR _7750_/X sky130_fd_sc_hd__and2_1
X_4962_ _4994_/A VGND VGND VPWR VPWR _4963_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_91_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7681_ _6399_/Y _7408_/X _6418_/Y _7410_/X VGND VGND VPWR VPWR _7681_/X sky130_fd_sc_hd__o22a_1
XFILLER_32_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4893_ _6111_/A _4917_/A VGND VGND VPWR VPWR _4893_/X sky130_fd_sc_hd__or2_4
X_6701_ _9330_/Q VGND VGND VPWR VPWR _6701_/Y sky130_fd_sc_hd__inv_2
X_9420_ _9684_/CLK _9420_/D _9685_/SET_B VGND VGND VPWR VPWR _9420_/Q sky130_fd_sc_hd__dfrtp_1
X_6632_ _9309_/Q VGND VGND VPWR VPWR _6632_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_149_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6563_ _9073_/Q VGND VGND VPWR VPWR _8783_/A sky130_fd_sc_hd__inv_8
XFILLER_177_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9351_ _9613_/CLK _9351_/D _9646_/SET_B VGND VGND VPWR VPWR _9351_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9282_ _9687_/CLK _9282_/D _9685_/SET_B VGND VGND VPWR VPWR _9282_/Q sky130_fd_sc_hd__dfrtp_1
X_5514_ _9367_/Q _5509_/A _8929_/A1 _5509_/Y VGND VGND VPWR VPWR _9367_/D sky130_fd_sc_hd__a22o_1
X_6494_ _8797_/A _6081_/B _7705_/A _5968_/B _6493_/X VGND VGND VPWR VPWR _6501_/C
+ sky130_fd_sc_hd__o221a_2
XFILLER_118_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8302_ _8498_/B VGND VGND VPWR VPWR _8302_/Y sky130_fd_sc_hd__inv_2
XFILLER_160_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5445_ _9415_/Q _5444_/A _5963_/B1 _5444_/Y VGND VGND VPWR VPWR _9415_/D sky130_fd_sc_hd__a22o_1
X_8233_ _8233_/A VGND VGND VPWR VPWR _8358_/B sky130_fd_sc_hd__inv_2
XFILLER_160_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8164_ _8164_/A _8168_/A VGND VGND VPWR VPWR _8708_/D sky130_fd_sc_hd__nor2_1
XFILLER_154_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5376_ _5376_/A VGND VGND VPWR VPWR _5376_/Y sky130_fd_sc_hd__inv_2
X_7115_ _7127_/C _7115_/B VGND VGND VPWR VPWR _7116_/A sky130_fd_sc_hd__or2_1
X_8095_ _8521_/A _8437_/B VGND VGND VPWR VPWR _8560_/A sky130_fd_sc_hd__nor2_1
XFILLER_113_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6039__1 _9709_/CLK VGND VGND VPWR VPWR _9058_/CLK sky130_fd_sc_hd__inv_4
X_7046_ _7125_/A _7127_/B _7073_/C VGND VGND VPWR VPWR _7047_/A sky130_fd_sc_hd__or3_1
XFILLER_86_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8997_ _9565_/Q _8771_/A VGND VGND VPWR VPWR mgmt_gpio_out[20] sky130_fd_sc_hd__ebufn_8
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7948_ _7948_/A VGND VGND VPWR VPWR _8378_/B sky130_fd_sc_hd__buf_12
XFILLER_103_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7879_ _7879_/A _7879_/B VGND VGND VPWR VPWR _7879_/Y sky130_fd_sc_hd__nor2_1
X_9618_ _9674_/CLK _9618_/D _9633_/SET_B VGND VGND VPWR VPWR _9618_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9549_ _9639_/CLK _9549_/D _9757_/SET_B VGND VGND VPWR VPWR _9549_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_7_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_8_csclk clkbuf_2_2_0_csclk/X VGND VGND VPWR VPWR _9358_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_73_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5230_ _5967_/B1 _9559_/Q _5230_/S VGND VGND VPWR VPWR _5231_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5161_ _9607_/Q _5158_/A _8844_/X _5158_/Y VGND VGND VPWR VPWR _9607_/D sky130_fd_sc_hd__a22o_1
XFILLER_142_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5092_ _9653_/Q _5091_/A _8846_/X _5091_/Y VGND VGND VPWR VPWR _9653_/D sky130_fd_sc_hd__a22o_1
XFILLER_110_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8920_ _9622_/Q _8925_/A1 _8955_/S VGND VGND VPWR VPWR _8920_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8851_ _8850_/X _9164_/Q _9054_/Q VGND VGND VPWR VPWR _8851_/X sky130_fd_sc_hd__mux2_1
X_8782_ _8782_/A VGND VGND VPWR VPWR _8782_/X sky130_fd_sc_hd__clkbuf_1
X_7802_ _7802_/A VGND VGND VPWR VPWR _8624_/B sky130_fd_sc_hd__buf_6
XFILLER_91_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5994_ _9051_/Q _5993_/X _6022_/B VGND VGND VPWR VPWR _5995_/A sky130_fd_sc_hd__o21ai_4
XFILLER_52_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7733_ _7733_/A _7734_/A _9066_/Q VGND VGND VPWR VPWR _7733_/X sky130_fd_sc_hd__and3_1
X_4945_ _7008_/A VGND VGND VPWR VPWR _5993_/B sky130_fd_sc_hd__clkinv_2
X_7664_ _6555_/Y _7400_/X _6497_/Y _7405_/X _7663_/X VGND VGND VPWR VPWR _7680_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_20_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4876_ _6111_/A _4876_/B VGND VGND VPWR VPWR _5110_/B sky130_fd_sc_hd__or2_4
XFILLER_192_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7595_ _6072_/Y _7427_/X _6141_/Y _5699_/X VGND VGND VPWR VPWR _7595_/X sky130_fd_sc_hd__o22a_1
X_6615_ _9487_/Q VGND VGND VPWR VPWR _6615_/Y sky130_fd_sc_hd__clkinv_4
X_9403_ _9758_/CLK _9403_/D _7011_/B VGND VGND VPWR VPWR _9403_/Q sky130_fd_sc_hd__dfrtp_1
X_9334_ _9532_/CLK _9334_/D _9647_/SET_B VGND VGND VPWR VPWR _9334_/Q sky130_fd_sc_hd__dfrtp_1
X_6546_ _9743_/Q VGND VGND VPWR VPWR _6546_/Y sky130_fd_sc_hd__inv_2
XFILLER_192_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9265_ _9789_/CLK _9265_/D _9685_/SET_B VGND VGND VPWR VPWR _9265_/Q sky130_fd_sc_hd__dfrtp_1
X_6477_ _9229_/Q VGND VGND VPWR VPWR _6477_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_160_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5428_ _9426_/Q _5422_/A _8841_/X _5422_/Y VGND VGND VPWR VPWR _9426_/D sky130_fd_sc_hd__a22o_1
X_8216_ _8510_/A _8341_/B VGND VGND VPWR VPWR _8216_/X sky130_fd_sc_hd__or2_2
X_9196_ _9653_/CLK _9196_/D _9646_/SET_B VGND VGND VPWR VPWR _9196_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput262 _9730_/Q VGND VGND VPWR VPWR pll90_sel[1] sky130_fd_sc_hd__buf_2
Xoutput251 _8837_/X VGND VGND VPWR VPWR pad_flash_clk sky130_fd_sc_hd__clkbuf_1
Xoutput240 _7704_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[4] sky130_fd_sc_hd__buf_2
X_5359_ _9474_/Q _5357_/A _8845_/X _5357_/Y VGND VGND VPWR VPWR _9474_/D sky130_fd_sc_hd__a22o_1
XFILLER_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8147_ _8213_/A _8551_/A VGND VGND VPWR VPWR _8577_/A sky130_fd_sc_hd__nor2_1
Xoutput295 _9736_/Q VGND VGND VPWR VPWR pll_trim[4] sky130_fd_sc_hd__buf_2
Xoutput273 _9727_/Q VGND VGND VPWR VPWR pll_sel[1] sky130_fd_sc_hd__buf_2
Xoutput284 _9750_/Q VGND VGND VPWR VPWR pll_trim[18] sky130_fd_sc_hd__buf_2
XFILLER_58_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8078_ _8078_/A _8672_/B VGND VGND VPWR VPWR _8082_/A sky130_fd_sc_hd__nor2_1
XFILLER_101_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7029_ _7073_/C _7123_/B VGND VGND VPWR VPWR _7030_/A sky130_fd_sc_hd__or2_1
XFILLER_114_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4730_ _4900_/B _4780_/B VGND VGND VPWR VPWR _5742_/B sky130_fd_sc_hd__or2_4
XFILLER_187_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4661_ _4665_/B _4665_/C _4661_/C VGND VGND VPWR VPWR _4662_/A sky130_fd_sc_hd__or3_1
XFILLER_174_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6400_ _6398_/Y _5534_/B _6399_/Y _5366_/B VGND VGND VPWR VPWR _6400_/X sky130_fd_sc_hd__o22a_1
XFILLER_80_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7380_ _6467_/Y _7048_/B _6416_/Y _7077_/A _7379_/X VGND VGND VPWR VPWR _7387_/A
+ sky130_fd_sc_hd__o221a_1
X_4592_ _4592_/A VGND VGND VPWR VPWR _4592_/Y sky130_fd_sc_hd__clkinv_2
X_6331_ _9124_/Q VGND VGND VPWR VPWR _6331_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_155_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6262_ _6262_/A VGND VGND VPWR VPWR _6262_/Y sky130_fd_sc_hd__clkinv_2
X_9050_ _8837_/A1 _9050_/D _6047_/X VGND VGND VPWR VPWR _9050_/Q sky130_fd_sc_hd__dfrtp_2
X_6193_ _6193_/A VGND VGND VPWR VPWR _6193_/Y sky130_fd_sc_hd__inv_2
XFILLER_142_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8001_ _8097_/B _8117_/A VGND VGND VPWR VPWR _8612_/A sky130_fd_sc_hd__nor2_1
X_5213_ _5213_/A VGND VGND VPWR VPWR _5213_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_142_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5144_ _9618_/Q _5136_/A _8916_/A1 _5136_/Y VGND VGND VPWR VPWR _9618_/D sky130_fd_sc_hd__a22o_1
XFILLER_96_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5075_ _5075_/A VGND VGND VPWR VPWR _9661_/D sky130_fd_sc_hd__clkbuf_1
X_8903_ _9619_/Q _8930_/A1 _8955_/S VGND VGND VPWR VPWR _8903_/X sky130_fd_sc_hd__mux2_1
X_8834_ _6485_/Y input90/X _8835_/S VGND VGND VPWR VPWR _8834_/X sky130_fd_sc_hd__mux2_2
XFILLER_71_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8765_ _8765_/A VGND VGND VPWR VPWR _8766_/A sky130_fd_sc_hd__clkbuf_1
X_5977_ _9094_/Q _5970_/A _8930_/A1 _5970_/Y VGND VGND VPWR VPWR _9094_/D sky130_fd_sc_hd__a22o_1
XFILLER_52_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8696_ _8696_/A _8696_/B _8696_/C _8727_/D VGND VGND VPWR VPWR _8697_/A sky130_fd_sc_hd__or4_1
X_4928_ _9398_/Q VGND VGND VPWR VPWR _4928_/Y sky130_fd_sc_hd__inv_2
X_7716_ _9086_/Q _7716_/B VGND VGND VPWR VPWR _7718_/A sky130_fd_sc_hd__nand2_1
XFILLER_193_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7647_ _6732_/Y _7419_/X _6762_/Y _7421_/X VGND VGND VPWR VPWR _7647_/X sky130_fd_sc_hd__o22a_1
XFILLER_165_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4859_ _4931_/A _4911_/A VGND VGND VPWR VPWR _5374_/B sky130_fd_sc_hd__or2_4
XFILLER_193_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7578_ _6171_/Y _7434_/X _6169_/Y _7436_/X VGND VGND VPWR VPWR _7578_/X sky130_fd_sc_hd__o22a_1
X_6529_ _9686_/Q VGND VGND VPWR VPWR _6529_/Y sky130_fd_sc_hd__clkinv_4
X_9317_ _9501_/CLK _9317_/D _9647_/SET_B VGND VGND VPWR VPWR _9317_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9248_ _9279_/CLK _9248_/D _9779_/SET_B VGND VGND VPWR VPWR _9248_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_192_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9179_ _9652_/CLK _9179_/D _9646_/SET_B VGND VGND VPWR VPWR _9179_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_121_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_11_csclk clkbuf_2_2_0_csclk/X VGND VGND VPWR VPWR _9527_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_169_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_26_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR _9613_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_140_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5900_ _9137_/Q _5899_/A _8843_/X _5899_/Y VGND VGND VPWR VPWR _9137_/D sky130_fd_sc_hd__a22o_1
XFILLER_75_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6880_ _9295_/Q VGND VGND VPWR VPWR _7150_/A sky130_fd_sc_hd__inv_2
XFILLER_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5831_ _5831_/A VGND VGND VPWR VPWR _5831_/Y sky130_fd_sc_hd__inv_2
X_5762_ _9236_/Q _5759_/A _8844_/X _5759_/Y VGND VGND VPWR VPWR _9236_/D sky130_fd_sc_hd__a22o_1
X_8550_ _8550_/A _8554_/B VGND VGND VPWR VPWR _8627_/D sky130_fd_sc_hd__nor2_1
X_7501_ _6736_/Y _7408_/X _6673_/Y _7410_/X VGND VGND VPWR VPWR _7501_/X sky130_fd_sc_hd__o22a_1
X_4713_ _4919_/A _4780_/B VGND VGND VPWR VPWR _5789_/B sky130_fd_sc_hd__or2_4
XFILLER_147_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8481_ _8481_/A _8706_/A VGND VGND VPWR VPWR _8483_/A sky130_fd_sc_hd__or2_1
X_5693_ _9252_/Q _9251_/Q VGND VGND VPWR VPWR _5694_/A sky130_fd_sc_hd__or2_1
X_4644_ _4994_/A VGND VGND VPWR VPWR _4645_/A sky130_fd_sc_hd__clkbuf_1
X_7432_ _7432_/A VGND VGND VPWR VPWR _7432_/X sky130_fd_sc_hd__buf_6
X_4575_ _4669_/A _4729_/D _4729_/A _8944_/X VGND VGND VPWR VPWR _4876_/B sky130_fd_sc_hd__or4_4
X_7363_ _6581_/Y _7068_/A _6597_/Y _7105_/X VGND VGND VPWR VPWR _7363_/X sky130_fd_sc_hd__o22a_1
X_6314_ _9651_/Q VGND VGND VPWR VPWR _6314_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7294_ _4924_/Y _7095_/X _4722_/Y _7068_/D _7293_/X VGND VGND VPWR VPWR _7299_/B
+ sky130_fd_sc_hd__o221a_1
X_9102_ _9775_/CLK _9102_/D _7011_/B VGND VGND VPWR VPWR _9102_/Q sky130_fd_sc_hd__dfrtp_1
X_9033_ _9664_/CLK _9033_/D VGND VGND VPWR VPWR _9033_/Q sky130_fd_sc_hd__dfxtp_1
X_6245_ _6245_/A VGND VGND VPWR VPWR _6245_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_115_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6176_ _9326_/Q VGND VGND VPWR VPWR _6176_/Y sky130_fd_sc_hd__clkinv_2
X_5127_ _9628_/Q _5123_/A _5966_/B1 _5123_/Y VGND VGND VPWR VPWR _9628_/D sky130_fd_sc_hd__a22o_1
X_5058_ _7734_/A _5058_/B VGND VGND VPWR VPWR _5058_/X sky130_fd_sc_hd__and2_1
XFILLER_84_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8817_ _8817_/A VGND VGND VPWR VPWR _8817_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_111_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8748_ _8748_/A VGND VGND VPWR VPWR _8748_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8679_ _8721_/A _8720_/C _8721_/C _8723_/C VGND VGND VPWR VPWR _8680_/C sky130_fd_sc_hd__or4_4
XFILLER_166_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_mgmt_gpio_in[4] clkbuf_2_3_0_mgmt_gpio_in[4]/A VGND VGND VPWR VPWR _9089_/CLK
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_90_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_3 _7155_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6030_ _9077_/Q _6029_/A _8846_/X _6029_/Y VGND VGND VPWR VPWR _9077_/D sky130_fd_sc_hd__a22o_1
XFILLER_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7981_ _7995_/B _7992_/B VGND VGND VPWR VPWR _7982_/A sky130_fd_sc_hd__or2_1
XFILLER_81_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9720_ _9770_/CLK _9720_/D _7011_/B VGND VGND VPWR VPWR _9720_/Q sky130_fd_sc_hd__dfstp_1
X_6932_ _9213_/Q VGND VGND VPWR VPWR _6932_/Y sky130_fd_sc_hd__inv_2
X_9651_ _9653_/CLK _9651_/D _9646_/SET_B VGND VGND VPWR VPWR _9651_/Q sky130_fd_sc_hd__dfrtp_1
X_6863_ _6861_/Y _4577_/B _8808_/A _5227_/B VGND VGND VPWR VPWR _6863_/X sky130_fd_sc_hd__o22a_2
XFILLER_179_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8602_ _8202_/A _8341_/A _8660_/C _7881_/A _8334_/X VGND VGND VPWR VPWR _8603_/D
+ sky130_fd_sc_hd__o221ai_1
X_5814_ _9201_/Q _5812_/A _5964_/B1 _5812_/Y VGND VGND VPWR VPWR _9201_/D sky130_fd_sc_hd__a22o_1
X_6794_ _6794_/A VGND VGND VPWR VPWR _6794_/Y sky130_fd_sc_hd__inv_2
X_9582_ _9674_/CLK _9582_/D _9633_/SET_B VGND VGND VPWR VPWR _9582_/Q sky130_fd_sc_hd__dfrtp_1
X_5745_ _9244_/Q _5744_/A _8843_/X _5744_/Y VGND VGND VPWR VPWR _9244_/D sky130_fd_sc_hd__a22o_1
X_8533_ _8516_/Y _8528_/Y _8518_/X _8464_/D VGND VGND VPWR VPWR _8615_/D sky130_fd_sc_hd__a31o_1
XFILLER_41_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5676_ _9266_/Q _5673_/A _8841_/X _5673_/Y VGND VGND VPWR VPWR _9266_/D sky130_fd_sc_hd__a22o_1
X_8464_ _8464_/A _8464_/B _8668_/A _8464_/D VGND VGND VPWR VPWR _8466_/A sky130_fd_sc_hd__or4_1
XFILLER_108_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4627_ _4627_/A VGND VGND VPWR VPWR _9719_/D sky130_fd_sc_hd__clkbuf_1
X_7415_ _7415_/A VGND VGND VPWR VPWR _7415_/X sky130_fd_sc_hd__buf_6
XFILLER_190_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8395_ _8496_/A _8395_/B VGND VGND VPWR VPWR _8395_/X sky130_fd_sc_hd__or2_1
XFILLER_190_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4558_ _5259_/A _4558_/B VGND VGND VPWR VPWR _4561_/S sky130_fd_sc_hd__or2_1
X_7346_ _6779_/Y _7118_/X _6668_/Y _7048_/C VGND VGND VPWR VPWR _7346_/X sky130_fd_sc_hd__o22a_1
XFILLER_143_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7277_ _7277_/A _7277_/B _7277_/C _7277_/D VGND VGND VPWR VPWR _7287_/B sky130_fd_sc_hd__and4_1
XFILLER_103_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4489_ _8934_/X _8932_/X _8946_/X _8944_/X VGND VGND VPWR VPWR _4805_/A sky130_fd_sc_hd__or4_4
X_9016_ _9039_/CLK _9016_/D VGND VGND VPWR VPWR _9016_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6228_ _6226_/Y _4524_/B _6227_/Y _4832_/X VGND VGND VPWR VPWR _6228_/X sky130_fd_sc_hd__o22a_2
X_6159_ _9456_/Q VGND VGND VPWR VPWR _6159_/Y sky130_fd_sc_hd__inv_2
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater370 _9779_/SET_B VGND VGND VPWR VPWR _9646_/SET_B sky130_fd_sc_hd__buf_12
XFILLER_82_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput151 wb_adr_i[27] VGND VGND VPWR VPWR _5930_/A sky130_fd_sc_hd__clkbuf_1
Xinput140 wb_adr_i[17] VGND VGND VPWR VPWR _7768_/A sky130_fd_sc_hd__clkbuf_1
Xinput162 wb_adr_i[8] VGND VGND VPWR VPWR _7774_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput184 wb_dat_i[27] VGND VGND VPWR VPWR _7743_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput173 wb_dat_i[17] VGND VGND VPWR VPWR _7738_/B sky130_fd_sc_hd__clkbuf_1
Xinput195 wb_dat_i[8] VGND VGND VPWR VPWR _7737_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5530_ _9357_/Q _5528_/A _8842_/X _5528_/Y VGND VGND VPWR VPWR _9357_/D sky130_fd_sc_hd__a22o_1
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5461_ _9405_/Q _5460_/A _8846_/X _5460_/Y VGND VGND VPWR VPWR _9405_/D sky130_fd_sc_hd__a22o_1
XFILLER_172_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7200_ _6415_/Y _7086_/X _6357_/Y _7088_/X VGND VGND VPWR VPWR _7200_/X sky130_fd_sc_hd__o22a_1
X_5392_ _9450_/Q _5384_/A _8916_/A1 _5384_/Y VGND VGND VPWR VPWR _9450_/D sky130_fd_sc_hd__a22o_1
XFILLER_172_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8180_ _8544_/A _8092_/Y _8179_/X VGND VGND VPWR VPWR _8180_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7131_ _7131_/A _7131_/B _7131_/C _7131_/D VGND VGND VPWR VPWR _7132_/C sky130_fd_sc_hd__and4_1
XFILLER_98_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7062_ _7075_/A _7087_/B VGND VGND VPWR VPWR _7063_/A sky130_fd_sc_hd__or2_1
XFILLER_98_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6013_ _6013_/A VGND VGND VPWR VPWR _6013_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_67_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7964_ _8189_/A _8099_/B _7966_/B VGND VGND VPWR VPWR _8091_/B sky130_fd_sc_hd__a21bo_2
XFILLER_82_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9703_ _4446_/A1 _9703_/D _4978_/X VGND VGND VPWR VPWR _9703_/Q sky130_fd_sc_hd__dfrtp_1
X_6915_ _9365_/Q VGND VGND VPWR VPWR _6915_/Y sky130_fd_sc_hd__clkinv_2
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7895_ _7895_/A VGND VGND VPWR VPWR _8341_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_35_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9634_ _9655_/CLK _9634_/D _9633_/SET_B VGND VGND VPWR VPWR _9634_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6846_ _6844_/Y _4491_/B _6845_/Y _5259_/B VGND VGND VPWR VPWR _6846_/X sky130_fd_sc_hd__o22a_1
X_9565_ _9617_/CLK _9565_/D _9295_/SET_B VGND VGND VPWR VPWR _9565_/Q sky130_fd_sc_hd__dfrtp_4
X_6777_ _6772_/Y _5941_/B _6773_/Y _5089_/B _6776_/X VGND VGND VPWR VPWR _6783_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_50_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8516_ _8525_/C _8516_/B VGND VGND VPWR VPWR _8516_/Y sky130_fd_sc_hd__nor2_4
X_5728_ _5728_/A VGND VGND VPWR VPWR _5728_/X sky130_fd_sc_hd__buf_8
X_9496_ _9532_/CLK _9496_/D _9647_/SET_B VGND VGND VPWR VPWR _9496_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8447_ _8496_/A _8447_/B VGND VGND VPWR VPWR _8447_/X sky130_fd_sc_hd__or2_1
XFILLER_108_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5659_ _5647_/A _5658_/A _9277_/Q _5658_/Y _5651_/X VGND VGND VPWR VPWR _9277_/D
+ sky130_fd_sc_hd__o221a_1
X_8378_ _8565_/A _8378_/B VGND VGND VPWR VPWR _8720_/C sky130_fd_sc_hd__nor2_1
XFILLER_163_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7329_ _6872_/Y _7124_/X _6885_/Y _7068_/B _7328_/X VGND VGND VPWR VPWR _7330_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_131_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4961_ _9092_/Q _9048_/Q _4949_/A _4958_/Y _4960_/X VGND VGND VPWR VPWR _9708_/D
+ sky130_fd_sc_hd__a41o_1
X_7680_ _7680_/A _7680_/B _7680_/C _7680_/D VGND VGND VPWR VPWR _7680_/Y sky130_fd_sc_hd__nand4_4
X_6700_ _9387_/Q VGND VGND VPWR VPWR _6700_/Y sky130_fd_sc_hd__inv_2
X_4892_ _4892_/A VGND VGND VPWR VPWR _4892_/Y sky130_fd_sc_hd__inv_2
X_6631_ _9296_/Q VGND VGND VPWR VPWR _7172_/A sky130_fd_sc_hd__inv_2
XFILLER_32_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9350_ _9352_/CLK _9350_/D _9646_/SET_B VGND VGND VPWR VPWR _9350_/Q sky130_fd_sc_hd__dfrtp_1
X_6562_ _9471_/Q VGND VGND VPWR VPWR _8791_/A sky130_fd_sc_hd__inv_12
X_8301_ _8301_/A VGND VGND VPWR VPWR _8498_/B sky130_fd_sc_hd__buf_6
X_9281_ _9687_/CLK _9281_/D _9528_/SET_B VGND VGND VPWR VPWR _9281_/Q sky130_fd_sc_hd__dfrtp_1
X_5513_ _9368_/Q _5509_/A _8925_/A1 _5509_/Y VGND VGND VPWR VPWR _9368_/D sky130_fd_sc_hd__a22o_1
X_6493_ _6491_/Y _5545_/B _8751_/A _5797_/B VGND VGND VPWR VPWR _6493_/X sky130_fd_sc_hd__o22a_1
XFILLER_133_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5444_ _5444_/A VGND VGND VPWR VPWR _5444_/Y sky130_fd_sc_hd__inv_2
X_8232_ _8341_/A _8232_/B VGND VGND VPWR VPWR _8233_/A sky130_fd_sc_hd__or2_1
XFILLER_172_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8163_ _8708_/B _8163_/B VGND VGND VPWR VPWR _8165_/A sky130_fd_sc_hd__or2_1
XFILLER_160_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5375_ _5375_/A VGND VGND VPWR VPWR _5376_/A sky130_fd_sc_hd__clkbuf_2
X_7114_ _4716_/Y _7040_/D _4804_/Y _7110_/X _7113_/X VGND VGND VPWR VPWR _7131_/A
+ sky130_fd_sc_hd__o221a_1
X_8094_ _8094_/A VGND VGND VPWR VPWR _8720_/A sky130_fd_sc_hd__inv_2
XFILLER_101_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7045_ _7045_/A VGND VGND VPWR VPWR _7048_/C sky130_fd_sc_hd__buf_8
XFILLER_170_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8996_ _9564_/Q _8769_/A VGND VGND VPWR VPWR mgmt_gpio_out[19] sky130_fd_sc_hd__ebufn_8
XFILLER_55_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7947_ _8379_/D _8379_/B _8079_/C VGND VGND VPWR VPWR _7948_/A sky130_fd_sc_hd__or3_1
XFILLER_82_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7878_ _7878_/A _8341_/A VGND VGND VPWR VPWR _7879_/B sky130_fd_sc_hd__or2_2
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9617_ _9617_/CLK _9617_/D _9295_/SET_B VGND VGND VPWR VPWR _9617_/Q sky130_fd_sc_hd__dfrtp_1
X_6829_ _6829_/A _6829_/B _6829_/C _6829_/D VGND VGND VPWR VPWR _6830_/D sky130_fd_sc_hd__and4_1
XFILLER_156_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9548_ _9639_/CLK _9548_/D _9633_/SET_B VGND VGND VPWR VPWR _9548_/Q sky130_fd_sc_hd__dfrtp_1
X_9479_ _9684_/CLK _9479_/D _9685_/SET_B VGND VGND VPWR VPWR _9479_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_183_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5160_ _9608_/Q _5158_/A _8845_/X _5158_/Y VGND VGND VPWR VPWR _9608_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5091_ _5091_/A VGND VGND VPWR VPWR _5091_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_68_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8850_ _7500_/Y _9633_/Q _8978_/S VGND VGND VPWR VPWR _8850_/X sky130_fd_sc_hd__mux2_1
X_8781_ _8781_/A VGND VGND VPWR VPWR _8782_/A sky130_fd_sc_hd__clkbuf_1
X_7801_ _8394_/B _8093_/A VGND VGND VPWR VPWR _7802_/A sky130_fd_sc_hd__or2_1
XFILLER_64_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5993_ _9050_/Q _5993_/B _7008_/B VGND VGND VPWR VPWR _5993_/X sky130_fd_sc_hd__and3_1
X_7732_ _7732_/A VGND VGND VPWR VPWR _8960_/S sky130_fd_sc_hd__clkbuf_1
X_4944_ _4944_/A VGND VGND VPWR VPWR _7008_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_149_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7663_ _6589_/Y _7408_/X _6529_/Y _7410_/X VGND VGND VPWR VPWR _7663_/X sky130_fd_sc_hd__o22a_1
X_4875_ _9632_/Q VGND VGND VPWR VPWR _4875_/Y sky130_fd_sc_hd__inv_2
X_9402_ _9758_/CLK _9402_/D _7011_/B VGND VGND VPWR VPWR _9402_/Q sky130_fd_sc_hd__dfrtp_1
X_7594_ _6126_/Y _7415_/X _6120_/Y _7417_/X _7593_/X VGND VGND VPWR VPWR _7608_/B
+ sky130_fd_sc_hd__o221a_1
X_6614_ _6609_/Y _5251_/B _8765_/A _5534_/B _6613_/X VGND VGND VPWR VPWR _6627_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_192_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9333_ _9535_/CLK _9333_/D _9528_/SET_B VGND VGND VPWR VPWR _9333_/Q sky130_fd_sc_hd__dfrtp_1
X_6545_ _9724_/Q VGND VGND VPWR VPWR _6545_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9264_ _9354_/CLK _9264_/D _9685_/SET_B VGND VGND VPWR VPWR _9264_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6476_ _6149_/A _6475_/Y _9040_/Q _6149_/Y VGND VGND VPWR VPWR _9040_/D sky130_fd_sc_hd__o22a_2
XFILLER_145_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8215_ _8660_/A _8498_/A VGND VGND VPWR VPWR _8215_/X sky130_fd_sc_hd__or2_2
XFILLER_133_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5427_ _9427_/Q _5422_/A _8929_/A1 _5422_/Y VGND VGND VPWR VPWR _9427_/D sky130_fd_sc_hd__a22o_1
X_9195_ _9653_/CLK _9195_/D _9646_/SET_B VGND VGND VPWR VPWR _9195_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput241 _8746_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[5] sky130_fd_sc_hd__buf_2
Xoutput252 _7011_/Y VGND VGND VPWR VPWR pad_flash_clk_oeb sky130_fd_sc_hd__buf_2
Xoutput230 _8744_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[2] sky130_fd_sc_hd__buf_2
X_5358_ _9475_/Q _5357_/A _8846_/X _5357_/Y VGND VGND VPWR VPWR _9475_/D sky130_fd_sc_hd__a22o_1
X_8146_ _7987_/Y _8544_/B _8145_/X VGND VGND VPWR VPWR _8148_/A sky130_fd_sc_hd__a21o_1
Xoutput263 _9731_/Q VGND VGND VPWR VPWR pll90_sel[2] sky130_fd_sc_hd__buf_2
Xoutput274 _9728_/Q VGND VGND VPWR VPWR pll_sel[2] sky130_fd_sc_hd__buf_2
Xoutput285 _9751_/Q VGND VGND VPWR VPWR pll_trim[19] sky130_fd_sc_hd__buf_2
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8077_ _8077_/A _8437_/B VGND VGND VPWR VPWR _8672_/B sky130_fd_sc_hd__nor2_1
XFILLER_101_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput296 _9737_/Q VGND VGND VPWR VPWR pll_trim[5] sky130_fd_sc_hd__buf_2
X_5289_ _6052_/A VGND VGND VPWR VPWR _5671_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_75_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7028_ _7104_/A _7111_/C VGND VGND VPWR VPWR _7123_/B sky130_fd_sc_hd__or2_1
XFILLER_74_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8979_ _9580_/Q _8743_/A VGND VGND VPWR VPWR mgmt_gpio_out[2] sky130_fd_sc_hd__ebufn_8
XFILLER_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xnet299_2 _4446_/A1 VGND VGND VPWR VPWR _7022_/A sky130_fd_sc_hd__inv_4
XFILLER_61_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4660_ _9333_/Q VGND VGND VPWR VPWR _4660_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6330_ _9519_/Q VGND VGND VPWR VPWR _6330_/Y sky130_fd_sc_hd__clkinv_2
X_4591_ _4591_/A VGND VGND VPWR VPWR _4592_/A sky130_fd_sc_hd__buf_2
XFILLER_127_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6261_ _6256_/Y _5355_/B _6257_/Y _4870_/X _6260_/X VGND VGND VPWR VPWR _6280_/A
+ sky130_fd_sc_hd__o221a_1
X_8000_ _8000_/A VGND VGND VPWR VPWR _8117_/A sky130_fd_sc_hd__buf_6
XFILLER_130_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6192_ _6188_/Y _6027_/B _6189_/Y _4491_/B _6191_/X VGND VGND VPWR VPWR _6211_/A
+ sky130_fd_sc_hd__o221a_1
X_5212_ _6040_/A VGND VGND VPWR VPWR _5213_/A sky130_fd_sc_hd__clkbuf_1
X_5143_ _9619_/Q _5136_/A _8930_/A1 _5136_/Y VGND VGND VPWR VPWR _9619_/D sky130_fd_sc_hd__a22o_1
XFILLER_57_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5074_ _8963_/X _9661_/Q _5078_/S VGND VGND VPWR VPWR _5075_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8902_ _7708_/Y _4949_/A _9051_/Q VGND VGND VPWR VPWR _8902_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8833_ _6491_/Y input82/X _8833_/S VGND VGND VPWR VPWR _8833_/X sky130_fd_sc_hd__mux2_4
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8764_ _8764_/A VGND VGND VPWR VPWR _8764_/X sky130_fd_sc_hd__clkbuf_1
X_5976_ _9095_/Q _5970_/A _8841_/X _5970_/Y VGND VGND VPWR VPWR _9095_/D sky130_fd_sc_hd__a22o_1
XFILLER_178_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8695_ _8695_/A _8695_/B _8695_/C _8695_/D VGND VGND VPWR VPWR _8727_/D sky130_fd_sc_hd__or4_1
X_4927_ _4927_/A _4931_/B VGND VGND VPWR VPWR _5306_/B sky130_fd_sc_hd__or2_4
X_7715_ _7716_/B _7715_/B VGND VGND VPWR VPWR _7715_/Y sky130_fd_sc_hd__nor2_1
XFILLER_52_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4858_ _9458_/Q VGND VGND VPWR VPWR _4858_/Y sky130_fd_sc_hd__inv_2
X_7646_ _6718_/Y _7400_/X _6645_/Y _7405_/X _7645_/X VGND VGND VPWR VPWR _7662_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_100_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9316_ _9534_/CLK _9316_/D _9647_/SET_B VGND VGND VPWR VPWR _9316_/Q sky130_fd_sc_hd__dfrtp_1
X_4789_ _4779_/Y _5757_/B _4781_/Y _6322_/A _4788_/X VGND VGND VPWR VPWR _4790_/D
+ sky130_fd_sc_hd__o221a_1
X_7577_ _6200_/Y _7427_/X _6176_/Y _5699_/X VGND VGND VPWR VPWR _7577_/X sky130_fd_sc_hd__o22a_1
X_6528_ _9136_/Q VGND VGND VPWR VPWR _6528_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_7_csclk clkbuf_2_2_0_csclk/X VGND VGND VPWR VPWR _9354_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_109_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6459_ _6457_/Y _5837_/B _6458_/Y _5960_/B VGND VGND VPWR VPWR _6459_/X sky130_fd_sc_hd__o22a_1
X_9247_ _9279_/CLK _9247_/D _9779_/SET_B VGND VGND VPWR VPWR _9247_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_9178_ _9613_/CLK _9178_/D _9646_/SET_B VGND VGND VPWR VPWR _9178_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_121_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8129_ _8130_/B _8378_/B VGND VGND VPWR VPWR _8357_/A sky130_fd_sc_hd__nor2_1
XFILLER_87_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5830_ _5830_/A VGND VGND VPWR VPWR _5831_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_34_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5761_ _9237_/Q _5759_/A _8845_/X _5759_/Y VGND VGND VPWR VPWR _9237_/D sky130_fd_sc_hd__a22o_1
X_8480_ _8515_/B _8437_/B _8521_/B _8437_/B VGND VGND VPWR VPWR _8706_/A sky130_fd_sc_hd__o22ai_4
X_7500_ _7500_/A _7500_/B _7500_/C _7500_/D VGND VGND VPWR VPWR _7500_/Y sky130_fd_sc_hd__nand4_4
XFILLER_30_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4712_ _9212_/Q VGND VGND VPWR VPWR _4712_/Y sky130_fd_sc_hd__inv_2
XFILLER_187_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5692_ _5692_/A VGND VGND VPWR VPWR _5692_/Y sky130_fd_sc_hd__inv_2
X_7431_ _7474_/C _7472_/A _7474_/D VGND VGND VPWR VPWR _7432_/A sky130_fd_sc_hd__or3_1
XFILLER_175_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4643_ hold1/A _4636_/A _8947_/X _4636_/Y VGND VGND VPWR VPWR _9716_/D sky130_fd_sc_hd__a22o_1
XFILLER_128_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7362_ _6522_/Y _7059_/B _6557_/Y _7068_/C _7361_/X VGND VGND VPWR VPWR _7365_/C
+ sky130_fd_sc_hd__o221a_1
X_4574_ _9748_/Q _4566_/A _5967_/B1 _4566_/Y VGND VGND VPWR VPWR _9748_/D sky130_fd_sc_hd__a22o_1
XFILLER_143_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6313_ _6308_/Y _5757_/B _6309_/Y _5679_/B _6312_/X VGND VGND VPWR VPWR _6325_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_115_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7293_ _4930_/Y _7097_/X _4883_/Y _7099_/X VGND VGND VPWR VPWR _7293_/X sky130_fd_sc_hd__o22a_1
X_9101_ _9777_/CLK _9101_/D _7011_/B VGND VGND VPWR VPWR _9101_/Q sky130_fd_sc_hd__dfrtp_1
X_9032_ _9039_/CLK _9032_/D VGND VGND VPWR VPWR _9032_/Q sky130_fd_sc_hd__dfxtp_1
X_6244_ _9499_/Q VGND VGND VPWR VPWR _6244_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_89_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6175_ _9196_/Q VGND VGND VPWR VPWR _6175_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_97_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5126_ _9629_/Q _5123_/A _5965_/B1 _5123_/Y VGND VGND VPWR VPWR _9629_/D sky130_fd_sc_hd__a22o_1
XFILLER_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5057_ _7734_/A _7734_/B _8813_/A VGND VGND VPWR VPWR _5062_/B sky130_fd_sc_hd__a21oi_1
XFILLER_111_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8816_ _8816_/A VGND VGND VPWR VPWR _8816_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5959_ _9106_/Q _5951_/A _8916_/A1 _5951_/Y VGND VGND VPWR VPWR _9106_/D sky130_fd_sc_hd__a22o_1
X_8747_ _8747_/A VGND VGND VPWR VPWR _8748_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_52_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8678_ _8678_/A _8678_/B _8678_/C VGND VGND VPWR VPWR _8723_/C sky130_fd_sc_hd__or3_2
XFILLER_166_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7629_ _6940_/Y _7419_/X _6868_/Y _7421_/X VGND VGND VPWR VPWR _7629_/X sky130_fd_sc_hd__o22a_1
XFILLER_193_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_4 _7177_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7980_ _8528_/A _7994_/A VGND VGND VPWR VPWR _7992_/B sky130_fd_sc_hd__or2_4
XFILLER_94_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6931_ _6926_/Y _5660_/B _6927_/Y _5742_/B _6930_/X VGND VGND VPWR VPWR _6944_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9650_ _9653_/CLK _9650_/D _9646_/SET_B VGND VGND VPWR VPWR _9650_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6862_ _9560_/Q VGND VGND VPWR VPWR _8808_/A sky130_fd_sc_hd__clkinv_2
XFILLER_50_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_8601_ _8601_/A _8696_/A _8662_/C _8601_/D VGND VGND VPWR VPWR _8603_/B sky130_fd_sc_hd__or4_1
X_5813_ _9202_/Q _5812_/A _8843_/X _5812_/Y VGND VGND VPWR VPWR _9202_/D sky130_fd_sc_hd__a22o_1
XFILLER_62_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9581_ _9620_/CLK _9581_/D _9633_/SET_B VGND VGND VPWR VPWR _9581_/Q sky130_fd_sc_hd__dfrtp_1
X_6793_ _9347_/Q VGND VGND VPWR VPWR _6793_/Y sky130_fd_sc_hd__clkinv_4
X_8532_ _8528_/Y _8525_/Y _8518_/X _8464_/B VGND VGND VPWR VPWR _8668_/C sky130_fd_sc_hd__a31o_1
X_5744_ _5744_/A VGND VGND VPWR VPWR _5744_/Y sky130_fd_sc_hd__inv_2
X_5675_ _9267_/Q _5673_/A _8842_/X _5673_/Y VGND VGND VPWR VPWR _9267_/D sky130_fd_sc_hd__a22o_1
X_8463_ _8463_/A _8685_/A VGND VGND VPWR VPWR _8464_/D sky130_fd_sc_hd__or2_1
X_8394_ _8394_/A _8394_/B _8394_/C _8394_/D VGND VGND VPWR VPWR _8395_/B sky130_fd_sc_hd__or4_2
XFILLER_135_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4626_ _5967_/B1 _9719_/Q _4626_/S VGND VGND VPWR VPWR _4627_/A sky130_fd_sc_hd__mux2_1
X_7414_ _7474_/C _7472_/A _9255_/Q VGND VGND VPWR VPWR _7415_/A sky130_fd_sc_hd__or3_1
XFILLER_163_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7345_ _6674_/Y _7040_/D _6662_/Y _7110_/X _7344_/X VGND VGND VPWR VPWR _7352_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_190_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4557_ _6111_/A _4805_/A VGND VGND VPWR VPWR _4558_/B sky130_fd_sc_hd__or2_2
XFILLER_171_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_7276_ _6121_/Y _7048_/D _6062_/Y _7040_/B _7275_/X VGND VGND VPWR VPWR _7277_/D
+ sky130_fd_sc_hd__o221a_1
X_4488_ _4488_/A VGND VGND VPWR VPWR _4911_/A sky130_fd_sc_hd__buf_6
X_9015_ _9039_/CLK _9015_/D VGND VGND VPWR VPWR _9015_/Q sky130_fd_sc_hd__dfxtp_1
X_6227_ _6227_/A VGND VGND VPWR VPWR _6227_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6158_ _6158_/A _6158_/B VGND VGND VPWR VPWR _6158_/X sky130_fd_sc_hd__or2_4
Xclkbuf_leaf_10_csclk clkbuf_2_2_0_csclk/X VGND VGND VPWR VPWR _9684_/CLK sky130_fd_sc_hd__clkbuf_16
X_5109_ _9640_/Q _5108_/X _7731_/A _5062_/D VGND VGND VPWR VPWR _9640_/D sky130_fd_sc_hd__o211a_2
XFILLER_111_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater360 _8843_/X VGND VGND VPWR VPWR _5963_/B1 sky130_fd_sc_hd__buf_12
X_6089_ _6083_/Y _5240_/B _6084_/Y _4590_/B _6088_/X VGND VGND VPWR VPWR _6096_/C
+ sky130_fd_sc_hd__o221a_2
Xrepeater371 _7011_/B VGND VGND VPWR VPWR _9779_/SET_B sky130_fd_sc_hd__buf_12
XFILLER_45_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_25_csclk clkbuf_2_3_0_csclk/X VGND VGND VPWR VPWR _9652_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_41_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9779_ _9779_/CLK _9779_/D _9779_/SET_B VGND VGND VPWR VPWR _9779_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_13_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput130 usr2_vcc_pwrgood VGND VGND VPWR VPWR _6676_/A sky130_fd_sc_hd__clkbuf_1
Xinput152 wb_adr_i[28] VGND VGND VPWR VPWR _5930_/B sky130_fd_sc_hd__clkbuf_1
Xinput141 wb_adr_i[18] VGND VGND VPWR VPWR _7768_/D sky130_fd_sc_hd__clkbuf_1
Xinput163 wb_adr_i[9] VGND VGND VPWR VPWR _7774_/C sky130_fd_sc_hd__clkbuf_1
Xinput185 wb_dat_i[28] VGND VGND VPWR VPWR _7745_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput174 wb_dat_i[18] VGND VGND VPWR VPWR _7740_/B sky130_fd_sc_hd__clkbuf_1
Xinput196 wb_dat_i[9] VGND VGND VPWR VPWR _7739_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5460_ _5460_/A VGND VGND VPWR VPWR _5460_/Y sky130_fd_sc_hd__inv_2
XFILLER_184_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5391_ _9451_/Q _5384_/A _8840_/X _5384_/Y VGND VGND VPWR VPWR _9451_/D sky130_fd_sc_hd__a22o_1
XFILLER_172_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7130_ _4928_/Y _7124_/X _4771_/Y _7068_/B _7129_/X VGND VGND VPWR VPWR _7131_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_125_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7061_ _7061_/A VGND VGND VPWR VPWR _7068_/A sky130_fd_sc_hd__buf_8
XFILLER_101_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6012_ _6040_/A VGND VGND VPWR VPWR _6013_/A sky130_fd_sc_hd__clkbuf_1
.ends

