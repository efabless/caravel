VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO open_source
  CLASS BLOCK ;
  FOREIGN open_source ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 25.000 ;
END open_source
END LIBRARY

