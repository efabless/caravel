magic
tech sky130A
magscale 1 2
timestamp 1666097791
<< viali >>
rect 1225 18377 1259 18411
rect 18429 18377 18463 18411
rect 4629 18241 4663 18275
rect 5457 18241 5491 18275
rect 10057 18241 10091 18275
rect 1593 18173 1627 18207
rect 1747 18173 1781 18207
rect 2237 18173 2271 18207
rect 2789 18173 2823 18207
rect 7021 18173 7055 18207
rect 7573 18173 7607 18207
rect 8309 18173 8343 18207
rect 9505 18173 9539 18207
rect 10333 18173 10367 18207
rect 11161 18173 11195 18207
rect 12449 18173 12483 18207
rect 12633 18173 12667 18207
rect 17969 18173 18003 18207
rect 5641 18105 5675 18139
rect 6653 18105 6687 18139
rect 8401 18105 8435 18139
rect 9597 18105 9631 18139
rect 11437 18105 11471 18139
rect 1961 18037 1995 18071
rect 2421 18037 2455 18071
rect 2973 18037 3007 18071
rect 4077 18037 4111 18071
rect 4445 18037 4479 18071
rect 4537 18037 4571 18071
rect 5549 18037 5583 18071
rect 6009 18037 6043 18071
rect 10241 18037 10275 18071
rect 10701 18037 10735 18071
rect 12541 18037 12575 18071
rect 17785 18037 17819 18071
rect 3249 17833 3283 17867
rect 11759 17833 11793 17867
rect 949 17765 983 17799
rect 5181 17765 5215 17799
rect 7849 17765 7883 17799
rect 4537 17697 4571 17731
rect 9965 17697 9999 17731
rect 12357 17697 12391 17731
rect 17509 17697 17543 17731
rect 673 17629 707 17663
rect 10333 17629 10367 17663
rect 14749 17629 14783 17663
rect 15117 17629 15151 17663
rect 16589 17629 16623 17663
rect 17601 17629 17635 17663
rect 17785 17629 17819 17663
rect 6469 17561 6503 17595
rect 2421 17493 2455 17527
rect 9321 17493 9355 17527
rect 13645 17493 13679 17527
rect 17141 17493 17175 17527
rect 1685 17289 1719 17323
rect 3617 17289 3651 17323
rect 5825 17289 5859 17323
rect 12449 17289 12483 17323
rect 17969 17289 18003 17323
rect 10563 17221 10597 17255
rect 2513 17153 2547 17187
rect 4353 17153 4387 17187
rect 6561 17153 6595 17187
rect 6929 17153 6963 17187
rect 8769 17153 8803 17187
rect 15577 17153 15611 17187
rect 16221 17153 16255 17187
rect 16497 17153 16531 17187
rect 1593 17085 1627 17119
rect 1777 17085 1811 17119
rect 1915 17085 1949 17119
rect 2053 17085 2087 17119
rect 2329 17085 2363 17119
rect 4077 17085 4111 17119
rect 9137 17085 9171 17119
rect 11161 17085 11195 17119
rect 15209 17085 15243 17119
rect 8355 17017 8389 17051
rect 13783 16949 13817 16983
rect 1685 16745 1719 16779
rect 4813 16745 4847 16779
rect 16037 16745 16071 16779
rect 17233 16745 17267 16779
rect 1593 16677 1627 16711
rect 3700 16677 3734 16711
rect 7021 16677 7055 16711
rect 9597 16677 9631 16711
rect 14749 16677 14783 16711
rect 1869 16609 1903 16643
rect 2973 16609 3007 16643
rect 3157 16609 3191 16643
rect 3433 16609 3467 16643
rect 14105 16609 14139 16643
rect 17601 16609 17635 16643
rect 18429 16609 18463 16643
rect 1777 16541 1811 16575
rect 1961 16541 1995 16575
rect 7849 16541 7883 16575
rect 10241 16541 10275 16575
rect 10517 16541 10551 16575
rect 13829 16541 13863 16575
rect 17693 16541 17727 16575
rect 17785 16541 17819 16575
rect 3157 16405 3191 16439
rect 5733 16405 5767 16439
rect 11989 16405 12023 16439
rect 12357 16405 12391 16439
rect 18245 16405 18279 16439
rect 5549 16201 5583 16235
rect 6837 16201 6871 16235
rect 12449 16201 12483 16235
rect 18429 16201 18463 16235
rect 17693 16133 17727 16167
rect 2053 16065 2087 16099
rect 2237 16065 2271 16099
rect 2789 16065 2823 16099
rect 13829 16065 13863 16099
rect 15945 16065 15979 16099
rect 17233 16065 17267 16099
rect 2881 15997 2915 16031
rect 4261 15997 4295 16031
rect 13553 15997 13587 16031
rect 16129 15997 16163 16031
rect 16221 15997 16255 16031
rect 17325 15997 17359 16031
rect 1961 15929 1995 15963
rect 8125 15929 8159 15963
rect 8769 15929 8803 15963
rect 11161 15929 11195 15963
rect 16589 15929 16623 15963
rect 16773 15929 16807 15963
rect 1593 15861 1627 15895
rect 3249 15861 3283 15895
rect 10057 15861 10091 15895
rect 15301 15861 15335 15895
rect 15945 15861 15979 15895
rect 7205 15657 7239 15691
rect 14749 15657 14783 15691
rect 16589 15657 16623 15691
rect 17233 15657 17267 15691
rect 857 15589 891 15623
rect 4537 15589 4571 15623
rect 10241 15589 10275 15623
rect 11989 15589 12023 15623
rect 12633 15589 12667 15623
rect 581 15521 615 15555
rect 4813 15521 4847 15555
rect 15117 15521 15151 15555
rect 16221 15521 16255 15555
rect 16497 15521 16531 15555
rect 16681 15521 16715 15555
rect 17141 15521 17175 15555
rect 17325 15521 17359 15555
rect 5457 15453 5491 15487
rect 5733 15453 5767 15487
rect 7849 15453 7883 15487
rect 8125 15453 8159 15487
rect 12357 15453 12391 15487
rect 15209 15453 15243 15487
rect 15301 15453 15335 15487
rect 15945 15453 15979 15487
rect 2329 15385 2363 15419
rect 14105 15385 14139 15419
rect 9597 15317 9631 15351
rect 17601 15317 17635 15351
rect 8309 15113 8343 15147
rect 15945 15113 15979 15147
rect 3525 15045 3559 15079
rect 5181 15045 5215 15079
rect 2237 14977 2271 15011
rect 4721 14977 4755 15011
rect 5365 14977 5399 15011
rect 7665 14977 7699 15011
rect 14289 14977 14323 15011
rect 16497 14977 16531 15011
rect 2053 14909 2087 14943
rect 2697 14909 2731 14943
rect 3433 14909 3467 14943
rect 3617 14909 3651 14943
rect 4537 14909 4571 14943
rect 4629 14909 4663 14943
rect 5089 14909 5123 14943
rect 5641 14909 5675 14943
rect 5825 14909 5859 14943
rect 7941 14909 7975 14943
rect 11161 14909 11195 14943
rect 11529 14909 11563 14943
rect 13553 14909 13587 14943
rect 17417 14909 17451 14943
rect 17601 14909 17635 14943
rect 4169 14841 4203 14875
rect 4353 14841 4387 14875
rect 5365 14841 5399 14875
rect 9045 14841 9079 14875
rect 1593 14773 1627 14807
rect 1961 14773 1995 14807
rect 2697 14773 2731 14807
rect 5733 14773 5767 14807
rect 6377 14773 6411 14807
rect 7849 14773 7883 14807
rect 10333 14773 10367 14807
rect 12955 14773 12989 14807
rect 16313 14773 16347 14807
rect 16405 14773 16439 14807
rect 17509 14773 17543 14807
rect 3249 14569 3283 14603
rect 3709 14569 3743 14603
rect 11069 14569 11103 14603
rect 14933 14569 14967 14603
rect 2421 14501 2455 14535
rect 11345 14501 11379 14535
rect 15669 14501 15703 14535
rect 581 14433 615 14467
rect 949 14433 983 14467
rect 3617 14433 3651 14467
rect 5365 14433 5399 14467
rect 5733 14433 5767 14467
rect 7757 14433 7791 14467
rect 10701 14433 10735 14467
rect 12357 14433 12391 14467
rect 12725 14433 12759 14467
rect 15025 14433 15059 14467
rect 15853 14433 15887 14467
rect 15945 14433 15979 14467
rect 17141 14433 17175 14467
rect 17601 14433 17635 14467
rect 17877 14433 17911 14467
rect 18245 14433 18279 14467
rect 3801 14365 3835 14399
rect 8125 14365 8159 14399
rect 10517 14365 10551 14399
rect 15485 14365 15519 14399
rect 16037 14365 16071 14399
rect 17233 14365 17267 14399
rect 18061 14297 18095 14331
rect 7159 14229 7193 14263
rect 9551 14229 9585 14263
rect 14151 14229 14185 14263
rect 17325 14229 17359 14263
rect 17463 14229 17497 14263
rect 17969 14229 18003 14263
rect 18245 14229 18279 14263
rect 2053 14025 2087 14059
rect 5641 14025 5675 14059
rect 8769 14025 8803 14059
rect 10253 14025 10287 14059
rect 17785 14025 17819 14059
rect 12725 13957 12759 13991
rect 2513 13889 2547 13923
rect 2697 13889 2731 13923
rect 10517 13889 10551 13923
rect 11897 13889 11931 13923
rect 14013 13889 14047 13923
rect 6745 13821 6779 13855
rect 7113 13821 7147 13855
rect 7481 13821 7515 13855
rect 11805 13821 11839 13855
rect 11989 13821 12023 13855
rect 12265 13821 12299 13855
rect 12633 13821 12667 13855
rect 12817 13821 12851 13855
rect 13093 13821 13127 13855
rect 15025 13821 15059 13855
rect 15301 13821 15335 13855
rect 15945 13821 15979 13855
rect 17416 13821 17450 13855
rect 17509 13821 17543 13855
rect 17969 13821 18003 13855
rect 18429 13821 18463 13855
rect 2421 13753 2455 13787
rect 6929 13753 6963 13787
rect 7757 13753 7791 13787
rect 8217 13753 8251 13787
rect 14105 13753 14139 13787
rect 14197 13753 14231 13787
rect 16221 13753 16255 13787
rect 6009 13685 6043 13719
rect 14565 13685 14599 13719
rect 17141 13685 17175 13719
rect 7803 13481 7837 13515
rect 10701 13481 10735 13515
rect 13093 13481 13127 13515
rect 15669 13481 15703 13515
rect 11989 13413 12023 13447
rect 3433 13345 3467 13379
rect 3700 13345 3734 13379
rect 5457 13345 5491 13379
rect 6193 13345 6227 13379
rect 6377 13345 6411 13379
rect 6653 13345 6687 13379
rect 7021 13345 7055 13379
rect 14381 13345 14415 13379
rect 14749 13345 14783 13379
rect 15209 13345 15243 13379
rect 15577 13345 15611 13379
rect 15761 13345 15795 13379
rect 16405 13345 16439 13379
rect 5733 13277 5767 13311
rect 6837 13277 6871 13311
rect 9229 13277 9263 13311
rect 9597 13277 9631 13311
rect 14841 13277 14875 13311
rect 4813 13209 4847 13243
rect 6929 13209 6963 13243
rect 5549 13141 5583 13175
rect 5641 13141 5675 13175
rect 6377 13141 6411 13175
rect 16129 13141 16163 13175
rect 4353 12937 4387 12971
rect 4997 12937 5031 12971
rect 7481 12937 7515 12971
rect 13553 12937 13587 12971
rect 17969 12937 18003 12971
rect 7757 12801 7791 12835
rect 10517 12801 10551 12835
rect 14197 12801 14231 12835
rect 16497 12801 16531 12835
rect 4169 12733 4203 12767
rect 4353 12733 4387 12767
rect 4721 12733 4755 12767
rect 4813 12733 4847 12767
rect 6653 12733 6687 12767
rect 6929 12733 6963 12767
rect 7113 12733 7147 12767
rect 7481 12733 7515 12767
rect 7941 12733 7975 12767
rect 11161 12733 11195 12767
rect 11529 12733 11563 12767
rect 13737 12733 13771 12767
rect 13921 12733 13955 12767
rect 16221 12733 16255 12767
rect 5641 12665 5675 12699
rect 10241 12665 10275 12699
rect 12955 12665 12989 12699
rect 14464 12665 14498 12699
rect 5365 12597 5399 12631
rect 8769 12597 8803 12631
rect 15577 12597 15611 12631
rect 7849 12393 7883 12427
rect 10793 12393 10827 12427
rect 17233 12393 17267 12427
rect 3157 12325 3191 12359
rect 3617 12325 3651 12359
rect 11253 12325 11287 12359
rect 14105 12325 14139 12359
rect 1041 12257 1075 12291
rect 1308 12257 1342 12291
rect 2789 12257 2823 12291
rect 2882 12257 2916 12291
rect 3433 12257 3467 12291
rect 3709 12257 3743 12291
rect 6929 12257 6963 12291
rect 10609 12257 10643 12291
rect 10793 12257 10827 12291
rect 11621 12257 11655 12291
rect 12817 12257 12851 12291
rect 13737 12257 13771 12291
rect 15209 12257 15243 12291
rect 15393 12257 15427 12291
rect 15853 12257 15887 12291
rect 16313 12257 16347 12291
rect 5181 12189 5215 12223
rect 9321 12189 9355 12223
rect 9597 12189 9631 12223
rect 13921 12189 13955 12223
rect 14749 12189 14783 12223
rect 15669 12189 15703 12223
rect 16589 12189 16623 12223
rect 2421 12121 2455 12155
rect 13829 12121 13863 12155
rect 15393 12121 15427 12155
rect 3709 12053 3743 12087
rect 12449 12053 12483 12087
rect 16037 12053 16071 12087
rect 16405 12053 16439 12087
rect 16497 12053 16531 12087
rect 4261 11849 4295 11883
rect 4721 11849 4755 11883
rect 5549 11849 5583 11883
rect 7113 11849 7147 11883
rect 8217 11849 8251 11883
rect 2605 11781 2639 11815
rect 11161 11781 11195 11815
rect 7573 11713 7607 11747
rect 7665 11713 7699 11747
rect 10517 11713 10551 11747
rect 11529 11713 11563 11747
rect 16129 11713 16163 11747
rect 2237 11645 2271 11679
rect 2391 11645 2425 11679
rect 4629 11645 4663 11679
rect 4905 11645 4939 11679
rect 4997 11645 5031 11679
rect 5733 11645 5767 11679
rect 5917 11645 5951 11679
rect 6009 11645 6043 11679
rect 6837 11645 6871 11679
rect 7481 11645 7515 11679
rect 11345 11645 11379 11679
rect 11437 11645 11471 11679
rect 11621 11645 11655 11679
rect 15577 11645 15611 11679
rect 16497 11645 16531 11679
rect 6561 11577 6595 11611
rect 10241 11577 10275 11611
rect 5181 11509 5215 11543
rect 8769 11509 8803 11543
rect 14289 11509 14323 11543
rect 17923 11509 17957 11543
rect 1961 11305 1995 11339
rect 6929 11305 6963 11339
rect 8309 11305 8343 11339
rect 10885 11305 10919 11339
rect 13737 11305 13771 11339
rect 14749 11305 14783 11339
rect 15209 11305 15243 11339
rect 16129 11305 16163 11339
rect 16589 11305 16623 11339
rect 18245 11305 18279 11339
rect 5457 11237 5491 11271
rect 9597 11237 9631 11271
rect 16405 11237 16439 11271
rect 17141 11237 17175 11271
rect 581 11169 615 11203
rect 848 11169 882 11203
rect 2973 11169 3007 11203
rect 5181 11169 5215 11203
rect 11069 11169 11103 11203
rect 11161 11169 11195 11203
rect 11437 11169 11471 11203
rect 13829 11169 13863 11203
rect 15117 11169 15151 11203
rect 15853 11169 15887 11203
rect 16681 11169 16715 11203
rect 17509 11169 17543 11203
rect 17969 11169 18003 11203
rect 18429 11169 18463 11203
rect 2881 11101 2915 11135
rect 10977 11101 11011 11135
rect 11253 11101 11287 11135
rect 14013 11101 14047 11135
rect 15301 11101 15335 11135
rect 16129 11101 16163 11135
rect 3341 11033 3375 11067
rect 15945 11033 15979 11067
rect 16405 11033 16439 11067
rect 4629 10965 4663 10999
rect 13369 10965 13403 10999
rect 12909 10761 12943 10795
rect 17969 10761 18003 10795
rect 4721 10693 4755 10727
rect 5273 10693 5307 10727
rect 14841 10693 14875 10727
rect 4353 10625 4387 10659
rect 14381 10625 14415 10659
rect 16221 10625 16255 10659
rect 1133 10557 1167 10591
rect 1225 10557 1259 10591
rect 1593 10557 1627 10591
rect 1961 10557 1995 10591
rect 4445 10557 4479 10591
rect 4721 10557 4755 10591
rect 4905 10557 4939 10591
rect 10333 10557 10367 10591
rect 12449 10557 12483 10591
rect 13001 10557 13035 10591
rect 14473 10557 14507 10591
rect 4169 10489 4203 10523
rect 6377 10489 6411 10523
rect 16497 10489 16531 10523
rect 3387 10421 3421 10455
rect 4445 10421 4479 10455
rect 10333 10421 10367 10455
rect 12541 10421 12575 10455
rect 12725 10421 12759 10455
rect 1593 10217 1627 10251
rect 6469 10217 6503 10251
rect 7205 10217 7239 10251
rect 12449 10217 12483 10251
rect 13093 10217 13127 10251
rect 17141 10217 17175 10251
rect 2789 10149 2823 10183
rect 4537 10149 4571 10183
rect 1961 10081 1995 10115
rect 2053 10081 2087 10115
rect 6377 10081 6411 10115
rect 6561 10081 6595 10115
rect 7021 10081 7055 10115
rect 7573 10081 7607 10115
rect 10149 10081 10183 10115
rect 10517 10081 10551 10115
rect 12724 10081 12758 10115
rect 12817 10081 12851 10115
rect 13093 10081 13127 10115
rect 13277 10081 13311 10115
rect 17345 10081 17379 10115
rect 17463 10081 17497 10115
rect 17693 10081 17727 10115
rect 2237 10013 2271 10047
rect 6837 10013 6871 10047
rect 7941 10013 7975 10047
rect 11943 10013 11977 10047
rect 17601 9945 17635 9979
rect 9367 9877 9401 9911
rect 16037 9877 16071 9911
rect 2881 9605 2915 9639
rect 8309 9605 8343 9639
rect 8769 9605 8803 9639
rect 3433 9537 3467 9571
rect 8401 9537 8435 9571
rect 2513 9469 2547 9503
rect 3249 9469 3283 9503
rect 5733 9469 5767 9503
rect 8125 9469 8159 9503
rect 8217 9469 8251 9503
rect 9045 9469 9079 9503
rect 14289 9469 14323 9503
rect 14657 9469 14691 9503
rect 15025 9469 15059 9503
rect 2237 9401 2271 9435
rect 3341 9401 3375 9435
rect 8769 9401 8803 9435
rect 4813 9333 4847 9367
rect 5457 9333 5491 9367
rect 8953 9333 8987 9367
rect 12081 9333 12115 9367
rect 12449 9333 12483 9367
rect 15025 9333 15059 9367
rect 1777 9129 1811 9163
rect 3157 9129 3191 9163
rect 3617 9129 3651 9163
rect 4169 9129 4203 9163
rect 17325 9129 17359 9163
rect 18245 9129 18279 9163
rect 14105 9061 14139 9095
rect 15393 9061 15427 9095
rect 17233 9061 17267 9095
rect 1685 8993 1719 9027
rect 3525 8993 3559 9027
rect 4353 8993 4387 9027
rect 5273 8993 5307 9027
rect 12541 8993 12575 9027
rect 12633 8993 12667 9027
rect 12725 8993 12759 9027
rect 14381 8993 14415 9027
rect 14749 8993 14783 9027
rect 14903 8993 14937 9027
rect 15669 8993 15703 9027
rect 17141 8993 17175 9027
rect 17417 8993 17451 9027
rect 18429 8993 18463 9027
rect 1961 8925 1995 8959
rect 3801 8925 3835 8959
rect 4629 8925 4663 8959
rect 5641 8925 5675 8959
rect 10241 8925 10275 8959
rect 10517 8925 10551 8959
rect 11989 8925 12023 8959
rect 15393 8925 15427 8959
rect 14289 8857 14323 8891
rect 14381 8857 14415 8891
rect 15117 8857 15151 8891
rect 17969 8857 18003 8891
rect 1317 8789 1351 8823
rect 4537 8789 4571 8823
rect 7067 8789 7101 8823
rect 12357 8789 12391 8823
rect 15577 8789 15611 8823
rect 3065 8585 3099 8619
rect 3985 8585 4019 8619
rect 4997 8585 5031 8619
rect 5365 8585 5399 8619
rect 11253 8585 11287 8619
rect 17969 8585 18003 8619
rect 13553 8517 13587 8551
rect 14565 8517 14599 8551
rect 16313 8517 16347 8551
rect 2973 8449 3007 8483
rect 11161 8449 11195 8483
rect 14105 8449 14139 8483
rect 3249 8381 3283 8415
rect 3433 8381 3467 8415
rect 4169 8381 4203 8415
rect 4445 8381 4479 8415
rect 5273 8381 5307 8415
rect 5457 8381 5491 8415
rect 6837 8381 6871 8415
rect 11345 8381 11379 8415
rect 11437 8381 11471 8415
rect 12357 8381 12391 8415
rect 12449 8381 12483 8415
rect 14013 8381 14047 8415
rect 15945 8381 15979 8415
rect 16099 8381 16133 8415
rect 16589 8381 16623 8415
rect 6377 8313 6411 8347
rect 16845 8313 16879 8347
rect 4353 8245 4387 8279
rect 13921 8245 13955 8279
rect 5365 8041 5399 8075
rect 14749 8041 14783 8075
rect 15117 8041 15151 8075
rect 17509 8041 17543 8075
rect 857 7973 891 8007
rect 4537 7973 4571 8007
rect 12817 7973 12851 8007
rect 14381 7973 14415 8007
rect 15209 7973 15243 8007
rect 15761 7973 15795 8007
rect 581 7905 615 7939
rect 2973 7905 3007 7939
rect 7573 7905 7607 7939
rect 10701 7905 10735 7939
rect 10793 7905 10827 7939
rect 10977 7905 11011 7939
rect 17141 7905 17175 7939
rect 17234 7905 17268 7939
rect 2329 7837 2363 7871
rect 5549 7837 5583 7871
rect 5641 7837 5675 7871
rect 5733 7837 5767 7871
rect 5825 7837 5859 7871
rect 7941 7837 7975 7871
rect 15301 7837 15335 7871
rect 10977 7769 11011 7803
rect 9321 7701 9355 7735
rect 3249 7497 3283 7531
rect 5641 7497 5675 7531
rect 11345 7497 11379 7531
rect 17785 7497 17819 7531
rect 9045 7429 9079 7463
rect 9597 7429 9631 7463
rect 13645 7429 13679 7463
rect 14105 7429 14139 7463
rect 2237 7361 2271 7395
rect 5089 7361 5123 7395
rect 5457 7361 5491 7395
rect 8769 7361 8803 7395
rect 9229 7361 9263 7395
rect 11161 7361 11195 7395
rect 11897 7361 11931 7395
rect 14657 7361 14691 7395
rect 16405 7361 16439 7395
rect 1961 7293 1995 7327
rect 3157 7293 3191 7327
rect 3985 7293 4019 7327
rect 4169 7293 4203 7327
rect 5549 7293 5583 7327
rect 6929 7293 6963 7327
rect 7113 7293 7147 7327
rect 8861 7293 8895 7327
rect 9045 7293 9079 7327
rect 9597 7293 9631 7327
rect 9781 7293 9815 7327
rect 11437 7293 11471 7327
rect 12081 7293 12115 7327
rect 12173 7293 12207 7327
rect 12301 7293 12335 7327
rect 13737 7293 13771 7327
rect 14565 7293 14599 7327
rect 4353 7225 4387 7259
rect 5273 7225 5307 7259
rect 5365 7225 5399 7259
rect 7757 7225 7791 7259
rect 16650 7225 16684 7259
rect 1593 7157 1627 7191
rect 2053 7157 2087 7191
rect 7113 7157 7147 7191
rect 7665 7157 7699 7191
rect 8309 7157 8343 7191
rect 9137 7157 9171 7191
rect 11161 7157 11195 7191
rect 14473 7157 14507 7191
rect 2329 6953 2363 6987
rect 2789 6953 2823 6987
rect 3157 6953 3191 6987
rect 8217 6953 8251 6987
rect 14749 6953 14783 6987
rect 4169 6885 4203 6919
rect 581 6817 615 6851
rect 6469 6817 6503 6851
rect 6744 6817 6778 6851
rect 6837 6817 6871 6851
rect 7665 6817 7699 6851
rect 7941 6817 7975 6851
rect 8493 6817 8527 6851
rect 8677 6817 8711 6851
rect 12909 6817 12943 6851
rect 13369 6817 13403 6851
rect 13737 6817 13771 6851
rect 15117 6817 15151 6851
rect 17233 6817 17267 6851
rect 17969 6817 18003 6851
rect 18429 6817 18463 6851
rect 857 6749 891 6783
rect 3249 6749 3283 6783
rect 3433 6749 3467 6783
rect 4261 6749 4295 6783
rect 4353 6749 4387 6783
rect 7573 6749 7607 6783
rect 8033 6749 8067 6783
rect 10149 6749 10183 6783
rect 10425 6749 10459 6783
rect 11897 6749 11931 6783
rect 13461 6749 13495 6783
rect 15209 6749 15243 6783
rect 15301 6749 15335 6783
rect 3801 6681 3835 6715
rect 12633 6681 12667 6715
rect 18245 6681 18279 6715
rect 8585 6613 8619 6647
rect 8953 6613 8987 6647
rect 17325 6613 17359 6647
rect 2237 6409 2271 6443
rect 2697 6409 2731 6443
rect 5825 6409 5859 6443
rect 14289 6409 14323 6443
rect 14933 6409 14967 6443
rect 2053 6273 2087 6307
rect 4077 6273 4111 6307
rect 4721 6273 4755 6307
rect 8125 6273 8159 6307
rect 16129 6273 16163 6307
rect 1961 6205 1995 6239
rect 2973 6205 3007 6239
rect 4445 6205 4479 6239
rect 4997 6205 5031 6239
rect 5457 6205 5491 6239
rect 7757 6205 7791 6239
rect 7849 6205 7883 6239
rect 12817 6205 12851 6239
rect 14749 6205 14783 6239
rect 16497 6205 16531 6239
rect 6377 6137 6411 6171
rect 8217 6137 8251 6171
rect 15577 6137 15611 6171
rect 17969 6137 18003 6171
rect 7573 6069 7607 6103
rect 12081 6069 12115 6103
rect 12909 6069 12943 6103
rect 4169 5865 4203 5899
rect 5365 5865 5399 5899
rect 17141 5865 17175 5899
rect 5181 5797 5215 5831
rect 8033 5797 8067 5831
rect 18061 5797 18095 5831
rect 1869 5729 1903 5763
rect 4261 5729 4295 5763
rect 5457 5729 5491 5763
rect 6193 5729 6227 5763
rect 7757 5729 7791 5763
rect 13093 5729 13127 5763
rect 13737 5729 13771 5763
rect 13830 5729 13864 5763
rect 15301 5729 15335 5763
rect 15485 5729 15519 5763
rect 15761 5729 15795 5763
rect 15945 5729 15979 5763
rect 16221 5729 16255 5763
rect 16405 5729 16439 5763
rect 16681 5729 16715 5763
rect 17325 5729 17359 5763
rect 17509 5729 17543 5763
rect 17601 5729 17635 5763
rect 6285 5661 6319 5695
rect 6469 5661 6503 5695
rect 10057 5661 10091 5695
rect 10333 5661 10367 5695
rect 13185 5661 13219 5695
rect 13277 5661 13311 5695
rect 15393 5661 15427 5695
rect 14105 5593 14139 5627
rect 15853 5593 15887 5627
rect 17417 5593 17451 5627
rect 2053 5525 2087 5559
rect 5181 5525 5215 5559
rect 6377 5525 6411 5559
rect 9505 5525 9539 5559
rect 11805 5525 11839 5559
rect 12449 5525 12483 5559
rect 12725 5525 12759 5559
rect 11161 5321 11195 5355
rect 17877 5321 17911 5355
rect 12265 5253 12299 5287
rect 12633 5253 12667 5287
rect 1685 5185 1719 5219
rect 4261 5185 4295 5219
rect 6377 5185 6411 5219
rect 8401 5185 8435 5219
rect 11805 5185 11839 5219
rect 13185 5185 13219 5219
rect 16129 5185 16163 5219
rect 2053 5117 2087 5151
rect 10425 5117 10459 5151
rect 13553 5117 13587 5151
rect 4537 5049 4571 5083
rect 6653 5049 6687 5083
rect 11529 5049 11563 5083
rect 13829 5049 13863 5083
rect 15577 5049 15611 5083
rect 16405 5049 16439 5083
rect 3479 4981 3513 5015
rect 6009 4981 6043 5015
rect 10149 4981 10183 5015
rect 11621 4981 11655 5015
rect 4537 4777 4571 4811
rect 6561 4777 6595 4811
rect 14749 4777 14783 4811
rect 16037 4777 16071 4811
rect 581 4641 615 4675
rect 3341 4641 3375 4675
rect 3433 4641 3467 4675
rect 3525 4641 3559 4675
rect 4813 4641 4847 4675
rect 6837 4641 6871 4675
rect 9965 4641 9999 4675
rect 14105 4641 14139 4675
rect 14933 4641 14967 4675
rect 15025 4641 15059 4675
rect 857 4573 891 4607
rect 2329 4573 2363 4607
rect 4537 4573 4571 4607
rect 4721 4573 4755 4607
rect 6561 4573 6595 4607
rect 10333 4573 10367 4607
rect 13829 4573 13863 4607
rect 14749 4573 14783 4607
rect 3157 4437 3191 4471
rect 6745 4437 6779 4471
rect 11759 4437 11793 4471
rect 12357 4437 12391 4471
rect 949 4233 983 4267
rect 4813 4233 4847 4267
rect 11161 4233 11195 4267
rect 14657 4233 14691 4267
rect 17325 4165 17359 4199
rect 857 4097 891 4131
rect 1041 4097 1075 4131
rect 8309 4097 8343 4131
rect 9321 4097 9355 4131
rect 11805 4097 11839 4131
rect 12357 4097 12391 4131
rect 14749 4097 14783 4131
rect 16497 4097 16531 4131
rect 17049 4097 17083 4131
rect 17417 4097 17451 4131
rect 765 4029 799 4063
rect 4445 4029 4479 4063
rect 4537 4029 4571 4063
rect 4629 4029 4663 4063
rect 11529 4029 11563 4063
rect 14473 4029 14507 4063
rect 14565 4029 14599 4063
rect 16405 4029 16439 4063
rect 17233 4029 17267 4063
rect 17509 4029 17543 4063
rect 8033 3961 8067 3995
rect 9229 3961 9263 3995
rect 12541 3961 12575 3995
rect 16313 3961 16347 3995
rect 7665 3893 7699 3927
rect 8125 3893 8159 3927
rect 8769 3893 8803 3927
rect 9137 3893 9171 3927
rect 11621 3893 11655 3927
rect 12633 3893 12667 3927
rect 13001 3893 13035 3927
rect 15945 3893 15979 3927
rect 1869 3689 1903 3723
rect 5273 3689 5307 3723
rect 6101 3689 6135 3723
rect 6469 3689 6503 3723
rect 8493 3689 8527 3723
rect 14197 3689 14231 3723
rect 14749 3689 14783 3723
rect 16313 3689 16347 3723
rect 17417 3689 17451 3723
rect 18245 3689 18279 3723
rect 1685 3621 1719 3655
rect 3157 3621 3191 3655
rect 6929 3621 6963 3655
rect 1593 3553 1627 3587
rect 2145 3553 2179 3587
rect 3432 3553 3466 3587
rect 3525 3553 3559 3587
rect 3801 3553 3835 3587
rect 3985 3553 4019 3587
rect 5181 3553 5215 3587
rect 6837 3553 6871 3587
rect 11253 3553 11287 3587
rect 11437 3553 11471 3587
rect 13737 3553 13771 3587
rect 14013 3553 14047 3587
rect 16129 3553 16163 3587
rect 16405 3553 16439 3587
rect 16589 3553 16623 3587
rect 17509 3553 17543 3587
rect 17693 3553 17727 3587
rect 18429 3553 18463 3587
rect 3893 3485 3927 3519
rect 7021 3485 7055 3519
rect 11437 3417 11471 3451
rect 13829 3417 13863 3451
rect 2053 3349 2087 3383
rect 17233 3349 17267 3383
rect 857 3145 891 3179
rect 4997 3145 5031 3179
rect 6653 3145 6687 3179
rect 6929 3145 6963 3179
rect 8769 3145 8803 3179
rect 11529 3145 11563 3179
rect 12449 3145 12483 3179
rect 14841 3145 14875 3179
rect 17141 3145 17175 3179
rect 18429 3145 18463 3179
rect 10333 3077 10367 3111
rect 5641 3009 5675 3043
rect 7389 3009 7423 3043
rect 7573 3009 7607 3043
rect 9321 3009 9355 3043
rect 11161 3009 11195 3043
rect 11621 3009 11655 3043
rect 13001 3009 13035 3043
rect 15393 3009 15427 3043
rect 17693 3009 17727 3043
rect 765 2941 799 2975
rect 7297 2941 7331 2975
rect 9229 2941 9263 2975
rect 10517 2941 10551 2975
rect 10793 2941 10827 2975
rect 11345 2941 11379 2975
rect 15301 2941 15335 2975
rect 5457 2873 5491 2907
rect 10701 2873 10735 2907
rect 12817 2873 12851 2907
rect 16865 2873 16899 2907
rect 17601 2873 17635 2907
rect 5365 2805 5399 2839
rect 9137 2805 9171 2839
rect 12909 2805 12943 2839
rect 15209 2805 15243 2839
rect 17509 2805 17543 2839
rect 581 2601 615 2635
rect 1593 2601 1627 2635
rect 2053 2601 2087 2635
rect 2789 2601 2823 2635
rect 5365 2601 5399 2635
rect 5825 2601 5859 2635
rect 8217 2601 8251 2635
rect 13185 2601 13219 2635
rect 14289 2601 14323 2635
rect 15209 2601 15243 2635
rect 15577 2601 15611 2635
rect 17233 2601 17267 2635
rect 17693 2601 17727 2635
rect 7849 2533 7883 2567
rect 8677 2533 8711 2567
rect 15669 2533 15703 2567
rect 16773 2533 16807 2567
rect 949 2465 983 2499
rect 1961 2465 1995 2499
rect 5733 2465 5767 2499
rect 8585 2465 8619 2499
rect 13185 2465 13219 2499
rect 13737 2465 13771 2499
rect 13921 2465 13955 2499
rect 17601 2465 17635 2499
rect 1041 2397 1075 2431
rect 1225 2397 1259 2431
rect 2145 2397 2179 2431
rect 5917 2397 5951 2431
rect 8769 2397 8803 2431
rect 13461 2397 13495 2431
rect 15853 2397 15887 2431
rect 17785 2397 17819 2431
rect 13277 2329 13311 2363
rect 13737 2261 13771 2295
rect 1593 2057 1627 2091
rect 2881 2057 2915 2091
rect 4077 2057 4111 2091
rect 12173 2057 12207 2091
rect 16681 2057 16715 2091
rect 11897 1989 11931 2023
rect 3341 1921 3375 1955
rect 3525 1921 3559 1955
rect 7205 1921 7239 1955
rect 9229 1921 9263 1955
rect 11345 1921 11379 1955
rect 12633 1921 12667 1955
rect 12725 1921 12759 1955
rect 14013 1921 14047 1955
rect 16129 1921 16163 1955
rect 4353 1853 4387 1887
rect 4629 1853 4663 1887
rect 5181 1853 5215 1887
rect 7389 1853 7423 1887
rect 7665 1853 7699 1887
rect 9597 1853 9631 1887
rect 13921 1853 13955 1887
rect 15025 1853 15059 1887
rect 15301 1853 15335 1887
rect 15393 1853 15427 1887
rect 15577 1853 15611 1887
rect 17693 1853 17727 1887
rect 17969 1853 18003 1887
rect 11437 1785 11471 1819
rect 3249 1717 3283 1751
rect 4445 1717 4479 1751
rect 7573 1717 7607 1751
rect 11529 1717 11563 1751
rect 12541 1717 12575 1751
rect 13553 1717 13587 1751
rect 16221 1717 16255 1751
rect 16313 1717 16347 1751
rect 18429 1717 18463 1751
rect 2237 1513 2271 1547
rect 3157 1513 3191 1547
rect 5641 1513 5675 1547
rect 11713 1513 11747 1547
rect 13185 1513 13219 1547
rect 14013 1513 14047 1547
rect 15485 1513 15519 1547
rect 17417 1513 17451 1547
rect 18061 1513 18095 1547
rect 3249 1445 3283 1479
rect 3801 1445 3835 1479
rect 4813 1445 4847 1479
rect 7573 1445 7607 1479
rect 10241 1445 10275 1479
rect 15761 1445 15795 1479
rect 2421 1377 2455 1411
rect 4537 1377 4571 1411
rect 5273 1377 5307 1411
rect 5366 1377 5400 1411
rect 6837 1377 6871 1411
rect 8033 1377 8067 1411
rect 9075 1377 9109 1411
rect 9229 1377 9263 1411
rect 9965 1377 9999 1411
rect 10977 1377 11011 1411
rect 11805 1377 11839 1411
rect 13369 1377 13403 1411
rect 13553 1377 13587 1411
rect 15117 1377 15151 1411
rect 15853 1377 15887 1411
rect 17631 1377 17665 1411
rect 17785 1377 17819 1411
rect 18061 1377 18095 1411
rect 18337 1377 18371 1411
rect 3433 1309 3467 1343
rect 4813 1309 4847 1343
rect 6745 1309 6779 1343
rect 10885 1309 10919 1343
rect 13645 1309 13679 1343
rect 15025 1309 15059 1343
rect 2789 1241 2823 1275
rect 7205 1241 7239 1275
rect 9965 1241 9999 1275
rect 10057 1241 10091 1275
rect 11345 1241 11379 1275
rect 18153 1241 18187 1275
rect 4629 1173 4663 1207
rect 9045 1173 9079 1207
rect 3249 969 3283 1003
rect 5273 969 5307 1003
rect 8953 969 8987 1003
rect 17509 969 17543 1003
rect 17601 969 17635 1003
rect 5365 901 5399 935
rect 9045 901 9079 935
rect 2881 833 2915 867
rect 8861 833 8895 867
rect 17417 833 17451 867
rect 2973 765 3007 799
rect 5181 765 5215 799
rect 5457 765 5491 799
rect 9137 765 9171 799
rect 17693 765 17727 799
<< metal1 >>
rect 184 18522 18860 18544
rect 184 18470 1556 18522
rect 1608 18470 1620 18522
rect 1672 18470 1684 18522
rect 1736 18470 1748 18522
rect 1800 18470 1812 18522
rect 1864 18470 4656 18522
rect 4708 18470 4720 18522
rect 4772 18470 4784 18522
rect 4836 18470 4848 18522
rect 4900 18470 4912 18522
rect 4964 18470 7756 18522
rect 7808 18470 7820 18522
rect 7872 18470 7884 18522
rect 7936 18470 7948 18522
rect 8000 18470 8012 18522
rect 8064 18470 10856 18522
rect 10908 18470 10920 18522
rect 10972 18470 10984 18522
rect 11036 18470 11048 18522
rect 11100 18470 11112 18522
rect 11164 18470 13956 18522
rect 14008 18470 14020 18522
rect 14072 18470 14084 18522
rect 14136 18470 14148 18522
rect 14200 18470 14212 18522
rect 14264 18470 17056 18522
rect 17108 18470 17120 18522
rect 17172 18470 17184 18522
rect 17236 18470 17248 18522
rect 17300 18470 17312 18522
rect 17364 18470 18860 18522
rect 184 18448 18860 18470
rect 1213 18411 1271 18417
rect 1213 18377 1225 18411
rect 1259 18408 1271 18411
rect 1394 18408 1400 18420
rect 1259 18380 1400 18408
rect 1259 18377 1271 18380
rect 1213 18371 1271 18377
rect 1394 18368 1400 18380
rect 1452 18368 1458 18420
rect 18414 18408 18420 18420
rect 18375 18380 18420 18408
rect 18414 18368 18420 18380
rect 18472 18368 18478 18420
rect 1412 18272 1440 18368
rect 11146 18340 11152 18352
rect 8220 18312 11152 18340
rect 1412 18244 2268 18272
rect 1394 18164 1400 18216
rect 1452 18204 1458 18216
rect 1581 18207 1639 18213
rect 1581 18204 1593 18207
rect 1452 18176 1593 18204
rect 1452 18164 1458 18176
rect 1581 18173 1593 18176
rect 1627 18173 1639 18207
rect 1581 18167 1639 18173
rect 1735 18207 1793 18213
rect 1735 18173 1747 18207
rect 1781 18204 1793 18207
rect 1946 18204 1952 18216
rect 1781 18176 1952 18204
rect 1781 18173 1793 18176
rect 1735 18167 1793 18173
rect 1946 18164 1952 18176
rect 2004 18164 2010 18216
rect 2240 18213 2268 18244
rect 4430 18232 4436 18284
rect 4488 18272 4494 18284
rect 4617 18275 4675 18281
rect 4617 18272 4629 18275
rect 4488 18244 4629 18272
rect 4488 18232 4494 18244
rect 4617 18241 4629 18244
rect 4663 18241 4675 18275
rect 4617 18235 4675 18241
rect 5445 18275 5503 18281
rect 5445 18241 5457 18275
rect 5491 18272 5503 18275
rect 5718 18272 5724 18284
rect 5491 18244 5724 18272
rect 5491 18241 5503 18244
rect 5445 18235 5503 18241
rect 5718 18232 5724 18244
rect 5776 18232 5782 18284
rect 2225 18207 2283 18213
rect 2225 18173 2237 18207
rect 2271 18173 2283 18207
rect 2777 18207 2835 18213
rect 2777 18204 2789 18207
rect 2225 18167 2283 18173
rect 2424 18176 2789 18204
rect 1210 18028 1216 18080
rect 1268 18068 1274 18080
rect 2424 18077 2452 18176
rect 2777 18173 2789 18176
rect 2823 18173 2835 18207
rect 7009 18207 7067 18213
rect 2777 18167 2835 18173
rect 2976 18176 6960 18204
rect 2976 18080 3004 18176
rect 5442 18096 5448 18148
rect 5500 18136 5506 18148
rect 5629 18139 5687 18145
rect 5629 18136 5641 18139
rect 5500 18108 5641 18136
rect 5500 18096 5506 18108
rect 5629 18105 5641 18108
rect 5675 18105 5687 18139
rect 5629 18099 5687 18105
rect 6546 18096 6552 18148
rect 6604 18136 6610 18148
rect 6641 18139 6699 18145
rect 6641 18136 6653 18139
rect 6604 18108 6653 18136
rect 6604 18096 6610 18108
rect 6641 18105 6653 18108
rect 6687 18105 6699 18139
rect 6932 18136 6960 18176
rect 7009 18173 7021 18207
rect 7055 18204 7067 18207
rect 7098 18204 7104 18216
rect 7055 18176 7104 18204
rect 7055 18173 7067 18176
rect 7009 18167 7067 18173
rect 7098 18164 7104 18176
rect 7156 18164 7162 18216
rect 7282 18164 7288 18216
rect 7340 18204 7346 18216
rect 7561 18207 7619 18213
rect 7561 18204 7573 18207
rect 7340 18176 7573 18204
rect 7340 18164 7346 18176
rect 7561 18173 7573 18176
rect 7607 18173 7619 18207
rect 7561 18167 7619 18173
rect 8220 18136 8248 18312
rect 11146 18300 11152 18312
rect 11204 18300 11210 18352
rect 9674 18232 9680 18284
rect 9732 18272 9738 18284
rect 10045 18275 10103 18281
rect 10045 18272 10057 18275
rect 9732 18244 10057 18272
rect 9732 18232 9738 18244
rect 10045 18241 10057 18244
rect 10091 18241 10103 18275
rect 16022 18272 16028 18284
rect 10045 18235 10103 18241
rect 10336 18244 16028 18272
rect 10336 18213 10364 18244
rect 16022 18232 16028 18244
rect 16080 18232 16086 18284
rect 8297 18207 8355 18213
rect 8297 18173 8309 18207
rect 8343 18204 8355 18207
rect 9493 18207 9551 18213
rect 9493 18204 9505 18207
rect 8343 18176 9505 18204
rect 8343 18173 8355 18176
rect 8297 18167 8355 18173
rect 9493 18173 9505 18176
rect 9539 18204 9551 18207
rect 10321 18207 10379 18213
rect 9539 18176 10088 18204
rect 9539 18173 9551 18176
rect 9493 18167 9551 18173
rect 8386 18136 8392 18148
rect 6932 18108 8248 18136
rect 8347 18108 8392 18136
rect 6641 18099 6699 18105
rect 1949 18071 2007 18077
rect 1949 18068 1961 18071
rect 1268 18040 1961 18068
rect 1268 18028 1274 18040
rect 1949 18037 1961 18040
rect 1995 18037 2007 18071
rect 1949 18031 2007 18037
rect 2409 18071 2467 18077
rect 2409 18037 2421 18071
rect 2455 18037 2467 18071
rect 2958 18068 2964 18080
rect 2919 18040 2964 18068
rect 2409 18031 2467 18037
rect 2958 18028 2964 18040
rect 3016 18028 3022 18080
rect 4062 18068 4068 18080
rect 4023 18040 4068 18068
rect 4062 18028 4068 18040
rect 4120 18028 4126 18080
rect 4338 18028 4344 18080
rect 4396 18068 4402 18080
rect 4433 18071 4491 18077
rect 4433 18068 4445 18071
rect 4396 18040 4445 18068
rect 4396 18028 4402 18040
rect 4433 18037 4445 18040
rect 4479 18037 4491 18071
rect 4433 18031 4491 18037
rect 4522 18028 4528 18080
rect 4580 18068 4586 18080
rect 5534 18068 5540 18080
rect 4580 18040 4625 18068
rect 5495 18040 5540 18068
rect 4580 18028 4586 18040
rect 5534 18028 5540 18040
rect 5592 18028 5598 18080
rect 5997 18071 6055 18077
rect 5997 18037 6009 18071
rect 6043 18068 6055 18071
rect 7834 18068 7840 18080
rect 6043 18040 7840 18068
rect 6043 18037 6055 18040
rect 5997 18031 6055 18037
rect 7834 18028 7840 18040
rect 7892 18028 7898 18080
rect 8220 18068 8248 18108
rect 8386 18096 8392 18108
rect 8444 18096 8450 18148
rect 9585 18139 9643 18145
rect 9585 18105 9597 18139
rect 9631 18136 9643 18139
rect 9950 18136 9956 18148
rect 9631 18108 9956 18136
rect 9631 18105 9643 18108
rect 9585 18099 9643 18105
rect 9950 18096 9956 18108
rect 10008 18096 10014 18148
rect 10060 18136 10088 18176
rect 10321 18173 10333 18207
rect 10367 18173 10379 18207
rect 11146 18204 11152 18216
rect 11107 18176 11152 18204
rect 10321 18167 10379 18173
rect 11146 18164 11152 18176
rect 11204 18164 11210 18216
rect 12434 18204 12440 18216
rect 12395 18176 12440 18204
rect 12434 18164 12440 18176
rect 12492 18164 12498 18216
rect 12621 18207 12679 18213
rect 12621 18173 12633 18207
rect 12667 18204 12679 18207
rect 17957 18207 18015 18213
rect 12667 18176 16574 18204
rect 12667 18173 12679 18176
rect 12621 18167 12679 18173
rect 11330 18136 11336 18148
rect 10060 18108 11336 18136
rect 11330 18096 11336 18108
rect 11388 18096 11394 18148
rect 11422 18096 11428 18148
rect 11480 18136 11486 18148
rect 11480 18108 11525 18136
rect 11480 18096 11486 18108
rect 8478 18068 8484 18080
rect 8220 18040 8484 18068
rect 8478 18028 8484 18040
rect 8536 18028 8542 18080
rect 10134 18028 10140 18080
rect 10192 18068 10198 18080
rect 10229 18071 10287 18077
rect 10229 18068 10241 18071
rect 10192 18040 10241 18068
rect 10192 18028 10198 18040
rect 10229 18037 10241 18040
rect 10275 18037 10287 18071
rect 10229 18031 10287 18037
rect 10689 18071 10747 18077
rect 10689 18037 10701 18071
rect 10735 18068 10747 18071
rect 11238 18068 11244 18080
rect 10735 18040 11244 18068
rect 10735 18037 10747 18040
rect 10689 18031 10747 18037
rect 11238 18028 11244 18040
rect 11296 18028 11302 18080
rect 12529 18071 12587 18077
rect 12529 18037 12541 18071
rect 12575 18068 12587 18071
rect 13446 18068 13452 18080
rect 12575 18040 13452 18068
rect 12575 18037 12587 18040
rect 12529 18031 12587 18037
rect 13446 18028 13452 18040
rect 13504 18028 13510 18080
rect 16546 18068 16574 18176
rect 17957 18173 17969 18207
rect 18003 18204 18015 18207
rect 18414 18204 18420 18216
rect 18003 18176 18420 18204
rect 18003 18173 18015 18176
rect 17957 18167 18015 18173
rect 18414 18164 18420 18176
rect 18472 18164 18478 18216
rect 17773 18071 17831 18077
rect 17773 18068 17785 18071
rect 16546 18040 17785 18068
rect 17773 18037 17785 18040
rect 17819 18037 17831 18071
rect 17773 18031 17831 18037
rect 184 17978 18920 18000
rect 184 17926 3106 17978
rect 3158 17926 3170 17978
rect 3222 17926 3234 17978
rect 3286 17926 3298 17978
rect 3350 17926 3362 17978
rect 3414 17926 6206 17978
rect 6258 17926 6270 17978
rect 6322 17926 6334 17978
rect 6386 17926 6398 17978
rect 6450 17926 6462 17978
rect 6514 17926 9306 17978
rect 9358 17926 9370 17978
rect 9422 17926 9434 17978
rect 9486 17926 9498 17978
rect 9550 17926 9562 17978
rect 9614 17926 12406 17978
rect 12458 17926 12470 17978
rect 12522 17926 12534 17978
rect 12586 17926 12598 17978
rect 12650 17926 12662 17978
rect 12714 17926 15506 17978
rect 15558 17926 15570 17978
rect 15622 17926 15634 17978
rect 15686 17926 15698 17978
rect 15750 17926 15762 17978
rect 15814 17926 18606 17978
rect 18658 17926 18670 17978
rect 18722 17926 18734 17978
rect 18786 17926 18798 17978
rect 18850 17926 18862 17978
rect 18914 17926 18920 17978
rect 184 17904 18920 17926
rect 3237 17867 3295 17873
rect 3237 17833 3249 17867
rect 3283 17864 3295 17867
rect 4522 17864 4528 17876
rect 3283 17836 4528 17864
rect 3283 17833 3295 17836
rect 3237 17827 3295 17833
rect 4522 17824 4528 17836
rect 4580 17824 4586 17876
rect 11747 17867 11805 17873
rect 11747 17833 11759 17867
rect 11793 17864 11805 17867
rect 12250 17864 12256 17876
rect 11793 17836 12256 17864
rect 11793 17833 11805 17836
rect 11747 17827 11805 17833
rect 12250 17824 12256 17836
rect 12308 17824 12314 17876
rect 13096 17836 15424 17864
rect 13096 17808 13124 17836
rect 937 17799 995 17805
rect 937 17765 949 17799
rect 983 17796 995 17799
rect 1210 17796 1216 17808
rect 983 17768 1216 17796
rect 983 17765 995 17768
rect 937 17759 995 17765
rect 1210 17756 1216 17768
rect 1268 17756 1274 17808
rect 2498 17796 2504 17808
rect 2162 17768 2504 17796
rect 2498 17756 2504 17768
rect 2556 17756 2562 17808
rect 4246 17756 4252 17808
rect 4304 17796 4310 17808
rect 5169 17799 5227 17805
rect 5169 17796 5181 17799
rect 4304 17768 5181 17796
rect 4304 17756 4310 17768
rect 5169 17765 5181 17768
rect 5215 17765 5227 17799
rect 7834 17796 7840 17808
rect 7795 17768 7840 17796
rect 5169 17759 5227 17765
rect 7834 17756 7840 17768
rect 7892 17756 7898 17808
rect 13078 17796 13084 17808
rect 11362 17768 13084 17796
rect 13078 17756 13084 17768
rect 13136 17756 13142 17808
rect 15396 17796 15424 17836
rect 15396 17768 15502 17796
rect 4525 17731 4583 17737
rect 4525 17697 4537 17731
rect 4571 17697 4583 17731
rect 9950 17728 9956 17740
rect 9911 17700 9956 17728
rect 4525 17691 4583 17697
rect 566 17620 572 17672
rect 624 17660 630 17672
rect 661 17663 719 17669
rect 661 17660 673 17663
rect 624 17632 673 17660
rect 624 17620 630 17632
rect 661 17629 673 17632
rect 707 17629 719 17663
rect 661 17623 719 17629
rect 4246 17620 4252 17672
rect 4304 17660 4310 17672
rect 4540 17660 4568 17691
rect 9950 17688 9956 17700
rect 10008 17688 10014 17740
rect 12250 17688 12256 17740
rect 12308 17728 12314 17740
rect 12345 17731 12403 17737
rect 12345 17728 12357 17731
rect 12308 17700 12357 17728
rect 12308 17688 12314 17700
rect 12345 17697 12357 17700
rect 12391 17697 12403 17731
rect 17494 17728 17500 17740
rect 17455 17700 17500 17728
rect 12345 17691 12403 17697
rect 17494 17688 17500 17700
rect 17552 17688 17558 17740
rect 10318 17660 10324 17672
rect 4304 17632 6500 17660
rect 10279 17632 10324 17660
rect 4304 17620 4310 17632
rect 6472 17601 6500 17632
rect 10318 17620 10324 17632
rect 10376 17620 10382 17672
rect 13814 17620 13820 17672
rect 13872 17660 13878 17672
rect 14734 17660 14740 17672
rect 13872 17632 14740 17660
rect 13872 17620 13878 17632
rect 14734 17620 14740 17632
rect 14792 17620 14798 17672
rect 15102 17660 15108 17672
rect 15063 17632 15108 17660
rect 15102 17620 15108 17632
rect 15160 17620 15166 17672
rect 16577 17663 16635 17669
rect 16577 17629 16589 17663
rect 16623 17660 16635 17663
rect 16942 17660 16948 17672
rect 16623 17632 16948 17660
rect 16623 17629 16635 17632
rect 16577 17623 16635 17629
rect 16942 17620 16948 17632
rect 17000 17620 17006 17672
rect 17589 17663 17647 17669
rect 17589 17629 17601 17663
rect 17635 17660 17647 17663
rect 17678 17660 17684 17672
rect 17635 17632 17684 17660
rect 17635 17629 17647 17632
rect 17589 17623 17647 17629
rect 17678 17620 17684 17632
rect 17736 17620 17742 17672
rect 17773 17663 17831 17669
rect 17773 17629 17785 17663
rect 17819 17660 17831 17663
rect 17862 17660 17868 17672
rect 17819 17632 17868 17660
rect 17819 17629 17831 17632
rect 17773 17623 17831 17629
rect 17862 17620 17868 17632
rect 17920 17620 17926 17672
rect 6457 17595 6515 17601
rect 6457 17561 6469 17595
rect 6503 17561 6515 17595
rect 14274 17592 14280 17604
rect 6457 17555 6515 17561
rect 11072 17564 14280 17592
rect 2406 17524 2412 17536
rect 2367 17496 2412 17524
rect 2406 17484 2412 17496
rect 2464 17484 2470 17536
rect 7006 17484 7012 17536
rect 7064 17524 7070 17536
rect 9309 17527 9367 17533
rect 9309 17524 9321 17527
rect 7064 17496 9321 17524
rect 7064 17484 7070 17496
rect 9309 17493 9321 17496
rect 9355 17524 9367 17527
rect 11072 17524 11100 17564
rect 14274 17552 14280 17564
rect 14332 17552 14338 17604
rect 9355 17496 11100 17524
rect 9355 17493 9367 17496
rect 9309 17487 9367 17493
rect 11974 17484 11980 17536
rect 12032 17524 12038 17536
rect 13633 17527 13691 17533
rect 13633 17524 13645 17527
rect 12032 17496 13645 17524
rect 12032 17484 12038 17496
rect 13633 17493 13645 17496
rect 13679 17493 13691 17527
rect 13633 17487 13691 17493
rect 16850 17484 16856 17536
rect 16908 17524 16914 17536
rect 17129 17527 17187 17533
rect 17129 17524 17141 17527
rect 16908 17496 17141 17524
rect 16908 17484 16914 17496
rect 17129 17493 17141 17496
rect 17175 17493 17187 17527
rect 17129 17487 17187 17493
rect 184 17434 18860 17456
rect 184 17382 1556 17434
rect 1608 17382 1620 17434
rect 1672 17382 1684 17434
rect 1736 17382 1748 17434
rect 1800 17382 1812 17434
rect 1864 17382 4656 17434
rect 4708 17382 4720 17434
rect 4772 17382 4784 17434
rect 4836 17382 4848 17434
rect 4900 17382 4912 17434
rect 4964 17382 7756 17434
rect 7808 17382 7820 17434
rect 7872 17382 7884 17434
rect 7936 17382 7948 17434
rect 8000 17382 8012 17434
rect 8064 17382 10856 17434
rect 10908 17382 10920 17434
rect 10972 17382 10984 17434
rect 11036 17382 11048 17434
rect 11100 17382 11112 17434
rect 11164 17382 13956 17434
rect 14008 17382 14020 17434
rect 14072 17382 14084 17434
rect 14136 17382 14148 17434
rect 14200 17382 14212 17434
rect 14264 17382 17056 17434
rect 17108 17382 17120 17434
rect 17172 17382 17184 17434
rect 17236 17382 17248 17434
rect 17300 17382 17312 17434
rect 17364 17382 18860 17434
rect 184 17360 18860 17382
rect 1673 17323 1731 17329
rect 1673 17289 1685 17323
rect 1719 17320 1731 17323
rect 1946 17320 1952 17332
rect 1719 17292 1952 17320
rect 1719 17289 1731 17292
rect 1673 17283 1731 17289
rect 1946 17280 1952 17292
rect 2004 17280 2010 17332
rect 3605 17323 3663 17329
rect 3605 17289 3617 17323
rect 3651 17320 3663 17323
rect 4154 17320 4160 17332
rect 3651 17292 4160 17320
rect 3651 17289 3663 17292
rect 3605 17283 3663 17289
rect 4154 17280 4160 17292
rect 4212 17280 4218 17332
rect 5534 17280 5540 17332
rect 5592 17320 5598 17332
rect 5813 17323 5871 17329
rect 5813 17320 5825 17323
rect 5592 17292 5825 17320
rect 5592 17280 5598 17292
rect 5813 17289 5825 17292
rect 5859 17289 5871 17323
rect 5813 17283 5871 17289
rect 10042 17280 10048 17332
rect 10100 17320 10106 17332
rect 12437 17323 12495 17329
rect 12437 17320 12449 17323
rect 10100 17292 12449 17320
rect 10100 17280 10106 17292
rect 12437 17289 12449 17292
rect 12483 17289 12495 17323
rect 12437 17283 12495 17289
rect 14200 17292 17632 17320
rect 10318 17212 10324 17264
rect 10376 17252 10382 17264
rect 10551 17255 10609 17261
rect 10551 17252 10563 17255
rect 10376 17224 10563 17252
rect 10376 17212 10382 17224
rect 10551 17221 10563 17224
rect 10597 17221 10609 17255
rect 10551 17215 10609 17221
rect 2498 17184 2504 17196
rect 2459 17156 2504 17184
rect 2498 17144 2504 17156
rect 2556 17144 2562 17196
rect 4338 17184 4344 17196
rect 4299 17156 4344 17184
rect 4338 17144 4344 17156
rect 4396 17144 4402 17196
rect 6546 17184 6552 17196
rect 6507 17156 6552 17184
rect 6546 17144 6552 17156
rect 6604 17144 6610 17196
rect 6917 17187 6975 17193
rect 6917 17153 6929 17187
rect 6963 17184 6975 17187
rect 7282 17184 7288 17196
rect 6963 17156 7288 17184
rect 6963 17153 6975 17156
rect 6917 17147 6975 17153
rect 7282 17144 7288 17156
rect 7340 17144 7346 17196
rect 8386 17144 8392 17196
rect 8444 17184 8450 17196
rect 8757 17187 8815 17193
rect 8757 17184 8769 17187
rect 8444 17156 8769 17184
rect 8444 17144 8450 17156
rect 8757 17153 8769 17156
rect 8803 17153 8815 17187
rect 8757 17147 8815 17153
rect 1578 17116 1584 17128
rect 1539 17088 1584 17116
rect 1578 17076 1584 17088
rect 1636 17076 1642 17128
rect 1762 17116 1768 17128
rect 1723 17088 1768 17116
rect 1762 17076 1768 17088
rect 1820 17076 1826 17128
rect 1854 17076 1860 17128
rect 1912 17125 1918 17128
rect 1912 17119 1961 17125
rect 1912 17085 1915 17119
rect 1949 17085 1961 17119
rect 1912 17079 1961 17085
rect 2041 17119 2099 17125
rect 2041 17085 2053 17119
rect 2087 17116 2099 17119
rect 2222 17116 2228 17128
rect 2087 17088 2228 17116
rect 2087 17085 2099 17088
rect 2041 17079 2099 17085
rect 1912 17076 1918 17079
rect 2222 17076 2228 17088
rect 2280 17076 2286 17128
rect 2314 17076 2320 17128
rect 2372 17116 2378 17128
rect 2958 17116 2964 17128
rect 2372 17088 2964 17116
rect 2372 17076 2378 17088
rect 2958 17076 2964 17088
rect 3016 17076 3022 17128
rect 3510 17076 3516 17128
rect 3568 17116 3574 17128
rect 4065 17119 4123 17125
rect 4065 17116 4077 17119
rect 3568 17088 4077 17116
rect 3568 17076 3574 17088
rect 4065 17085 4077 17088
rect 4111 17085 4123 17119
rect 9125 17119 9183 17125
rect 9125 17116 9137 17119
rect 4065 17079 4123 17085
rect 8772 17088 9137 17116
rect 2498 17008 2504 17060
rect 2556 17048 2562 17060
rect 4430 17048 4436 17060
rect 2556 17020 4436 17048
rect 2556 17008 2562 17020
rect 4430 17008 4436 17020
rect 4488 17048 4494 17060
rect 8343 17051 8401 17057
rect 4488 17020 4830 17048
rect 7208 17020 7314 17048
rect 4488 17008 4494 17020
rect 4724 16980 4752 17020
rect 6822 16980 6828 16992
rect 4724 16952 6828 16980
rect 6822 16940 6828 16952
rect 6880 16980 6886 16992
rect 7208 16980 7236 17020
rect 8343 17017 8355 17051
rect 8389 17048 8401 17051
rect 8772 17048 8800 17088
rect 9125 17085 9137 17088
rect 9171 17085 9183 17119
rect 9125 17079 9183 17085
rect 11149 17119 11207 17125
rect 11149 17085 11161 17119
rect 11195 17116 11207 17119
rect 11238 17116 11244 17128
rect 11195 17088 11244 17116
rect 11195 17085 11207 17088
rect 11149 17079 11207 17085
rect 11238 17076 11244 17088
rect 11296 17076 11302 17128
rect 8389 17020 8800 17048
rect 9416 17020 9522 17048
rect 8389 17017 8401 17020
rect 8343 17011 8401 17017
rect 9416 16980 9444 17020
rect 13078 17008 13084 17060
rect 13136 17048 13142 17060
rect 14200 17048 14228 17292
rect 14734 17144 14740 17196
rect 14792 17184 14798 17196
rect 15565 17187 15623 17193
rect 15565 17184 15577 17187
rect 14792 17156 15577 17184
rect 14792 17144 14798 17156
rect 15565 17153 15577 17156
rect 15611 17184 15623 17187
rect 16209 17187 16267 17193
rect 16209 17184 16221 17187
rect 15611 17156 16221 17184
rect 15611 17153 15623 17156
rect 15565 17147 15623 17153
rect 16209 17153 16221 17156
rect 16255 17153 16267 17187
rect 16209 17147 16267 17153
rect 16485 17187 16543 17193
rect 16485 17153 16497 17187
rect 16531 17184 16543 17187
rect 16850 17184 16856 17196
rect 16531 17156 16856 17184
rect 16531 17153 16543 17156
rect 16485 17147 16543 17153
rect 16850 17144 16856 17156
rect 16908 17144 16914 17196
rect 15197 17119 15255 17125
rect 15197 17085 15209 17119
rect 15243 17116 15255 17119
rect 15243 17088 15884 17116
rect 17604 17102 17632 17292
rect 17678 17280 17684 17332
rect 17736 17320 17742 17332
rect 17957 17323 18015 17329
rect 17957 17320 17969 17323
rect 17736 17292 17969 17320
rect 17736 17280 17742 17292
rect 17957 17289 17969 17292
rect 18003 17289 18015 17323
rect 17957 17283 18015 17289
rect 15243 17085 15255 17088
rect 15197 17079 15255 17085
rect 13136 17034 14228 17048
rect 15856 17048 15884 17088
rect 16574 17048 16580 17060
rect 13136 17020 14214 17034
rect 15856 17020 16580 17048
rect 13136 17008 13142 17020
rect 16574 17008 16580 17020
rect 16632 17008 16638 17060
rect 6880 16952 9444 16980
rect 13771 16983 13829 16989
rect 6880 16940 6886 16952
rect 13771 16949 13783 16983
rect 13817 16980 13829 16983
rect 15930 16980 15936 16992
rect 13817 16952 15936 16980
rect 13817 16949 13829 16952
rect 13771 16943 13829 16949
rect 15930 16940 15936 16952
rect 15988 16940 15994 16992
rect 184 16890 18920 16912
rect 184 16838 3106 16890
rect 3158 16838 3170 16890
rect 3222 16838 3234 16890
rect 3286 16838 3298 16890
rect 3350 16838 3362 16890
rect 3414 16838 6206 16890
rect 6258 16838 6270 16890
rect 6322 16838 6334 16890
rect 6386 16838 6398 16890
rect 6450 16838 6462 16890
rect 6514 16838 9306 16890
rect 9358 16838 9370 16890
rect 9422 16838 9434 16890
rect 9486 16838 9498 16890
rect 9550 16838 9562 16890
rect 9614 16838 12406 16890
rect 12458 16838 12470 16890
rect 12522 16838 12534 16890
rect 12586 16838 12598 16890
rect 12650 16838 12662 16890
rect 12714 16838 15506 16890
rect 15558 16838 15570 16890
rect 15622 16838 15634 16890
rect 15686 16838 15698 16890
rect 15750 16838 15762 16890
rect 15814 16838 18606 16890
rect 18658 16838 18670 16890
rect 18722 16838 18734 16890
rect 18786 16838 18798 16890
rect 18850 16838 18862 16890
rect 18914 16838 18920 16890
rect 184 16816 18920 16838
rect 1670 16776 1676 16788
rect 1631 16748 1676 16776
rect 1670 16736 1676 16748
rect 1728 16736 1734 16788
rect 2406 16776 2412 16788
rect 1780 16748 2412 16776
rect 1578 16708 1584 16720
rect 1491 16680 1584 16708
rect 1578 16668 1584 16680
rect 1636 16708 1642 16720
rect 1780 16708 1808 16748
rect 2406 16736 2412 16748
rect 2464 16776 2470 16788
rect 2464 16748 3188 16776
rect 2464 16736 2470 16748
rect 1636 16680 1808 16708
rect 1636 16668 1642 16680
rect 1854 16640 1860 16652
rect 1767 16612 1860 16640
rect 1854 16600 1860 16612
rect 1912 16640 1918 16652
rect 3160 16649 3188 16748
rect 4338 16736 4344 16788
rect 4396 16776 4402 16788
rect 4801 16779 4859 16785
rect 4801 16776 4813 16779
rect 4396 16748 4813 16776
rect 4396 16736 4402 16748
rect 4801 16745 4813 16748
rect 4847 16745 4859 16779
rect 4801 16739 4859 16745
rect 12158 16736 12164 16788
rect 12216 16776 12222 16788
rect 16022 16776 16028 16788
rect 12216 16748 14136 16776
rect 15983 16748 16028 16776
rect 12216 16736 12222 16748
rect 3688 16711 3746 16717
rect 3688 16677 3700 16711
rect 3734 16708 3746 16711
rect 4062 16708 4068 16720
rect 3734 16680 4068 16708
rect 3734 16677 3746 16680
rect 3688 16671 3746 16677
rect 4062 16668 4068 16680
rect 4120 16668 4126 16720
rect 7006 16708 7012 16720
rect 6967 16680 7012 16708
rect 7006 16668 7012 16680
rect 7064 16668 7070 16720
rect 9585 16711 9643 16717
rect 9585 16677 9597 16711
rect 9631 16708 9643 16711
rect 10226 16708 10232 16720
rect 9631 16680 10232 16708
rect 9631 16677 9643 16680
rect 9585 16671 9643 16677
rect 10226 16668 10232 16680
rect 10284 16668 10290 16720
rect 12526 16708 12532 16720
rect 11730 16680 12532 16708
rect 12526 16668 12532 16680
rect 12584 16668 12590 16720
rect 13078 16668 13084 16720
rect 13136 16668 13142 16720
rect 2961 16643 3019 16649
rect 2961 16640 2973 16643
rect 1912 16612 2973 16640
rect 1912 16600 1918 16612
rect 2961 16609 2973 16612
rect 3007 16609 3019 16643
rect 2961 16603 3019 16609
rect 3145 16643 3203 16649
rect 3145 16609 3157 16643
rect 3191 16609 3203 16643
rect 3145 16603 3203 16609
rect 3421 16643 3479 16649
rect 3421 16609 3433 16643
rect 3467 16640 3479 16643
rect 3510 16640 3516 16652
rect 3467 16612 3516 16640
rect 3467 16609 3479 16612
rect 3421 16603 3479 16609
rect 1762 16572 1768 16584
rect 1723 16544 1768 16572
rect 1762 16532 1768 16544
rect 1820 16532 1826 16584
rect 1949 16575 2007 16581
rect 1949 16541 1961 16575
rect 1995 16572 2007 16575
rect 2222 16572 2228 16584
rect 1995 16544 2228 16572
rect 1995 16541 2007 16544
rect 1949 16535 2007 16541
rect 2222 16532 2228 16544
rect 2280 16532 2286 16584
rect 566 16464 572 16516
rect 624 16504 630 16516
rect 3436 16504 3464 16603
rect 3510 16600 3516 16612
rect 3568 16600 3574 16652
rect 14108 16649 14136 16748
rect 16022 16736 16028 16748
rect 16080 16736 16086 16788
rect 17221 16779 17279 16785
rect 17221 16745 17233 16779
rect 17267 16776 17279 16779
rect 17494 16776 17500 16788
rect 17267 16748 17500 16776
rect 17267 16745 17279 16748
rect 17221 16739 17279 16745
rect 17494 16736 17500 16748
rect 17552 16736 17558 16788
rect 14274 16668 14280 16720
rect 14332 16708 14338 16720
rect 14737 16711 14795 16717
rect 14737 16708 14749 16711
rect 14332 16680 14749 16708
rect 14332 16668 14338 16680
rect 14737 16677 14749 16680
rect 14783 16677 14795 16711
rect 14737 16671 14795 16677
rect 14093 16643 14151 16649
rect 14093 16609 14105 16643
rect 14139 16609 14151 16643
rect 14093 16603 14151 16609
rect 17494 16600 17500 16652
rect 17552 16640 17558 16652
rect 17589 16643 17647 16649
rect 17589 16640 17601 16643
rect 17552 16612 17601 16640
rect 17552 16600 17558 16612
rect 17589 16609 17601 16612
rect 17635 16609 17647 16643
rect 18414 16640 18420 16652
rect 18375 16612 18420 16640
rect 17589 16603 17647 16609
rect 18414 16600 18420 16612
rect 18472 16600 18478 16652
rect 7650 16532 7656 16584
rect 7708 16572 7714 16584
rect 7837 16575 7895 16581
rect 7837 16572 7849 16575
rect 7708 16544 7849 16572
rect 7708 16532 7714 16544
rect 7837 16541 7849 16544
rect 7883 16541 7895 16575
rect 7837 16535 7895 16541
rect 10134 16532 10140 16584
rect 10192 16572 10198 16584
rect 10229 16575 10287 16581
rect 10229 16572 10241 16575
rect 10192 16544 10241 16572
rect 10192 16532 10198 16544
rect 10229 16541 10241 16544
rect 10275 16541 10287 16575
rect 10229 16535 10287 16541
rect 10505 16575 10563 16581
rect 10505 16541 10517 16575
rect 10551 16572 10563 16575
rect 13817 16575 13875 16581
rect 10551 16544 12848 16572
rect 10551 16541 10563 16544
rect 10505 16535 10563 16541
rect 624 16476 3464 16504
rect 624 16464 630 16476
rect 1762 16396 1768 16448
rect 1820 16436 1826 16448
rect 2038 16436 2044 16448
rect 1820 16408 2044 16436
rect 1820 16396 1826 16408
rect 2038 16396 2044 16408
rect 2096 16436 2102 16448
rect 2774 16436 2780 16448
rect 2096 16408 2780 16436
rect 2096 16396 2102 16408
rect 2774 16396 2780 16408
rect 2832 16396 2838 16448
rect 3145 16439 3203 16445
rect 3145 16405 3157 16439
rect 3191 16436 3203 16439
rect 3418 16436 3424 16448
rect 3191 16408 3424 16436
rect 3191 16405 3203 16408
rect 3145 16399 3203 16405
rect 3418 16396 3424 16408
rect 3476 16396 3482 16448
rect 5721 16439 5779 16445
rect 5721 16405 5733 16439
rect 5767 16436 5779 16439
rect 7466 16436 7472 16448
rect 5767 16408 7472 16436
rect 5767 16405 5779 16408
rect 5721 16399 5779 16405
rect 7466 16396 7472 16408
rect 7524 16396 7530 16448
rect 11977 16439 12035 16445
rect 11977 16405 11989 16439
rect 12023 16436 12035 16439
rect 12066 16436 12072 16448
rect 12023 16408 12072 16436
rect 12023 16405 12035 16408
rect 11977 16399 12035 16405
rect 12066 16396 12072 16408
rect 12124 16396 12130 16448
rect 12345 16439 12403 16445
rect 12345 16405 12357 16439
rect 12391 16436 12403 16439
rect 12710 16436 12716 16448
rect 12391 16408 12716 16436
rect 12391 16405 12403 16408
rect 12345 16399 12403 16405
rect 12710 16396 12716 16408
rect 12768 16396 12774 16448
rect 12820 16436 12848 16544
rect 13817 16541 13829 16575
rect 13863 16572 13875 16575
rect 17678 16572 17684 16584
rect 13863 16544 16574 16572
rect 17639 16544 17684 16572
rect 13863 16541 13875 16544
rect 13817 16535 13875 16541
rect 16546 16504 16574 16544
rect 17678 16532 17684 16544
rect 17736 16532 17742 16584
rect 17770 16532 17776 16584
rect 17828 16572 17834 16584
rect 17828 16544 17873 16572
rect 17828 16532 17834 16544
rect 18046 16504 18052 16516
rect 16546 16476 18052 16504
rect 18046 16464 18052 16476
rect 18104 16464 18110 16516
rect 18233 16439 18291 16445
rect 18233 16436 18245 16439
rect 12820 16408 18245 16436
rect 18233 16405 18245 16408
rect 18279 16405 18291 16439
rect 18233 16399 18291 16405
rect 184 16346 18860 16368
rect 184 16294 1556 16346
rect 1608 16294 1620 16346
rect 1672 16294 1684 16346
rect 1736 16294 1748 16346
rect 1800 16294 1812 16346
rect 1864 16294 4656 16346
rect 4708 16294 4720 16346
rect 4772 16294 4784 16346
rect 4836 16294 4848 16346
rect 4900 16294 4912 16346
rect 4964 16294 7756 16346
rect 7808 16294 7820 16346
rect 7872 16294 7884 16346
rect 7936 16294 7948 16346
rect 8000 16294 8012 16346
rect 8064 16294 10856 16346
rect 10908 16294 10920 16346
rect 10972 16294 10984 16346
rect 11036 16294 11048 16346
rect 11100 16294 11112 16346
rect 11164 16294 13956 16346
rect 14008 16294 14020 16346
rect 14072 16294 14084 16346
rect 14136 16294 14148 16346
rect 14200 16294 14212 16346
rect 14264 16294 17056 16346
rect 17108 16294 17120 16346
rect 17172 16294 17184 16346
rect 17236 16294 17248 16346
rect 17300 16294 17312 16346
rect 17364 16294 18860 16346
rect 184 16272 18860 16294
rect 5442 16192 5448 16244
rect 5500 16232 5506 16244
rect 5537 16235 5595 16241
rect 5537 16232 5549 16235
rect 5500 16204 5549 16232
rect 5500 16192 5506 16204
rect 5537 16201 5549 16204
rect 5583 16201 5595 16235
rect 5537 16195 5595 16201
rect 6825 16235 6883 16241
rect 6825 16201 6837 16235
rect 6871 16232 6883 16235
rect 7098 16232 7104 16244
rect 6871 16204 7104 16232
rect 6871 16201 6883 16204
rect 6825 16195 6883 16201
rect 7098 16192 7104 16204
rect 7156 16192 7162 16244
rect 11330 16192 11336 16244
rect 11388 16232 11394 16244
rect 12437 16235 12495 16241
rect 12437 16232 12449 16235
rect 11388 16204 12449 16232
rect 11388 16192 11394 16204
rect 12437 16201 12449 16204
rect 12483 16201 12495 16235
rect 12437 16195 12495 16201
rect 16114 16192 16120 16244
rect 16172 16232 16178 16244
rect 17770 16232 17776 16244
rect 16172 16204 17776 16232
rect 16172 16192 16178 16204
rect 17770 16192 17776 16204
rect 17828 16192 17834 16244
rect 18414 16232 18420 16244
rect 18375 16204 18420 16232
rect 18414 16192 18420 16204
rect 18472 16192 18478 16244
rect 17678 16164 17684 16176
rect 17639 16136 17684 16164
rect 17678 16124 17684 16136
rect 17736 16124 17742 16176
rect 1946 16056 1952 16108
rect 2004 16096 2010 16108
rect 2041 16099 2099 16105
rect 2041 16096 2053 16099
rect 2004 16068 2053 16096
rect 2004 16056 2010 16068
rect 2041 16065 2053 16068
rect 2087 16065 2099 16099
rect 2222 16096 2228 16108
rect 2183 16068 2228 16096
rect 2041 16059 2099 16065
rect 2056 16028 2084 16059
rect 2222 16056 2228 16068
rect 2280 16056 2286 16108
rect 2774 16096 2780 16108
rect 2735 16068 2780 16096
rect 2774 16056 2780 16068
rect 2832 16056 2838 16108
rect 12066 16056 12072 16108
rect 12124 16096 12130 16108
rect 13817 16099 13875 16105
rect 13817 16096 13829 16099
rect 12124 16068 13829 16096
rect 12124 16056 12130 16068
rect 13817 16065 13829 16068
rect 13863 16065 13875 16099
rect 13817 16059 13875 16065
rect 15933 16099 15991 16105
rect 15933 16065 15945 16099
rect 15979 16096 15991 16099
rect 16022 16096 16028 16108
rect 15979 16068 16028 16096
rect 15979 16065 15991 16068
rect 15933 16059 15991 16065
rect 16022 16056 16028 16068
rect 16080 16056 16086 16108
rect 16942 16056 16948 16108
rect 17000 16096 17006 16108
rect 17221 16099 17279 16105
rect 17221 16096 17233 16099
rect 17000 16068 17233 16096
rect 17000 16056 17006 16068
rect 17221 16065 17233 16068
rect 17267 16065 17279 16099
rect 17221 16059 17279 16065
rect 2869 16031 2927 16037
rect 2869 16028 2881 16031
rect 2056 16000 2881 16028
rect 2869 15997 2881 16000
rect 2915 15997 2927 16031
rect 4246 16028 4252 16040
rect 4207 16000 4252 16028
rect 2869 15991 2927 15997
rect 4246 15988 4252 16000
rect 4304 15988 4310 16040
rect 10134 15988 10140 16040
rect 10192 16028 10198 16040
rect 13541 16031 13599 16037
rect 13541 16028 13553 16031
rect 10192 16000 13553 16028
rect 10192 15988 10198 16000
rect 13541 15997 13553 16000
rect 13587 15997 13599 16031
rect 16114 16028 16120 16040
rect 16075 16000 16120 16028
rect 13541 15991 13599 15997
rect 16114 15988 16120 16000
rect 16172 15988 16178 16040
rect 16209 16031 16267 16037
rect 16209 15997 16221 16031
rect 16255 16028 16267 16031
rect 17313 16031 17371 16037
rect 16255 16000 16804 16028
rect 16255 15997 16267 16000
rect 16209 15991 16267 15997
rect 1949 15963 2007 15969
rect 1949 15929 1961 15963
rect 1995 15960 2007 15963
rect 2958 15960 2964 15972
rect 1995 15932 2964 15960
rect 1995 15929 2007 15932
rect 1949 15923 2007 15929
rect 2958 15920 2964 15932
rect 3016 15920 3022 15972
rect 8113 15963 8171 15969
rect 8113 15929 8125 15963
rect 8159 15929 8171 15963
rect 8754 15960 8760 15972
rect 8715 15932 8760 15960
rect 8113 15923 8171 15929
rect 842 15852 848 15904
rect 900 15892 906 15904
rect 1581 15895 1639 15901
rect 1581 15892 1593 15895
rect 900 15864 1593 15892
rect 900 15852 906 15864
rect 1581 15861 1593 15864
rect 1627 15861 1639 15895
rect 1581 15855 1639 15861
rect 3237 15895 3295 15901
rect 3237 15861 3249 15895
rect 3283 15892 3295 15895
rect 3694 15892 3700 15904
rect 3283 15864 3700 15892
rect 3283 15861 3295 15864
rect 3237 15855 3295 15861
rect 3694 15852 3700 15864
rect 3752 15852 3758 15904
rect 8128 15892 8156 15923
rect 8754 15920 8760 15932
rect 8812 15920 8818 15972
rect 11149 15963 11207 15969
rect 11149 15929 11161 15963
rect 11195 15929 11207 15963
rect 11149 15923 11207 15929
rect 10045 15895 10103 15901
rect 10045 15892 10057 15895
rect 8128 15864 10057 15892
rect 10045 15861 10057 15864
rect 10091 15892 10103 15895
rect 11164 15892 11192 15923
rect 12526 15920 12532 15972
rect 12584 15960 12590 15972
rect 13078 15960 13084 15972
rect 12584 15932 13084 15960
rect 12584 15920 12590 15932
rect 13078 15920 13084 15932
rect 13136 15960 13142 15972
rect 13136 15932 14306 15960
rect 13136 15920 13142 15932
rect 15194 15920 15200 15972
rect 15252 15960 15258 15972
rect 16224 15960 16252 15991
rect 15252 15932 16252 15960
rect 15252 15920 15258 15932
rect 16298 15920 16304 15972
rect 16356 15960 16362 15972
rect 16776 15969 16804 16000
rect 17313 15997 17325 16031
rect 17359 16028 17371 16031
rect 17586 16028 17592 16040
rect 17359 16000 17592 16028
rect 17359 15997 17371 16000
rect 17313 15991 17371 15997
rect 17586 15988 17592 16000
rect 17644 15988 17650 16040
rect 16577 15963 16635 15969
rect 16577 15960 16589 15963
rect 16356 15932 16589 15960
rect 16356 15920 16362 15932
rect 16577 15929 16589 15932
rect 16623 15929 16635 15963
rect 16577 15923 16635 15929
rect 16761 15963 16819 15969
rect 16761 15929 16773 15963
rect 16807 15960 16819 15963
rect 17862 15960 17868 15972
rect 16807 15932 17868 15960
rect 16807 15929 16819 15932
rect 16761 15923 16819 15929
rect 17862 15920 17868 15932
rect 17920 15920 17926 15972
rect 15286 15892 15292 15904
rect 10091 15864 11192 15892
rect 15247 15864 15292 15892
rect 10091 15861 10103 15864
rect 10045 15855 10103 15861
rect 15286 15852 15292 15864
rect 15344 15852 15350 15904
rect 15930 15892 15936 15904
rect 15891 15864 15936 15892
rect 15930 15852 15936 15864
rect 15988 15852 15994 15904
rect 184 15802 18920 15824
rect 184 15750 3106 15802
rect 3158 15750 3170 15802
rect 3222 15750 3234 15802
rect 3286 15750 3298 15802
rect 3350 15750 3362 15802
rect 3414 15750 6206 15802
rect 6258 15750 6270 15802
rect 6322 15750 6334 15802
rect 6386 15750 6398 15802
rect 6450 15750 6462 15802
rect 6514 15750 9306 15802
rect 9358 15750 9370 15802
rect 9422 15750 9434 15802
rect 9486 15750 9498 15802
rect 9550 15750 9562 15802
rect 9614 15750 12406 15802
rect 12458 15750 12470 15802
rect 12522 15750 12534 15802
rect 12586 15750 12598 15802
rect 12650 15750 12662 15802
rect 12714 15750 15506 15802
rect 15558 15750 15570 15802
rect 15622 15750 15634 15802
rect 15686 15750 15698 15802
rect 15750 15750 15762 15802
rect 15814 15750 18606 15802
rect 18658 15750 18670 15802
rect 18722 15750 18734 15802
rect 18786 15750 18798 15802
rect 18850 15750 18862 15802
rect 18914 15750 18920 15802
rect 184 15728 18920 15750
rect 7193 15691 7251 15697
rect 6840 15660 7052 15688
rect 842 15620 848 15632
rect 803 15592 848 15620
rect 842 15580 848 15592
rect 900 15580 906 15632
rect 2130 15620 2136 15632
rect 2043 15592 2136 15620
rect 2130 15580 2136 15592
rect 2188 15620 2194 15632
rect 2498 15620 2504 15632
rect 2188 15592 2504 15620
rect 2188 15580 2194 15592
rect 2498 15580 2504 15592
rect 2556 15580 2562 15632
rect 4154 15580 4160 15632
rect 4212 15620 4218 15632
rect 4525 15623 4583 15629
rect 4525 15620 4537 15623
rect 4212 15592 4537 15620
rect 4212 15580 4218 15592
rect 4525 15589 4537 15592
rect 4571 15620 4583 15623
rect 5810 15620 5816 15632
rect 4571 15592 5816 15620
rect 4571 15589 4583 15592
rect 4525 15583 4583 15589
rect 5810 15580 5816 15592
rect 5868 15580 5874 15632
rect 6840 15564 6868 15660
rect 7024 15620 7052 15660
rect 7193 15657 7205 15691
rect 7239 15688 7251 15691
rect 7558 15688 7564 15700
rect 7239 15660 7564 15688
rect 7239 15657 7251 15660
rect 7193 15651 7251 15657
rect 7558 15648 7564 15660
rect 7616 15688 7622 15700
rect 9674 15688 9680 15700
rect 7616 15660 9680 15688
rect 7616 15648 7622 15660
rect 9674 15648 9680 15660
rect 9732 15648 9738 15700
rect 12802 15648 12808 15700
rect 12860 15648 12866 15700
rect 12894 15648 12900 15700
rect 12952 15688 12958 15700
rect 14274 15688 14280 15700
rect 12952 15660 14280 15688
rect 12952 15648 12958 15660
rect 14274 15648 14280 15660
rect 14332 15648 14338 15700
rect 14737 15691 14795 15697
rect 14737 15657 14749 15691
rect 14783 15688 14795 15691
rect 15102 15688 15108 15700
rect 14783 15660 15108 15688
rect 14783 15657 14795 15660
rect 14737 15651 14795 15657
rect 15102 15648 15108 15660
rect 15160 15648 15166 15700
rect 16298 15688 16304 15700
rect 15304 15660 16304 15688
rect 7024 15592 8602 15620
rect 10134 15580 10140 15632
rect 10192 15620 10198 15632
rect 10229 15623 10287 15629
rect 10229 15620 10241 15623
rect 10192 15592 10241 15620
rect 10192 15580 10198 15592
rect 10229 15589 10241 15592
rect 10275 15589 10287 15623
rect 11974 15620 11980 15632
rect 11935 15592 11980 15620
rect 10229 15583 10287 15589
rect 11974 15580 11980 15592
rect 12032 15580 12038 15632
rect 12621 15623 12679 15629
rect 12621 15589 12633 15623
rect 12667 15620 12679 15623
rect 12820 15620 12848 15648
rect 12667 15592 12848 15620
rect 12667 15589 12679 15592
rect 12621 15583 12679 15589
rect 13078 15580 13084 15632
rect 13136 15580 13142 15632
rect 15304 15620 15332 15660
rect 16298 15648 16304 15660
rect 16356 15648 16362 15700
rect 16574 15648 16580 15700
rect 16632 15688 16638 15700
rect 17221 15691 17279 15697
rect 16632 15660 16677 15688
rect 16632 15648 16638 15660
rect 17221 15657 17233 15691
rect 17267 15688 17279 15691
rect 17770 15688 17776 15700
rect 17267 15660 17776 15688
rect 17267 15657 17279 15660
rect 17221 15651 17279 15657
rect 17770 15648 17776 15660
rect 17828 15648 17834 15700
rect 14108 15592 15332 15620
rect 566 15552 572 15564
rect 527 15524 572 15552
rect 566 15512 572 15524
rect 624 15512 630 15564
rect 4801 15555 4859 15561
rect 4801 15521 4813 15555
rect 4847 15521 4859 15555
rect 4801 15515 4859 15521
rect 1946 15376 1952 15428
rect 2004 15416 2010 15428
rect 2317 15419 2375 15425
rect 2317 15416 2329 15419
rect 2004 15388 2329 15416
rect 2004 15376 2010 15388
rect 2317 15385 2329 15388
rect 2363 15385 2375 15419
rect 2317 15379 2375 15385
rect 4816 15348 4844 15515
rect 6822 15512 6828 15564
rect 6880 15512 6886 15564
rect 5442 15484 5448 15496
rect 5403 15456 5448 15484
rect 5442 15444 5448 15456
rect 5500 15444 5506 15496
rect 5718 15484 5724 15496
rect 5631 15456 5724 15484
rect 5718 15444 5724 15456
rect 5776 15484 5782 15496
rect 7282 15484 7288 15496
rect 5776 15456 7288 15484
rect 5776 15444 5782 15456
rect 7282 15444 7288 15456
rect 7340 15444 7346 15496
rect 7650 15444 7656 15496
rect 7708 15484 7714 15496
rect 7837 15487 7895 15493
rect 7837 15484 7849 15487
rect 7708 15456 7849 15484
rect 7708 15444 7714 15456
rect 7837 15453 7849 15456
rect 7883 15453 7895 15487
rect 7837 15447 7895 15453
rect 8113 15487 8171 15493
rect 8113 15453 8125 15487
rect 8159 15484 8171 15487
rect 11330 15484 11336 15496
rect 8159 15456 11336 15484
rect 8159 15453 8171 15456
rect 8113 15447 8171 15453
rect 11330 15444 11336 15456
rect 11388 15444 11394 15496
rect 12158 15444 12164 15496
rect 12216 15484 12222 15496
rect 12345 15487 12403 15493
rect 12345 15484 12357 15487
rect 12216 15456 12357 15484
rect 12216 15444 12222 15456
rect 12345 15453 12357 15456
rect 12391 15453 12403 15487
rect 12345 15447 12403 15453
rect 14108 15425 14136 15592
rect 15930 15580 15936 15632
rect 15988 15620 15994 15632
rect 15988 15592 16712 15620
rect 15988 15580 15994 15592
rect 15105 15555 15163 15561
rect 15105 15521 15117 15555
rect 15151 15552 15163 15555
rect 15838 15552 15844 15564
rect 15151 15524 15844 15552
rect 15151 15521 15163 15524
rect 15105 15515 15163 15521
rect 15838 15512 15844 15524
rect 15896 15512 15902 15564
rect 16206 15552 16212 15564
rect 16167 15524 16212 15552
rect 16206 15512 16212 15524
rect 16264 15512 16270 15564
rect 16482 15552 16488 15564
rect 16443 15524 16488 15552
rect 16482 15512 16488 15524
rect 16540 15512 16546 15564
rect 16684 15561 16712 15592
rect 16669 15555 16727 15561
rect 16669 15521 16681 15555
rect 16715 15521 16727 15555
rect 16669 15515 16727 15521
rect 16942 15512 16948 15564
rect 17000 15552 17006 15564
rect 17129 15555 17187 15561
rect 17129 15552 17141 15555
rect 17000 15524 17141 15552
rect 17000 15512 17006 15524
rect 17129 15521 17141 15524
rect 17175 15521 17187 15555
rect 17129 15515 17187 15521
rect 17313 15555 17371 15561
rect 17313 15521 17325 15555
rect 17359 15552 17371 15555
rect 17402 15552 17408 15564
rect 17359 15524 17408 15552
rect 17359 15521 17371 15524
rect 17313 15515 17371 15521
rect 17402 15512 17408 15524
rect 17460 15512 17466 15564
rect 15010 15444 15016 15496
rect 15068 15484 15074 15496
rect 15197 15487 15255 15493
rect 15197 15484 15209 15487
rect 15068 15456 15209 15484
rect 15068 15444 15074 15456
rect 15197 15453 15209 15456
rect 15243 15453 15255 15487
rect 15197 15447 15255 15453
rect 15289 15487 15347 15493
rect 15289 15453 15301 15487
rect 15335 15453 15347 15487
rect 15930 15484 15936 15496
rect 15891 15456 15936 15484
rect 15289 15447 15347 15453
rect 14093 15419 14151 15425
rect 14093 15385 14105 15419
rect 14139 15385 14151 15419
rect 14093 15379 14151 15385
rect 8662 15348 8668 15360
rect 4816 15320 8668 15348
rect 8662 15308 8668 15320
rect 8720 15308 8726 15360
rect 9585 15351 9643 15357
rect 9585 15317 9597 15351
rect 9631 15348 9643 15351
rect 10134 15348 10140 15360
rect 9631 15320 10140 15348
rect 9631 15317 9643 15320
rect 9585 15311 9643 15317
rect 10134 15308 10140 15320
rect 10192 15308 10198 15360
rect 15102 15308 15108 15360
rect 15160 15348 15166 15360
rect 15304 15348 15332 15447
rect 15930 15444 15936 15456
rect 15988 15444 15994 15496
rect 15160 15320 15332 15348
rect 15160 15308 15166 15320
rect 16942 15308 16948 15360
rect 17000 15348 17006 15360
rect 17494 15348 17500 15360
rect 17000 15320 17500 15348
rect 17000 15308 17006 15320
rect 17494 15308 17500 15320
rect 17552 15348 17558 15360
rect 17589 15351 17647 15357
rect 17589 15348 17601 15351
rect 17552 15320 17601 15348
rect 17552 15308 17558 15320
rect 17589 15317 17601 15320
rect 17635 15317 17647 15351
rect 17589 15311 17647 15317
rect 184 15258 18860 15280
rect 184 15206 1556 15258
rect 1608 15206 1620 15258
rect 1672 15206 1684 15258
rect 1736 15206 1748 15258
rect 1800 15206 1812 15258
rect 1864 15206 4656 15258
rect 4708 15206 4720 15258
rect 4772 15206 4784 15258
rect 4836 15206 4848 15258
rect 4900 15206 4912 15258
rect 4964 15206 7756 15258
rect 7808 15206 7820 15258
rect 7872 15206 7884 15258
rect 7936 15206 7948 15258
rect 8000 15206 8012 15258
rect 8064 15206 10856 15258
rect 10908 15206 10920 15258
rect 10972 15206 10984 15258
rect 11036 15206 11048 15258
rect 11100 15206 11112 15258
rect 11164 15206 13956 15258
rect 14008 15206 14020 15258
rect 14072 15206 14084 15258
rect 14136 15206 14148 15258
rect 14200 15206 14212 15258
rect 14264 15206 17056 15258
rect 17108 15206 17120 15258
rect 17172 15206 17184 15258
rect 17236 15206 17248 15258
rect 17300 15206 17312 15258
rect 17364 15206 18860 15258
rect 184 15184 18860 15206
rect 5074 15144 5080 15156
rect 3436 15116 5080 15144
rect 2222 15008 2228 15020
rect 2135 14980 2228 15008
rect 2222 14968 2228 14980
rect 2280 15008 2286 15020
rect 3436 15008 3464 15116
rect 5074 15104 5080 15116
rect 5132 15104 5138 15156
rect 8297 15147 8355 15153
rect 8297 15113 8309 15147
rect 8343 15144 8355 15147
rect 8754 15144 8760 15156
rect 8343 15116 8760 15144
rect 8343 15113 8355 15116
rect 8297 15107 8355 15113
rect 8754 15104 8760 15116
rect 8812 15104 8818 15156
rect 15838 15104 15844 15156
rect 15896 15144 15902 15156
rect 15933 15147 15991 15153
rect 15933 15144 15945 15147
rect 15896 15116 15945 15144
rect 15896 15104 15902 15116
rect 15933 15113 15945 15116
rect 15979 15113 15991 15147
rect 15933 15107 15991 15113
rect 3513 15079 3571 15085
rect 3513 15045 3525 15079
rect 3559 15076 3571 15079
rect 3786 15076 3792 15088
rect 3559 15048 3792 15076
rect 3559 15045 3571 15048
rect 3513 15039 3571 15045
rect 3786 15036 3792 15048
rect 3844 15076 3850 15088
rect 5169 15079 5227 15085
rect 5169 15076 5181 15079
rect 3844 15048 5181 15076
rect 3844 15036 3850 15048
rect 5169 15045 5181 15048
rect 5215 15045 5227 15079
rect 5169 15039 5227 15045
rect 4709 15011 4767 15017
rect 2280 14980 3464 15008
rect 3528 14980 4563 15008
rect 2280 14968 2286 14980
rect 3528 14952 3556 14980
rect 2038 14940 2044 14952
rect 1999 14912 2044 14940
rect 2038 14900 2044 14912
rect 2096 14940 2102 14952
rect 2406 14940 2412 14952
rect 2096 14912 2412 14940
rect 2096 14900 2102 14912
rect 2406 14900 2412 14912
rect 2464 14940 2470 14952
rect 2685 14943 2743 14949
rect 2685 14940 2697 14943
rect 2464 14912 2697 14940
rect 2464 14900 2470 14912
rect 2685 14909 2697 14912
rect 2731 14940 2743 14943
rect 3421 14943 3479 14949
rect 2731 14912 3096 14940
rect 2731 14909 2743 14912
rect 2685 14903 2743 14909
rect 3068 14872 3096 14912
rect 3421 14909 3433 14943
rect 3467 14940 3479 14943
rect 3510 14940 3516 14952
rect 3467 14912 3516 14940
rect 3467 14909 3479 14912
rect 3421 14903 3479 14909
rect 3510 14900 3516 14912
rect 3568 14900 3574 14952
rect 3605 14943 3663 14949
rect 3605 14909 3617 14943
rect 3651 14940 3663 14943
rect 4430 14940 4436 14952
rect 3651 14912 4436 14940
rect 3651 14909 3663 14912
rect 3605 14903 3663 14909
rect 3620 14872 3648 14903
rect 4430 14900 4436 14912
rect 4488 14900 4494 14952
rect 4535 14949 4563 14980
rect 4709 14977 4721 15011
rect 4755 15008 4767 15011
rect 5353 15011 5411 15017
rect 5353 15008 5365 15011
rect 4755 14980 5365 15008
rect 4755 14977 4767 14980
rect 4709 14971 4767 14977
rect 5353 14977 5365 14980
rect 5399 15008 5411 15011
rect 7006 15008 7012 15020
rect 5399 14980 7012 15008
rect 5399 14977 5411 14980
rect 5353 14971 5411 14977
rect 7006 14968 7012 14980
rect 7064 14968 7070 15020
rect 7558 14968 7564 15020
rect 7616 15008 7622 15020
rect 7653 15011 7711 15017
rect 7653 15008 7665 15011
rect 7616 14980 7665 15008
rect 7616 14968 7622 14980
rect 7653 14977 7665 14980
rect 7699 14977 7711 15011
rect 14274 15008 14280 15020
rect 14235 14980 14280 15008
rect 7653 14971 7711 14977
rect 14274 14968 14280 14980
rect 14332 14968 14338 15020
rect 16114 14968 16120 15020
rect 16172 15008 16178 15020
rect 16485 15011 16543 15017
rect 16485 15008 16497 15011
rect 16172 14980 16497 15008
rect 16172 14968 16178 14980
rect 16485 14977 16497 14980
rect 16531 14977 16543 15011
rect 16485 14971 16543 14977
rect 4525 14943 4583 14949
rect 4525 14909 4537 14943
rect 4571 14909 4583 14943
rect 4525 14903 4583 14909
rect 4614 14900 4620 14952
rect 4672 14940 4678 14952
rect 5074 14940 5080 14952
rect 4672 14912 4717 14940
rect 5035 14912 5080 14940
rect 4672 14900 4678 14912
rect 5074 14900 5080 14912
rect 5132 14900 5138 14952
rect 5629 14943 5687 14949
rect 5629 14940 5641 14943
rect 5276 14912 5641 14940
rect 4154 14872 4160 14884
rect 3068 14844 3648 14872
rect 4115 14844 4160 14872
rect 4154 14832 4160 14844
rect 4212 14832 4218 14884
rect 4341 14875 4399 14881
rect 4341 14841 4353 14875
rect 4387 14872 4399 14875
rect 5276 14872 5304 14912
rect 5629 14909 5641 14912
rect 5675 14909 5687 14943
rect 5629 14903 5687 14909
rect 5813 14943 5871 14949
rect 5813 14909 5825 14943
rect 5859 14909 5871 14943
rect 5813 14903 5871 14909
rect 4387 14844 5304 14872
rect 5353 14875 5411 14881
rect 4387 14841 4399 14844
rect 4341 14835 4399 14841
rect 5353 14841 5365 14875
rect 5399 14872 5411 14875
rect 5828 14872 5856 14903
rect 7466 14900 7472 14952
rect 7524 14940 7530 14952
rect 7929 14943 7987 14949
rect 7929 14940 7941 14943
rect 7524 14912 7941 14940
rect 7524 14900 7530 14912
rect 7929 14909 7941 14912
rect 7975 14909 7987 14943
rect 7929 14903 7987 14909
rect 11149 14943 11207 14949
rect 11149 14909 11161 14943
rect 11195 14940 11207 14943
rect 11238 14940 11244 14952
rect 11195 14912 11244 14940
rect 11195 14909 11207 14912
rect 11149 14903 11207 14909
rect 11238 14900 11244 14912
rect 11296 14900 11302 14952
rect 11514 14940 11520 14952
rect 11475 14912 11520 14940
rect 11514 14900 11520 14912
rect 11572 14900 11578 14952
rect 13446 14900 13452 14952
rect 13504 14940 13510 14952
rect 13541 14943 13599 14949
rect 13541 14940 13553 14943
rect 13504 14912 13553 14940
rect 13504 14900 13510 14912
rect 13541 14909 13553 14912
rect 13587 14909 13599 14943
rect 13541 14903 13599 14909
rect 17405 14943 17463 14949
rect 17405 14909 17417 14943
rect 17451 14909 17463 14943
rect 17586 14940 17592 14952
rect 17547 14912 17592 14940
rect 17405 14903 17463 14909
rect 9030 14872 9036 14884
rect 5399 14844 5856 14872
rect 8991 14844 9036 14872
rect 5399 14841 5411 14844
rect 5353 14835 5411 14841
rect 9030 14832 9036 14844
rect 9088 14832 9094 14884
rect 11882 14872 11888 14884
rect 11808 14844 11888 14872
rect 934 14764 940 14816
rect 992 14804 998 14816
rect 1581 14807 1639 14813
rect 1581 14804 1593 14807
rect 992 14776 1593 14804
rect 992 14764 998 14776
rect 1581 14773 1593 14776
rect 1627 14773 1639 14807
rect 1946 14804 1952 14816
rect 1907 14776 1952 14804
rect 1581 14767 1639 14773
rect 1946 14764 1952 14776
rect 2004 14764 2010 14816
rect 2498 14764 2504 14816
rect 2556 14804 2562 14816
rect 2685 14807 2743 14813
rect 2685 14804 2697 14807
rect 2556 14776 2697 14804
rect 2556 14764 2562 14776
rect 2685 14773 2697 14776
rect 2731 14773 2743 14807
rect 5718 14804 5724 14816
rect 5679 14776 5724 14804
rect 2685 14767 2743 14773
rect 5718 14764 5724 14776
rect 5776 14764 5782 14816
rect 5810 14764 5816 14816
rect 5868 14804 5874 14816
rect 6365 14807 6423 14813
rect 6365 14804 6377 14807
rect 5868 14776 6377 14804
rect 5868 14764 5874 14776
rect 6365 14773 6377 14776
rect 6411 14773 6423 14807
rect 7834 14804 7840 14816
rect 7795 14776 7840 14804
rect 6365 14767 6423 14773
rect 7834 14764 7840 14776
rect 7892 14764 7898 14816
rect 10318 14804 10324 14816
rect 10279 14776 10324 14804
rect 10318 14764 10324 14776
rect 10376 14764 10382 14816
rect 11146 14764 11152 14816
rect 11204 14804 11210 14816
rect 11808 14804 11836 14844
rect 11882 14832 11888 14844
rect 11940 14832 11946 14884
rect 17420 14872 17448 14903
rect 17586 14900 17592 14912
rect 17644 14900 17650 14952
rect 17954 14872 17960 14884
rect 17420 14844 17960 14872
rect 17954 14832 17960 14844
rect 18012 14832 18018 14884
rect 11204 14776 11836 14804
rect 11204 14764 11210 14776
rect 12802 14764 12808 14816
rect 12860 14804 12866 14816
rect 12943 14807 13001 14813
rect 12943 14804 12955 14807
rect 12860 14776 12955 14804
rect 12860 14764 12866 14776
rect 12943 14773 12955 14776
rect 12989 14773 13001 14807
rect 12943 14767 13001 14773
rect 15930 14764 15936 14816
rect 15988 14804 15994 14816
rect 16114 14804 16120 14816
rect 15988 14776 16120 14804
rect 15988 14764 15994 14776
rect 16114 14764 16120 14776
rect 16172 14804 16178 14816
rect 16301 14807 16359 14813
rect 16301 14804 16313 14807
rect 16172 14776 16313 14804
rect 16172 14764 16178 14776
rect 16301 14773 16313 14776
rect 16347 14773 16359 14807
rect 16301 14767 16359 14773
rect 16390 14764 16396 14816
rect 16448 14804 16454 14816
rect 16448 14776 16493 14804
rect 16448 14764 16454 14776
rect 17126 14764 17132 14816
rect 17184 14804 17190 14816
rect 17402 14804 17408 14816
rect 17184 14776 17408 14804
rect 17184 14764 17190 14776
rect 17402 14764 17408 14776
rect 17460 14804 17466 14816
rect 17497 14807 17555 14813
rect 17497 14804 17509 14807
rect 17460 14776 17509 14804
rect 17460 14764 17466 14776
rect 17497 14773 17509 14776
rect 17543 14773 17555 14807
rect 17497 14767 17555 14773
rect 184 14714 18920 14736
rect 184 14662 3106 14714
rect 3158 14662 3170 14714
rect 3222 14662 3234 14714
rect 3286 14662 3298 14714
rect 3350 14662 3362 14714
rect 3414 14662 6206 14714
rect 6258 14662 6270 14714
rect 6322 14662 6334 14714
rect 6386 14662 6398 14714
rect 6450 14662 6462 14714
rect 6514 14662 9306 14714
rect 9358 14662 9370 14714
rect 9422 14662 9434 14714
rect 9486 14662 9498 14714
rect 9550 14662 9562 14714
rect 9614 14662 12406 14714
rect 12458 14662 12470 14714
rect 12522 14662 12534 14714
rect 12586 14662 12598 14714
rect 12650 14662 12662 14714
rect 12714 14662 15506 14714
rect 15558 14662 15570 14714
rect 15622 14662 15634 14714
rect 15686 14662 15698 14714
rect 15750 14662 15762 14714
rect 15814 14662 18606 14714
rect 18658 14662 18670 14714
rect 18722 14662 18734 14714
rect 18786 14662 18798 14714
rect 18850 14662 18862 14714
rect 18914 14662 18920 14714
rect 184 14640 18920 14662
rect 2958 14560 2964 14612
rect 3016 14600 3022 14612
rect 3237 14603 3295 14609
rect 3237 14600 3249 14603
rect 3016 14572 3249 14600
rect 3016 14560 3022 14572
rect 3237 14569 3249 14572
rect 3283 14569 3295 14603
rect 3694 14600 3700 14612
rect 3655 14572 3700 14600
rect 3237 14563 3295 14569
rect 3694 14560 3700 14572
rect 3752 14560 3758 14612
rect 11057 14603 11115 14609
rect 11057 14569 11069 14603
rect 11103 14600 11115 14603
rect 11422 14600 11428 14612
rect 11103 14572 11428 14600
rect 11103 14569 11115 14572
rect 11057 14563 11115 14569
rect 2130 14532 2136 14544
rect 1978 14504 2136 14532
rect 2130 14492 2136 14504
rect 2188 14492 2194 14544
rect 2406 14532 2412 14544
rect 2367 14504 2412 14532
rect 2406 14492 2412 14504
rect 2464 14492 2470 14544
rect 6730 14492 6736 14544
rect 6788 14492 6794 14544
rect 8478 14492 8484 14544
rect 8536 14492 8542 14544
rect 566 14464 572 14476
rect 527 14436 572 14464
rect 566 14424 572 14436
rect 624 14424 630 14476
rect 934 14464 940 14476
rect 895 14436 940 14464
rect 934 14424 940 14436
rect 992 14424 998 14476
rect 3605 14467 3663 14473
rect 3605 14433 3617 14467
rect 3651 14464 3663 14467
rect 3694 14464 3700 14476
rect 3651 14436 3700 14464
rect 3651 14433 3663 14436
rect 3605 14427 3663 14433
rect 3694 14424 3700 14436
rect 3752 14424 3758 14476
rect 4522 14424 4528 14476
rect 4580 14464 4586 14476
rect 5353 14467 5411 14473
rect 5353 14464 5365 14467
rect 4580 14436 5365 14464
rect 4580 14424 4586 14436
rect 5353 14433 5365 14436
rect 5399 14464 5411 14467
rect 5442 14464 5448 14476
rect 5399 14436 5448 14464
rect 5399 14433 5411 14436
rect 5353 14427 5411 14433
rect 5442 14424 5448 14436
rect 5500 14424 5506 14476
rect 5718 14464 5724 14476
rect 5679 14436 5724 14464
rect 5718 14424 5724 14436
rect 5776 14424 5782 14476
rect 7745 14467 7803 14473
rect 7745 14433 7757 14467
rect 7791 14464 7803 14467
rect 7834 14464 7840 14476
rect 7791 14436 7840 14464
rect 7791 14433 7803 14436
rect 7745 14427 7803 14433
rect 7834 14424 7840 14436
rect 7892 14464 7898 14476
rect 8202 14464 8208 14476
rect 7892 14436 8208 14464
rect 7892 14424 7898 14436
rect 8202 14424 8208 14436
rect 8260 14424 8266 14476
rect 10689 14467 10747 14473
rect 10689 14433 10701 14467
rect 10735 14464 10747 14467
rect 11072 14464 11100 14563
rect 11422 14560 11428 14572
rect 11480 14560 11486 14612
rect 11882 14560 11888 14612
rect 11940 14600 11946 14612
rect 14921 14603 14979 14609
rect 11940 14572 13032 14600
rect 11940 14560 11946 14572
rect 11330 14532 11336 14544
rect 11291 14504 11336 14532
rect 11330 14492 11336 14504
rect 11388 14492 11394 14544
rect 13004 14532 13032 14572
rect 14921 14569 14933 14603
rect 14967 14600 14979 14603
rect 16390 14600 16396 14612
rect 14967 14572 16396 14600
rect 14967 14569 14979 14572
rect 14921 14563 14979 14569
rect 16390 14560 16396 14572
rect 16448 14560 16454 14612
rect 13078 14532 13084 14544
rect 13004 14504 13084 14532
rect 13078 14492 13084 14504
rect 13136 14492 13142 14544
rect 15657 14535 15715 14541
rect 15657 14501 15669 14535
rect 15703 14532 15715 14535
rect 16482 14532 16488 14544
rect 15703 14504 16488 14532
rect 15703 14501 15715 14504
rect 15657 14495 15715 14501
rect 16482 14492 16488 14504
rect 16540 14492 16546 14544
rect 17144 14504 18000 14532
rect 10735 14436 11100 14464
rect 10735 14433 10747 14436
rect 10689 14427 10747 14433
rect 11238 14424 11244 14476
rect 11296 14464 11302 14476
rect 12158 14464 12164 14476
rect 11296 14436 12164 14464
rect 11296 14424 11302 14436
rect 12158 14424 12164 14436
rect 12216 14464 12222 14476
rect 12345 14467 12403 14473
rect 12345 14464 12357 14467
rect 12216 14436 12357 14464
rect 12216 14424 12222 14436
rect 12345 14433 12357 14436
rect 12391 14433 12403 14467
rect 12345 14427 12403 14433
rect 12713 14467 12771 14473
rect 12713 14433 12725 14467
rect 12759 14464 12771 14467
rect 12802 14464 12808 14476
rect 12759 14436 12808 14464
rect 12759 14433 12771 14436
rect 12713 14427 12771 14433
rect 12802 14424 12808 14436
rect 12860 14424 12866 14476
rect 15010 14464 15016 14476
rect 14971 14436 15016 14464
rect 15010 14424 15016 14436
rect 15068 14464 15074 14476
rect 15746 14464 15752 14476
rect 15068 14436 15752 14464
rect 15068 14424 15074 14436
rect 15746 14424 15752 14436
rect 15804 14424 15810 14476
rect 15841 14467 15899 14473
rect 15841 14433 15853 14467
rect 15887 14433 15899 14467
rect 15841 14427 15899 14433
rect 3786 14396 3792 14408
rect 3747 14368 3792 14396
rect 3786 14356 3792 14368
rect 3844 14356 3850 14408
rect 8110 14396 8116 14408
rect 8071 14368 8116 14396
rect 8110 14356 8116 14368
rect 8168 14356 8174 14408
rect 10505 14399 10563 14405
rect 10505 14365 10517 14399
rect 10551 14396 10563 14399
rect 11146 14396 11152 14408
rect 10551 14368 11152 14396
rect 10551 14365 10563 14368
rect 10505 14359 10563 14365
rect 11146 14356 11152 14368
rect 11204 14356 11210 14408
rect 11330 14356 11336 14408
rect 11388 14396 11394 14408
rect 11388 14368 13492 14396
rect 11388 14356 11394 14368
rect 13464 14328 13492 14368
rect 15194 14356 15200 14408
rect 15252 14396 15258 14408
rect 15473 14399 15531 14405
rect 15473 14396 15485 14399
rect 15252 14368 15485 14396
rect 15252 14356 15258 14368
rect 15473 14365 15485 14368
rect 15519 14365 15531 14399
rect 15473 14359 15531 14365
rect 15562 14328 15568 14340
rect 13464 14300 15568 14328
rect 15562 14288 15568 14300
rect 15620 14288 15626 14340
rect 15856 14328 15884 14427
rect 15930 14424 15936 14476
rect 15988 14464 15994 14476
rect 17144 14473 17172 14504
rect 17972 14476 18000 14504
rect 17129 14467 17187 14473
rect 15988 14436 16574 14464
rect 15988 14424 15994 14436
rect 16022 14396 16028 14408
rect 15983 14368 16028 14396
rect 16022 14356 16028 14368
rect 16080 14356 16086 14408
rect 16546 14396 16574 14436
rect 17129 14433 17141 14467
rect 17175 14433 17187 14467
rect 17129 14427 17187 14433
rect 17589 14467 17647 14473
rect 17589 14433 17601 14467
rect 17635 14464 17647 14467
rect 17862 14464 17868 14476
rect 17635 14436 17868 14464
rect 17635 14433 17647 14436
rect 17589 14427 17647 14433
rect 17862 14424 17868 14436
rect 17920 14424 17926 14476
rect 17954 14424 17960 14476
rect 18012 14464 18018 14476
rect 18233 14467 18291 14473
rect 18233 14464 18245 14467
rect 18012 14436 18245 14464
rect 18012 14424 18018 14436
rect 18233 14433 18245 14436
rect 18279 14433 18291 14467
rect 18233 14427 18291 14433
rect 16850 14396 16856 14408
rect 16546 14368 16856 14396
rect 16850 14356 16856 14368
rect 16908 14356 16914 14408
rect 17221 14399 17279 14405
rect 17221 14365 17233 14399
rect 17267 14396 17279 14399
rect 17402 14396 17408 14408
rect 17267 14368 17408 14396
rect 17267 14365 17279 14368
rect 17221 14359 17279 14365
rect 17402 14356 17408 14368
rect 17460 14356 17466 14408
rect 17126 14328 17132 14340
rect 15856 14300 17132 14328
rect 17126 14288 17132 14300
rect 17184 14288 17190 14340
rect 18049 14331 18107 14337
rect 18049 14328 18061 14331
rect 17328 14300 18061 14328
rect 7006 14220 7012 14272
rect 7064 14260 7070 14272
rect 7147 14263 7205 14269
rect 7147 14260 7159 14263
rect 7064 14232 7159 14260
rect 7064 14220 7070 14232
rect 7147 14229 7159 14232
rect 7193 14260 7205 14263
rect 7374 14260 7380 14272
rect 7193 14232 7380 14260
rect 7193 14229 7205 14232
rect 7147 14223 7205 14229
rect 7374 14220 7380 14232
rect 7432 14220 7438 14272
rect 7466 14220 7472 14272
rect 7524 14260 7530 14272
rect 9539 14263 9597 14269
rect 9539 14260 9551 14263
rect 7524 14232 9551 14260
rect 7524 14220 7530 14232
rect 9539 14229 9551 14232
rect 9585 14229 9597 14263
rect 9539 14223 9597 14229
rect 11790 14220 11796 14272
rect 11848 14260 11854 14272
rect 12894 14260 12900 14272
rect 11848 14232 12900 14260
rect 11848 14220 11854 14232
rect 12894 14220 12900 14232
rect 12952 14220 12958 14272
rect 14139 14263 14197 14269
rect 14139 14229 14151 14263
rect 14185 14260 14197 14263
rect 15010 14260 15016 14272
rect 14185 14232 15016 14260
rect 14185 14229 14197 14232
rect 14139 14223 14197 14229
rect 15010 14220 15016 14232
rect 15068 14260 15074 14272
rect 16206 14260 16212 14272
rect 15068 14232 16212 14260
rect 15068 14220 15074 14232
rect 16206 14220 16212 14232
rect 16264 14220 16270 14272
rect 16850 14220 16856 14272
rect 16908 14260 16914 14272
rect 17328 14269 17356 14300
rect 18049 14297 18061 14300
rect 18095 14297 18107 14331
rect 18049 14291 18107 14297
rect 17313 14263 17371 14269
rect 17313 14260 17325 14263
rect 16908 14232 17325 14260
rect 16908 14220 16914 14232
rect 17313 14229 17325 14232
rect 17359 14229 17371 14263
rect 17313 14223 17371 14229
rect 17451 14263 17509 14269
rect 17451 14229 17463 14263
rect 17497 14260 17509 14263
rect 17586 14260 17592 14272
rect 17497 14232 17592 14260
rect 17497 14229 17509 14232
rect 17451 14223 17509 14229
rect 17586 14220 17592 14232
rect 17644 14260 17650 14272
rect 17957 14263 18015 14269
rect 17957 14260 17969 14263
rect 17644 14232 17969 14260
rect 17644 14220 17650 14232
rect 17957 14229 17969 14232
rect 18003 14229 18015 14263
rect 18230 14260 18236 14272
rect 18191 14232 18236 14260
rect 17957 14223 18015 14229
rect 18230 14220 18236 14232
rect 18288 14220 18294 14272
rect 184 14170 18860 14192
rect 184 14118 1556 14170
rect 1608 14118 1620 14170
rect 1672 14118 1684 14170
rect 1736 14118 1748 14170
rect 1800 14118 1812 14170
rect 1864 14118 4656 14170
rect 4708 14118 4720 14170
rect 4772 14118 4784 14170
rect 4836 14118 4848 14170
rect 4900 14118 4912 14170
rect 4964 14118 7756 14170
rect 7808 14118 7820 14170
rect 7872 14118 7884 14170
rect 7936 14118 7948 14170
rect 8000 14118 8012 14170
rect 8064 14118 10856 14170
rect 10908 14118 10920 14170
rect 10972 14118 10984 14170
rect 11036 14118 11048 14170
rect 11100 14118 11112 14170
rect 11164 14118 13956 14170
rect 14008 14118 14020 14170
rect 14072 14118 14084 14170
rect 14136 14118 14148 14170
rect 14200 14118 14212 14170
rect 14264 14118 17056 14170
rect 17108 14118 17120 14170
rect 17172 14118 17184 14170
rect 17236 14118 17248 14170
rect 17300 14118 17312 14170
rect 17364 14118 18860 14170
rect 184 14096 18860 14118
rect 1946 14016 1952 14068
rect 2004 14056 2010 14068
rect 2041 14059 2099 14065
rect 2041 14056 2053 14059
rect 2004 14028 2053 14056
rect 2004 14016 2010 14028
rect 2041 14025 2053 14028
rect 2087 14025 2099 14059
rect 2041 14019 2099 14025
rect 5629 14059 5687 14065
rect 5629 14025 5641 14059
rect 5675 14056 5687 14059
rect 5810 14056 5816 14068
rect 5675 14028 5816 14056
rect 5675 14025 5687 14028
rect 5629 14019 5687 14025
rect 5810 14016 5816 14028
rect 5868 14056 5874 14068
rect 6638 14056 6644 14068
rect 5868 14028 6644 14056
rect 5868 14016 5874 14028
rect 6638 14016 6644 14028
rect 6696 14016 6702 14068
rect 8662 14016 8668 14068
rect 8720 14056 8726 14068
rect 8757 14059 8815 14065
rect 8757 14056 8769 14059
rect 8720 14028 8769 14056
rect 8720 14016 8726 14028
rect 8757 14025 8769 14028
rect 8803 14025 8815 14059
rect 8757 14019 8815 14025
rect 10134 14016 10140 14068
rect 10192 14056 10198 14068
rect 10241 14059 10299 14065
rect 10241 14056 10253 14059
rect 10192 14028 10253 14056
rect 10192 14016 10198 14028
rect 10241 14025 10253 14028
rect 10287 14025 10299 14059
rect 10241 14019 10299 14025
rect 11514 14016 11520 14068
rect 11572 14056 11578 14068
rect 17773 14059 17831 14065
rect 17773 14056 17785 14059
rect 11572 14028 17785 14056
rect 11572 14016 11578 14028
rect 17773 14025 17785 14028
rect 17819 14025 17831 14059
rect 17773 14019 17831 14025
rect 12250 13948 12256 14000
rect 12308 13988 12314 14000
rect 12713 13991 12771 13997
rect 12713 13988 12725 13991
rect 12308 13960 12725 13988
rect 12308 13948 12314 13960
rect 12713 13957 12725 13960
rect 12759 13957 12771 13991
rect 14274 13988 14280 14000
rect 12713 13951 12771 13957
rect 12820 13960 14280 13988
rect 2498 13920 2504 13932
rect 2459 13892 2504 13920
rect 2498 13880 2504 13892
rect 2556 13880 2562 13932
rect 2685 13923 2743 13929
rect 2685 13889 2697 13923
rect 2731 13920 2743 13923
rect 3786 13920 3792 13932
rect 2731 13892 3792 13920
rect 2731 13889 2743 13892
rect 2685 13883 2743 13889
rect 3786 13880 3792 13892
rect 3844 13880 3850 13932
rect 6656 13892 7236 13920
rect 2590 13852 2596 13864
rect 2424 13824 2596 13852
rect 2424 13793 2452 13824
rect 2590 13812 2596 13824
rect 2648 13852 2654 13864
rect 6656 13852 6684 13892
rect 2648 13824 6684 13852
rect 6733 13855 6791 13861
rect 2648 13812 2654 13824
rect 6733 13821 6745 13855
rect 6779 13852 6791 13855
rect 6822 13852 6828 13864
rect 6779 13824 6828 13852
rect 6779 13821 6791 13824
rect 6733 13815 6791 13821
rect 2409 13787 2467 13793
rect 2409 13753 2421 13787
rect 2455 13753 2467 13787
rect 2409 13747 2467 13753
rect 5074 13744 5080 13796
rect 5132 13784 5138 13796
rect 6748 13784 6776 13815
rect 6822 13812 6828 13824
rect 6880 13812 6886 13864
rect 7098 13852 7104 13864
rect 7059 13824 7104 13852
rect 7098 13812 7104 13824
rect 7156 13812 7162 13864
rect 7208 13852 7236 13892
rect 8202 13880 8208 13932
rect 8260 13920 8266 13932
rect 10505 13923 10563 13929
rect 10505 13920 10517 13923
rect 8260 13892 10517 13920
rect 8260 13880 8266 13892
rect 10505 13889 10517 13892
rect 10551 13889 10563 13923
rect 10505 13883 10563 13889
rect 11885 13923 11943 13929
rect 11885 13889 11897 13923
rect 11931 13920 11943 13923
rect 12820 13920 12848 13960
rect 14274 13948 14280 13960
rect 14332 13948 14338 14000
rect 15286 13948 15292 14000
rect 15344 13948 15350 14000
rect 15562 13948 15568 14000
rect 15620 13988 15626 14000
rect 18138 13988 18144 14000
rect 15620 13960 18144 13988
rect 15620 13948 15626 13960
rect 18138 13948 18144 13960
rect 18196 13948 18202 14000
rect 11931 13892 12296 13920
rect 11931 13889 11943 13892
rect 11885 13883 11943 13889
rect 7466 13852 7472 13864
rect 7208 13824 7472 13852
rect 7466 13812 7472 13824
rect 7524 13812 7530 13864
rect 11790 13852 11796 13864
rect 11751 13824 11796 13852
rect 11790 13812 11796 13824
rect 11848 13812 11854 13864
rect 12268 13861 12296 13892
rect 12636 13892 12848 13920
rect 14001 13923 14059 13929
rect 12636 13861 12664 13892
rect 14001 13889 14013 13923
rect 14047 13920 14059 13923
rect 15194 13920 15200 13932
rect 14047 13892 15200 13920
rect 14047 13889 14059 13892
rect 14001 13883 14059 13889
rect 15194 13880 15200 13892
rect 15252 13880 15258 13932
rect 15304 13920 15332 13948
rect 16942 13920 16948 13932
rect 15304 13892 15976 13920
rect 11977 13855 12035 13861
rect 11977 13821 11989 13855
rect 12023 13821 12035 13855
rect 11977 13815 12035 13821
rect 12253 13855 12311 13861
rect 12253 13821 12265 13855
rect 12299 13821 12311 13855
rect 12253 13815 12311 13821
rect 12621 13855 12679 13861
rect 12621 13821 12633 13855
rect 12667 13821 12679 13855
rect 12802 13852 12808 13864
rect 12763 13824 12808 13852
rect 12621 13815 12679 13821
rect 5132 13756 6776 13784
rect 6917 13787 6975 13793
rect 5132 13744 5138 13756
rect 6917 13753 6929 13787
rect 6963 13784 6975 13787
rect 7190 13784 7196 13796
rect 6963 13756 7196 13784
rect 6963 13753 6975 13756
rect 6917 13747 6975 13753
rect 7190 13744 7196 13756
rect 7248 13744 7254 13796
rect 7745 13787 7803 13793
rect 7745 13753 7757 13787
rect 7791 13784 7803 13787
rect 8205 13787 8263 13793
rect 8205 13784 8217 13787
rect 7791 13756 8217 13784
rect 7791 13753 7803 13756
rect 7745 13747 7803 13753
rect 8205 13753 8217 13756
rect 8251 13753 8263 13787
rect 8205 13747 8263 13753
rect 5997 13719 6055 13725
rect 5997 13685 6009 13719
rect 6043 13716 6055 13719
rect 6822 13716 6828 13728
rect 6043 13688 6828 13716
rect 6043 13685 6055 13688
rect 5997 13679 6055 13685
rect 6822 13676 6828 13688
rect 6880 13716 6886 13728
rect 7760 13716 7788 13747
rect 8478 13744 8484 13796
rect 8536 13784 8542 13796
rect 8938 13784 8944 13796
rect 8536 13756 8944 13784
rect 8536 13744 8542 13756
rect 8938 13744 8944 13756
rect 8996 13784 9002 13796
rect 11992 13784 12020 13815
rect 12802 13812 12808 13824
rect 12860 13812 12866 13864
rect 13081 13855 13139 13861
rect 13081 13821 13093 13855
rect 13127 13852 13139 13855
rect 14826 13852 14832 13864
rect 13127 13824 14832 13852
rect 13127 13821 13139 13824
rect 13081 13815 13139 13821
rect 14826 13812 14832 13824
rect 14884 13812 14890 13864
rect 14918 13812 14924 13864
rect 14976 13852 14982 13864
rect 15948 13861 15976 13892
rect 16546 13892 16948 13920
rect 15013 13855 15071 13861
rect 15013 13852 15025 13855
rect 14976 13824 15025 13852
rect 14976 13812 14982 13824
rect 15013 13821 15025 13824
rect 15059 13821 15071 13855
rect 15013 13815 15071 13821
rect 15289 13855 15347 13861
rect 15289 13821 15301 13855
rect 15335 13852 15347 13855
rect 15933 13855 15991 13861
rect 15335 13824 15884 13852
rect 15335 13821 15347 13824
rect 15289 13815 15347 13821
rect 13722 13784 13728 13796
rect 8996 13756 9062 13784
rect 11992 13756 13728 13784
rect 8996 13744 9002 13756
rect 13722 13744 13728 13756
rect 13780 13744 13786 13796
rect 13814 13744 13820 13796
rect 13872 13784 13878 13796
rect 14093 13787 14151 13793
rect 14093 13784 14105 13787
rect 13872 13756 14105 13784
rect 13872 13744 13878 13756
rect 14093 13753 14105 13756
rect 14139 13753 14151 13787
rect 14093 13747 14151 13753
rect 14185 13787 14243 13793
rect 14185 13753 14197 13787
rect 14231 13784 14243 13787
rect 15856 13784 15884 13824
rect 15933 13821 15945 13855
rect 15979 13821 15991 13855
rect 16298 13852 16304 13864
rect 15933 13815 15991 13821
rect 16040 13824 16304 13852
rect 16040 13784 16068 13824
rect 16298 13812 16304 13824
rect 16356 13812 16362 13864
rect 16206 13784 16212 13796
rect 14231 13756 14964 13784
rect 15856 13756 16068 13784
rect 16167 13756 16212 13784
rect 14231 13753 14243 13756
rect 14185 13747 14243 13753
rect 6880 13688 7788 13716
rect 14553 13719 14611 13725
rect 6880 13676 6886 13688
rect 14553 13685 14565 13719
rect 14599 13716 14611 13719
rect 14734 13716 14740 13728
rect 14599 13688 14740 13716
rect 14599 13685 14611 13688
rect 14553 13679 14611 13685
rect 14734 13676 14740 13688
rect 14792 13676 14798 13728
rect 14936 13716 14964 13756
rect 16206 13744 16212 13756
rect 16264 13784 16270 13796
rect 16546 13784 16574 13892
rect 16942 13880 16948 13892
rect 17000 13880 17006 13932
rect 18230 13920 18236 13932
rect 17512 13892 18236 13920
rect 17402 13852 17408 13864
rect 17363 13824 17408 13852
rect 17402 13812 17408 13824
rect 17460 13812 17466 13864
rect 17512 13861 17540 13892
rect 18230 13880 18236 13892
rect 18288 13880 18294 13932
rect 17497 13855 17555 13861
rect 17497 13821 17509 13855
rect 17543 13821 17555 13855
rect 17497 13815 17555 13821
rect 17957 13855 18015 13861
rect 17957 13821 17969 13855
rect 18003 13852 18015 13855
rect 18417 13855 18475 13861
rect 18417 13852 18429 13855
rect 18003 13824 18429 13852
rect 18003 13821 18015 13824
rect 17957 13815 18015 13821
rect 18417 13821 18429 13824
rect 18463 13852 18475 13855
rect 19058 13852 19064 13864
rect 18463 13824 19064 13852
rect 18463 13821 18475 13824
rect 18417 13815 18475 13821
rect 19058 13812 19064 13824
rect 19116 13812 19122 13864
rect 16264 13756 16574 13784
rect 16264 13744 16270 13756
rect 16022 13716 16028 13728
rect 14936 13688 16028 13716
rect 16022 13676 16028 13688
rect 16080 13676 16086 13728
rect 16850 13676 16856 13728
rect 16908 13716 16914 13728
rect 17129 13719 17187 13725
rect 17129 13716 17141 13719
rect 16908 13688 17141 13716
rect 16908 13676 16914 13688
rect 17129 13685 17141 13688
rect 17175 13685 17187 13719
rect 17129 13679 17187 13685
rect 184 13626 18920 13648
rect 184 13574 3106 13626
rect 3158 13574 3170 13626
rect 3222 13574 3234 13626
rect 3286 13574 3298 13626
rect 3350 13574 3362 13626
rect 3414 13574 6206 13626
rect 6258 13574 6270 13626
rect 6322 13574 6334 13626
rect 6386 13574 6398 13626
rect 6450 13574 6462 13626
rect 6514 13574 9306 13626
rect 9358 13574 9370 13626
rect 9422 13574 9434 13626
rect 9486 13574 9498 13626
rect 9550 13574 9562 13626
rect 9614 13574 12406 13626
rect 12458 13574 12470 13626
rect 12522 13574 12534 13626
rect 12586 13574 12598 13626
rect 12650 13574 12662 13626
rect 12714 13574 15506 13626
rect 15558 13574 15570 13626
rect 15622 13574 15634 13626
rect 15686 13574 15698 13626
rect 15750 13574 15762 13626
rect 15814 13574 18606 13626
rect 18658 13574 18670 13626
rect 18722 13574 18734 13626
rect 18786 13574 18798 13626
rect 18850 13574 18862 13626
rect 18914 13574 18920 13626
rect 184 13552 18920 13574
rect 7791 13515 7849 13521
rect 7791 13481 7803 13515
rect 7837 13512 7849 13515
rect 8018 13512 8024 13524
rect 7837 13484 8024 13512
rect 7837 13481 7849 13484
rect 7791 13475 7849 13481
rect 8018 13472 8024 13484
rect 8076 13472 8082 13524
rect 10689 13515 10747 13521
rect 10689 13481 10701 13515
rect 10735 13512 10747 13515
rect 11238 13512 11244 13524
rect 10735 13484 11244 13512
rect 10735 13481 10747 13484
rect 10689 13475 10747 13481
rect 11238 13472 11244 13484
rect 11296 13472 11302 13524
rect 13081 13515 13139 13521
rect 13081 13481 13093 13515
rect 13127 13512 13139 13515
rect 13814 13512 13820 13524
rect 13127 13484 13820 13512
rect 13127 13481 13139 13484
rect 13081 13475 13139 13481
rect 13814 13472 13820 13484
rect 13872 13472 13878 13524
rect 15194 13472 15200 13524
rect 15252 13512 15258 13524
rect 15657 13515 15715 13521
rect 15657 13512 15669 13515
rect 15252 13484 15669 13512
rect 15252 13472 15258 13484
rect 15657 13481 15669 13484
rect 15703 13481 15715 13515
rect 15657 13475 15715 13481
rect 4522 13444 4528 13456
rect 3436 13416 4528 13444
rect 3436 13385 3464 13416
rect 4522 13404 4528 13416
rect 4580 13404 4586 13456
rect 6086 13444 6092 13456
rect 5276 13416 6092 13444
rect 3694 13385 3700 13388
rect 3421 13379 3479 13385
rect 3421 13376 3433 13379
rect 2746 13348 3433 13376
rect 566 13268 572 13320
rect 624 13308 630 13320
rect 2746 13308 2774 13348
rect 3421 13345 3433 13348
rect 3467 13345 3479 13379
rect 3688 13376 3700 13385
rect 3655 13348 3700 13376
rect 3421 13339 3479 13345
rect 3688 13339 3700 13348
rect 3752 13376 3758 13388
rect 5276 13376 5304 13416
rect 6086 13404 6092 13416
rect 6144 13444 6150 13456
rect 6546 13444 6552 13456
rect 6144 13416 6224 13444
rect 6144 13404 6150 13416
rect 5442 13376 5448 13388
rect 3752 13348 5304 13376
rect 5403 13348 5448 13376
rect 3694 13336 3700 13339
rect 3752 13336 3758 13348
rect 5442 13336 5448 13348
rect 5500 13336 5506 13388
rect 6196 13385 6224 13416
rect 6380 13416 6552 13444
rect 6380 13385 6408 13416
rect 6546 13404 6552 13416
rect 6604 13444 6610 13456
rect 6822 13444 6828 13456
rect 6604 13416 6828 13444
rect 6604 13404 6610 13416
rect 6822 13404 6828 13416
rect 6880 13444 6886 13456
rect 11974 13444 11980 13456
rect 6880 13416 7052 13444
rect 6880 13404 6886 13416
rect 6181 13379 6239 13385
rect 6181 13345 6193 13379
rect 6227 13345 6239 13379
rect 6181 13339 6239 13345
rect 6365 13379 6423 13385
rect 6365 13345 6377 13379
rect 6411 13345 6423 13379
rect 6638 13376 6644 13388
rect 6599 13348 6644 13376
rect 6365 13339 6423 13345
rect 6638 13336 6644 13348
rect 6696 13336 6702 13388
rect 6730 13336 6736 13388
rect 6788 13376 6794 13388
rect 7024 13385 7052 13416
rect 7009 13379 7067 13385
rect 6788 13348 6960 13376
rect 6788 13336 6794 13348
rect 5718 13308 5724 13320
rect 624 13280 2774 13308
rect 5679 13280 5724 13308
rect 624 13268 630 13280
rect 5718 13268 5724 13280
rect 5776 13268 5782 13320
rect 5994 13268 6000 13320
rect 6052 13308 6058 13320
rect 6825 13311 6883 13317
rect 6825 13308 6837 13311
rect 6052 13280 6837 13308
rect 6052 13268 6058 13280
rect 6825 13277 6837 13280
rect 6871 13277 6883 13311
rect 6932 13308 6960 13348
rect 7009 13345 7021 13379
rect 7055 13345 7067 13379
rect 7009 13339 7067 13345
rect 8220 13308 8248 13430
rect 11935 13416 11980 13444
rect 11974 13404 11980 13416
rect 12032 13404 12038 13456
rect 14642 13404 14648 13456
rect 14700 13444 14706 13456
rect 14700 13416 15792 13444
rect 14700 13404 14706 13416
rect 14366 13376 14372 13388
rect 14327 13348 14372 13376
rect 14366 13336 14372 13348
rect 14424 13336 14430 13388
rect 14734 13376 14740 13388
rect 14695 13348 14740 13376
rect 14734 13336 14740 13348
rect 14792 13336 14798 13388
rect 14918 13336 14924 13388
rect 14976 13376 14982 13388
rect 15764 13385 15792 13416
rect 15197 13379 15255 13385
rect 15197 13376 15209 13379
rect 14976 13348 15209 13376
rect 14976 13336 14982 13348
rect 15197 13345 15209 13348
rect 15243 13345 15255 13379
rect 15197 13339 15255 13345
rect 15565 13379 15623 13385
rect 15565 13345 15577 13379
rect 15611 13345 15623 13379
rect 15565 13339 15623 13345
rect 15749 13379 15807 13385
rect 15749 13345 15761 13379
rect 15795 13376 15807 13379
rect 16206 13376 16212 13388
rect 15795 13348 16212 13376
rect 15795 13345 15807 13348
rect 15749 13339 15807 13345
rect 6932 13280 8248 13308
rect 6825 13271 6883 13277
rect 8846 13268 8852 13320
rect 8904 13308 8910 13320
rect 9217 13311 9275 13317
rect 9217 13308 9229 13311
rect 8904 13280 9229 13308
rect 8904 13268 8910 13280
rect 9217 13277 9229 13280
rect 9263 13277 9275 13311
rect 9217 13271 9275 13277
rect 9306 13268 9312 13320
rect 9364 13308 9370 13320
rect 9585 13311 9643 13317
rect 9585 13308 9597 13311
rect 9364 13280 9597 13308
rect 9364 13268 9370 13280
rect 9585 13277 9597 13280
rect 9631 13277 9643 13311
rect 14826 13308 14832 13320
rect 14787 13280 14832 13308
rect 9585 13271 9643 13277
rect 14826 13268 14832 13280
rect 14884 13268 14890 13320
rect 15010 13268 15016 13320
rect 15068 13308 15074 13320
rect 15580 13308 15608 13339
rect 16206 13336 16212 13348
rect 16264 13376 16270 13388
rect 16393 13379 16451 13385
rect 16393 13376 16405 13379
rect 16264 13348 16405 13376
rect 16264 13336 16270 13348
rect 16393 13345 16405 13348
rect 16439 13345 16451 13379
rect 16393 13339 16451 13345
rect 16298 13308 16304 13320
rect 15068 13280 16304 13308
rect 15068 13268 15074 13280
rect 16298 13268 16304 13280
rect 16356 13268 16362 13320
rect 4801 13243 4859 13249
rect 4801 13209 4813 13243
rect 4847 13240 4859 13243
rect 5074 13240 5080 13252
rect 4847 13212 5080 13240
rect 4847 13209 4859 13212
rect 4801 13203 4859 13209
rect 5074 13200 5080 13212
rect 5132 13200 5138 13252
rect 6914 13240 6920 13252
rect 6875 13212 6920 13240
rect 6914 13200 6920 13212
rect 6972 13200 6978 13252
rect 4982 13132 4988 13184
rect 5040 13172 5046 13184
rect 5537 13175 5595 13181
rect 5537 13172 5549 13175
rect 5040 13144 5549 13172
rect 5040 13132 5046 13144
rect 5537 13141 5549 13144
rect 5583 13141 5595 13175
rect 5537 13135 5595 13141
rect 5626 13132 5632 13184
rect 5684 13172 5690 13184
rect 6365 13175 6423 13181
rect 5684 13144 5729 13172
rect 5684 13132 5690 13144
rect 6365 13141 6377 13175
rect 6411 13172 6423 13175
rect 7650 13172 7656 13184
rect 6411 13144 7656 13172
rect 6411 13141 6423 13144
rect 6365 13135 6423 13141
rect 7650 13132 7656 13144
rect 7708 13132 7714 13184
rect 16117 13175 16175 13181
rect 16117 13141 16129 13175
rect 16163 13172 16175 13175
rect 16206 13172 16212 13184
rect 16163 13144 16212 13172
rect 16163 13141 16175 13144
rect 16117 13135 16175 13141
rect 16206 13132 16212 13144
rect 16264 13132 16270 13184
rect 184 13082 18860 13104
rect 184 13030 1556 13082
rect 1608 13030 1620 13082
rect 1672 13030 1684 13082
rect 1736 13030 1748 13082
rect 1800 13030 1812 13082
rect 1864 13030 4656 13082
rect 4708 13030 4720 13082
rect 4772 13030 4784 13082
rect 4836 13030 4848 13082
rect 4900 13030 4912 13082
rect 4964 13030 7756 13082
rect 7808 13030 7820 13082
rect 7872 13030 7884 13082
rect 7936 13030 7948 13082
rect 8000 13030 8012 13082
rect 8064 13030 10856 13082
rect 10908 13030 10920 13082
rect 10972 13030 10984 13082
rect 11036 13030 11048 13082
rect 11100 13030 11112 13082
rect 11164 13030 13956 13082
rect 14008 13030 14020 13082
rect 14072 13030 14084 13082
rect 14136 13030 14148 13082
rect 14200 13030 14212 13082
rect 14264 13030 17056 13082
rect 17108 13030 17120 13082
rect 17172 13030 17184 13082
rect 17236 13030 17248 13082
rect 17300 13030 17312 13082
rect 17364 13030 18860 13082
rect 184 13008 18860 13030
rect 4341 12971 4399 12977
rect 4341 12937 4353 12971
rect 4387 12937 4399 12971
rect 4982 12968 4988 12980
rect 4943 12940 4988 12968
rect 4341 12931 4399 12937
rect 4356 12900 4384 12931
rect 4982 12928 4988 12940
rect 5040 12928 5046 12980
rect 7006 12928 7012 12980
rect 7064 12968 7070 12980
rect 7469 12971 7527 12977
rect 7064 12940 7420 12968
rect 7064 12928 7070 12940
rect 5442 12900 5448 12912
rect 4356 12872 5448 12900
rect 5442 12860 5448 12872
rect 5500 12860 5506 12912
rect 7282 12832 7288 12844
rect 4356 12804 4844 12832
rect 4356 12773 4384 12804
rect 4816 12773 4844 12804
rect 6932 12804 7288 12832
rect 6932 12776 6960 12804
rect 7282 12792 7288 12804
rect 7340 12792 7346 12844
rect 7392 12832 7420 12940
rect 7469 12937 7481 12971
rect 7515 12968 7527 12971
rect 9030 12968 9036 12980
rect 7515 12940 9036 12968
rect 7515 12937 7527 12940
rect 7469 12931 7527 12937
rect 9030 12928 9036 12940
rect 9088 12928 9094 12980
rect 12802 12928 12808 12980
rect 12860 12968 12866 12980
rect 13541 12971 13599 12977
rect 13541 12968 13553 12971
rect 12860 12940 13553 12968
rect 12860 12928 12866 12940
rect 13541 12937 13553 12940
rect 13587 12937 13599 12971
rect 17954 12968 17960 12980
rect 17915 12940 17960 12968
rect 13541 12931 13599 12937
rect 17954 12928 17960 12940
rect 18012 12928 18018 12980
rect 7745 12835 7803 12841
rect 7745 12832 7757 12835
rect 7392 12804 7757 12832
rect 7745 12801 7757 12804
rect 7791 12801 7803 12835
rect 7745 12795 7803 12801
rect 9214 12792 9220 12844
rect 9272 12832 9278 12844
rect 10505 12835 10563 12841
rect 10505 12832 10517 12835
rect 9272 12804 10517 12832
rect 9272 12792 9278 12804
rect 10505 12801 10517 12804
rect 10551 12801 10563 12835
rect 10505 12795 10563 12801
rect 13814 12792 13820 12844
rect 13872 12832 13878 12844
rect 14185 12835 14243 12841
rect 14185 12832 14197 12835
rect 13872 12804 14197 12832
rect 13872 12792 13878 12804
rect 14185 12801 14197 12804
rect 14231 12801 14243 12835
rect 14185 12795 14243 12801
rect 16485 12835 16543 12841
rect 16485 12801 16497 12835
rect 16531 12832 16543 12835
rect 16850 12832 16856 12844
rect 16531 12804 16856 12832
rect 16531 12801 16543 12804
rect 16485 12795 16543 12801
rect 4157 12767 4215 12773
rect 4157 12733 4169 12767
rect 4203 12733 4215 12767
rect 4157 12727 4215 12733
rect 4341 12767 4399 12773
rect 4341 12733 4353 12767
rect 4387 12733 4399 12767
rect 4341 12727 4399 12733
rect 4709 12767 4767 12773
rect 4709 12733 4721 12767
rect 4755 12733 4767 12767
rect 4709 12727 4767 12733
rect 4801 12767 4859 12773
rect 4801 12733 4813 12767
rect 4847 12764 4859 12767
rect 5074 12764 5080 12776
rect 4847 12736 5080 12764
rect 4847 12733 4859 12736
rect 4801 12727 4859 12733
rect 4172 12696 4200 12727
rect 4724 12696 4752 12727
rect 5074 12724 5080 12736
rect 5132 12724 5138 12776
rect 5994 12764 6000 12776
rect 5276 12736 6000 12764
rect 5276 12696 5304 12736
rect 5994 12724 6000 12736
rect 6052 12724 6058 12776
rect 6638 12764 6644 12776
rect 6599 12736 6644 12764
rect 6638 12724 6644 12736
rect 6696 12724 6702 12776
rect 6914 12764 6920 12776
rect 6875 12736 6920 12764
rect 6914 12724 6920 12736
rect 6972 12724 6978 12776
rect 7006 12724 7012 12776
rect 7064 12764 7070 12776
rect 7101 12767 7159 12773
rect 7101 12764 7113 12767
rect 7064 12736 7113 12764
rect 7064 12724 7070 12736
rect 7101 12733 7113 12736
rect 7147 12733 7159 12767
rect 7101 12727 7159 12733
rect 7190 12724 7196 12776
rect 7248 12764 7254 12776
rect 7469 12767 7527 12773
rect 7469 12764 7481 12767
rect 7248 12736 7481 12764
rect 7248 12724 7254 12736
rect 7469 12733 7481 12736
rect 7515 12733 7527 12767
rect 7469 12727 7527 12733
rect 7929 12767 7987 12773
rect 7929 12733 7941 12767
rect 7975 12764 7987 12767
rect 8662 12764 8668 12776
rect 7975 12736 8668 12764
rect 7975 12733 7987 12736
rect 7929 12727 7987 12733
rect 8662 12724 8668 12736
rect 8720 12724 8726 12776
rect 11146 12764 11152 12776
rect 11107 12736 11152 12764
rect 11146 12724 11152 12736
rect 11204 12724 11210 12776
rect 11514 12764 11520 12776
rect 11475 12736 11520 12764
rect 11514 12724 11520 12736
rect 11572 12724 11578 12776
rect 13722 12764 13728 12776
rect 13683 12736 13728 12764
rect 13722 12724 13728 12736
rect 13780 12724 13786 12776
rect 13909 12767 13967 12773
rect 13909 12733 13921 12767
rect 13955 12733 13967 12767
rect 14200 12764 14228 12795
rect 16850 12792 16856 12804
rect 16908 12792 16914 12844
rect 16114 12764 16120 12776
rect 14200 12736 16120 12764
rect 13909 12727 13967 12733
rect 4172 12668 5304 12696
rect 5629 12699 5687 12705
rect 5629 12665 5641 12699
rect 5675 12696 5687 12699
rect 5675 12668 6960 12696
rect 5675 12665 5687 12668
rect 5629 12659 5687 12665
rect 6932 12640 6960 12668
rect 8938 12656 8944 12708
rect 8996 12696 9002 12708
rect 8996 12668 9062 12696
rect 8996 12656 9002 12668
rect 9950 12656 9956 12708
rect 10008 12696 10014 12708
rect 10229 12699 10287 12705
rect 10229 12696 10241 12699
rect 10008 12668 10241 12696
rect 10008 12656 10014 12668
rect 10229 12665 10241 12668
rect 10275 12665 10287 12699
rect 11882 12696 11888 12708
rect 10229 12659 10287 12665
rect 11808 12668 11888 12696
rect 4338 12588 4344 12640
rect 4396 12628 4402 12640
rect 5353 12631 5411 12637
rect 5353 12628 5365 12631
rect 4396 12600 5365 12628
rect 4396 12588 4402 12600
rect 5353 12597 5365 12600
rect 5399 12597 5411 12631
rect 5353 12591 5411 12597
rect 6914 12588 6920 12640
rect 6972 12588 6978 12640
rect 8662 12588 8668 12640
rect 8720 12628 8726 12640
rect 8757 12631 8815 12637
rect 8757 12628 8769 12631
rect 8720 12600 8769 12628
rect 8720 12588 8726 12600
rect 8757 12597 8769 12600
rect 8803 12597 8815 12631
rect 11808 12628 11836 12668
rect 11882 12656 11888 12668
rect 11940 12656 11946 12708
rect 12894 12696 12900 12708
rect 12853 12668 12900 12696
rect 12894 12656 12900 12668
rect 12952 12705 12958 12708
rect 12952 12699 13001 12705
rect 12952 12665 12955 12699
rect 12989 12696 13001 12699
rect 13924 12696 13952 12727
rect 16114 12724 16120 12736
rect 16172 12764 16178 12776
rect 16209 12767 16267 12773
rect 16209 12764 16221 12767
rect 16172 12736 16221 12764
rect 16172 12724 16178 12736
rect 16209 12733 16221 12736
rect 16255 12733 16267 12767
rect 16209 12727 16267 12733
rect 12989 12668 13952 12696
rect 14452 12699 14510 12705
rect 12989 12665 13001 12668
rect 12952 12659 13001 12665
rect 14452 12665 14464 12699
rect 14498 12696 14510 12699
rect 15194 12696 15200 12708
rect 14498 12668 15200 12696
rect 14498 12665 14510 12668
rect 14452 12659 14510 12665
rect 12952 12656 12958 12659
rect 15194 12656 15200 12668
rect 15252 12656 15258 12708
rect 16224 12668 16974 12696
rect 16224 12640 16252 12668
rect 12250 12628 12256 12640
rect 11808 12600 12256 12628
rect 8757 12591 8815 12597
rect 12250 12588 12256 12600
rect 12308 12588 12314 12640
rect 15286 12588 15292 12640
rect 15344 12628 15350 12640
rect 15565 12631 15623 12637
rect 15565 12628 15577 12631
rect 15344 12600 15577 12628
rect 15344 12588 15350 12600
rect 15565 12597 15577 12600
rect 15611 12597 15623 12631
rect 15565 12591 15623 12597
rect 16206 12588 16212 12640
rect 16264 12588 16270 12640
rect 184 12538 18920 12560
rect 184 12486 3106 12538
rect 3158 12486 3170 12538
rect 3222 12486 3234 12538
rect 3286 12486 3298 12538
rect 3350 12486 3362 12538
rect 3414 12486 6206 12538
rect 6258 12486 6270 12538
rect 6322 12486 6334 12538
rect 6386 12486 6398 12538
rect 6450 12486 6462 12538
rect 6514 12486 9306 12538
rect 9358 12486 9370 12538
rect 9422 12486 9434 12538
rect 9486 12486 9498 12538
rect 9550 12486 9562 12538
rect 9614 12486 12406 12538
rect 12458 12486 12470 12538
rect 12522 12486 12534 12538
rect 12586 12486 12598 12538
rect 12650 12486 12662 12538
rect 12714 12486 15506 12538
rect 15558 12486 15570 12538
rect 15622 12486 15634 12538
rect 15686 12486 15698 12538
rect 15750 12486 15762 12538
rect 15814 12486 18606 12538
rect 18658 12486 18670 12538
rect 18722 12486 18734 12538
rect 18786 12486 18798 12538
rect 18850 12486 18862 12538
rect 18914 12486 18920 12538
rect 184 12464 18920 12486
rect 7558 12384 7564 12436
rect 7616 12424 7622 12436
rect 7837 12427 7895 12433
rect 7837 12424 7849 12427
rect 7616 12396 7849 12424
rect 7616 12384 7622 12396
rect 7837 12393 7849 12396
rect 7883 12393 7895 12427
rect 7837 12387 7895 12393
rect 10781 12427 10839 12433
rect 10781 12393 10793 12427
rect 10827 12424 10839 12427
rect 11514 12424 11520 12436
rect 10827 12396 11520 12424
rect 10827 12393 10839 12396
rect 10781 12387 10839 12393
rect 11514 12384 11520 12396
rect 11572 12384 11578 12436
rect 12250 12384 12256 12436
rect 12308 12424 12314 12436
rect 16850 12424 16856 12436
rect 12308 12396 16856 12424
rect 12308 12384 12314 12396
rect 16850 12384 16856 12396
rect 16908 12384 16914 12436
rect 17221 12427 17279 12433
rect 17221 12393 17233 12427
rect 17267 12424 17279 12427
rect 17954 12424 17960 12436
rect 17267 12396 17960 12424
rect 17267 12393 17279 12396
rect 17221 12387 17279 12393
rect 17954 12384 17960 12396
rect 18012 12424 18018 12436
rect 18506 12424 18512 12436
rect 18012 12396 18512 12424
rect 18012 12384 18018 12396
rect 18506 12384 18512 12396
rect 18564 12384 18570 12436
rect 3145 12359 3203 12365
rect 2608 12328 2912 12356
rect 2608 12300 2636 12328
rect 566 12248 572 12300
rect 624 12288 630 12300
rect 1029 12291 1087 12297
rect 1029 12288 1041 12291
rect 624 12260 1041 12288
rect 624 12248 630 12260
rect 1029 12257 1041 12260
rect 1075 12288 1087 12291
rect 1118 12288 1124 12300
rect 1075 12260 1124 12288
rect 1075 12257 1087 12260
rect 1029 12251 1087 12257
rect 1118 12248 1124 12260
rect 1176 12248 1182 12300
rect 1296 12291 1354 12297
rect 1296 12257 1308 12291
rect 1342 12288 1354 12291
rect 2222 12288 2228 12300
rect 1342 12260 2228 12288
rect 1342 12257 1354 12260
rect 1296 12251 1354 12257
rect 2222 12248 2228 12260
rect 2280 12288 2286 12300
rect 2590 12288 2596 12300
rect 2280 12260 2596 12288
rect 2280 12248 2286 12260
rect 2590 12248 2596 12260
rect 2648 12248 2654 12300
rect 2884 12297 2912 12328
rect 3145 12325 3157 12359
rect 3191 12356 3203 12359
rect 3605 12359 3663 12365
rect 3605 12356 3617 12359
rect 3191 12328 3617 12356
rect 3191 12325 3203 12328
rect 3145 12319 3203 12325
rect 3605 12325 3617 12328
rect 3651 12325 3663 12359
rect 3605 12319 3663 12325
rect 8570 12316 8576 12368
rect 8628 12316 8634 12368
rect 11146 12316 11152 12368
rect 11204 12356 11210 12368
rect 11241 12359 11299 12365
rect 11241 12356 11253 12359
rect 11204 12328 11253 12356
rect 11204 12316 11210 12328
rect 11241 12325 11253 12328
rect 11287 12325 11299 12359
rect 13814 12356 13820 12368
rect 11241 12319 11299 12325
rect 11624 12328 13820 12356
rect 2777 12291 2835 12297
rect 2777 12257 2789 12291
rect 2823 12257 2835 12291
rect 2777 12251 2835 12257
rect 2870 12291 2928 12297
rect 2870 12257 2882 12291
rect 2916 12257 2928 12291
rect 2870 12251 2928 12257
rect 2406 12152 2412 12164
rect 2319 12124 2412 12152
rect 2406 12112 2412 12124
rect 2464 12152 2470 12164
rect 2792 12152 2820 12251
rect 2958 12248 2964 12300
rect 3016 12288 3022 12300
rect 3421 12291 3479 12297
rect 3421 12288 3433 12291
rect 3016 12260 3433 12288
rect 3016 12248 3022 12260
rect 3421 12257 3433 12260
rect 3467 12257 3479 12291
rect 3421 12251 3479 12257
rect 3510 12248 3516 12300
rect 3568 12288 3574 12300
rect 3697 12291 3755 12297
rect 3697 12288 3709 12291
rect 3568 12260 3709 12288
rect 3568 12248 3574 12260
rect 3697 12257 3709 12260
rect 3743 12257 3755 12291
rect 3697 12251 3755 12257
rect 6917 12291 6975 12297
rect 6917 12257 6929 12291
rect 6963 12288 6975 12291
rect 7190 12288 7196 12300
rect 6963 12260 7196 12288
rect 6963 12257 6975 12260
rect 6917 12251 6975 12257
rect 7190 12248 7196 12260
rect 7248 12248 7254 12300
rect 10594 12288 10600 12300
rect 10555 12260 10600 12288
rect 10594 12248 10600 12260
rect 10652 12248 10658 12300
rect 10778 12288 10784 12300
rect 10739 12260 10784 12288
rect 10778 12248 10784 12260
rect 10836 12248 10842 12300
rect 11624 12297 11652 12328
rect 13814 12316 13820 12328
rect 13872 12316 13878 12368
rect 14093 12359 14151 12365
rect 14093 12325 14105 12359
rect 14139 12356 14151 12359
rect 15102 12356 15108 12368
rect 14139 12328 15108 12356
rect 14139 12325 14151 12328
rect 14093 12319 14151 12325
rect 15102 12316 15108 12328
rect 15160 12316 15166 12368
rect 11609 12291 11667 12297
rect 11609 12257 11621 12291
rect 11655 12257 11667 12291
rect 11609 12251 11667 12257
rect 12805 12291 12863 12297
rect 12805 12257 12817 12291
rect 12851 12288 12863 12291
rect 12894 12288 12900 12300
rect 12851 12260 12900 12288
rect 12851 12257 12863 12260
rect 12805 12251 12863 12257
rect 12894 12248 12900 12260
rect 12952 12248 12958 12300
rect 13725 12291 13783 12297
rect 13725 12257 13737 12291
rect 13771 12288 13783 12291
rect 15010 12288 15016 12300
rect 13771 12260 15016 12288
rect 13771 12257 13783 12260
rect 13725 12251 13783 12257
rect 15010 12248 15016 12260
rect 15068 12248 15074 12300
rect 15194 12288 15200 12300
rect 15155 12260 15200 12288
rect 15194 12248 15200 12260
rect 15252 12248 15258 12300
rect 15286 12248 15292 12300
rect 15344 12288 15350 12300
rect 15381 12291 15439 12297
rect 15381 12288 15393 12291
rect 15344 12260 15393 12288
rect 15344 12248 15350 12260
rect 15381 12257 15393 12260
rect 15427 12288 15439 12291
rect 15841 12291 15899 12297
rect 15841 12288 15853 12291
rect 15427 12260 15853 12288
rect 15427 12257 15439 12260
rect 15381 12251 15439 12257
rect 15841 12257 15853 12260
rect 15887 12257 15899 12291
rect 16301 12291 16359 12297
rect 16301 12288 16313 12291
rect 15841 12251 15899 12257
rect 15948 12260 16313 12288
rect 5166 12220 5172 12232
rect 5127 12192 5172 12220
rect 5166 12180 5172 12192
rect 5224 12180 5230 12232
rect 8570 12180 8576 12232
rect 8628 12220 8634 12232
rect 9309 12223 9367 12229
rect 9309 12220 9321 12223
rect 8628 12192 9321 12220
rect 8628 12180 8634 12192
rect 9309 12189 9321 12192
rect 9355 12189 9367 12223
rect 9309 12183 9367 12189
rect 9585 12223 9643 12229
rect 9585 12189 9597 12223
rect 9631 12189 9643 12223
rect 9585 12183 9643 12189
rect 13909 12223 13967 12229
rect 13909 12189 13921 12223
rect 13955 12220 13967 12223
rect 14642 12220 14648 12232
rect 13955 12192 14648 12220
rect 13955 12189 13967 12192
rect 13909 12183 13967 12189
rect 2464 12124 2820 12152
rect 2464 12112 2470 12124
rect 3694 12084 3700 12096
rect 3655 12056 3700 12084
rect 3694 12044 3700 12056
rect 3752 12044 3758 12096
rect 7558 12044 7564 12096
rect 7616 12084 7622 12096
rect 9600 12084 9628 12183
rect 14642 12180 14648 12192
rect 14700 12220 14706 12232
rect 14737 12223 14795 12229
rect 14737 12220 14749 12223
rect 14700 12192 14749 12220
rect 14700 12180 14706 12192
rect 14737 12189 14749 12192
rect 14783 12189 14795 12223
rect 15212 12220 15240 12248
rect 15657 12223 15715 12229
rect 15657 12220 15669 12223
rect 15212 12192 15669 12220
rect 14737 12183 14795 12189
rect 15657 12189 15669 12192
rect 15703 12189 15715 12223
rect 15657 12183 15715 12189
rect 13814 12152 13820 12164
rect 13775 12124 13820 12152
rect 13814 12112 13820 12124
rect 13872 12152 13878 12164
rect 14274 12152 14280 12164
rect 13872 12124 14280 12152
rect 13872 12112 13878 12124
rect 14274 12112 14280 12124
rect 14332 12112 14338 12164
rect 15381 12155 15439 12161
rect 15381 12121 15393 12155
rect 15427 12152 15439 12155
rect 15948 12152 15976 12260
rect 16301 12257 16313 12260
rect 16347 12257 16359 12291
rect 16301 12251 16359 12257
rect 16574 12220 16580 12232
rect 16535 12192 16580 12220
rect 16574 12180 16580 12192
rect 16632 12180 16638 12232
rect 15427 12124 15976 12152
rect 15427 12121 15439 12124
rect 15381 12115 15439 12121
rect 7616 12056 9628 12084
rect 7616 12044 7622 12056
rect 11606 12044 11612 12096
rect 11664 12084 11670 12096
rect 12437 12087 12495 12093
rect 12437 12084 12449 12087
rect 11664 12056 12449 12084
rect 11664 12044 11670 12056
rect 12437 12053 12449 12056
rect 12483 12053 12495 12087
rect 12437 12047 12495 12053
rect 16025 12087 16083 12093
rect 16025 12053 16037 12087
rect 16071 12084 16083 12087
rect 16393 12087 16451 12093
rect 16393 12084 16405 12087
rect 16071 12056 16405 12084
rect 16071 12053 16083 12056
rect 16025 12047 16083 12053
rect 16393 12053 16405 12056
rect 16439 12053 16451 12087
rect 16393 12047 16451 12053
rect 16485 12087 16543 12093
rect 16485 12053 16497 12087
rect 16531 12084 16543 12087
rect 16942 12084 16948 12096
rect 16531 12056 16948 12084
rect 16531 12053 16543 12056
rect 16485 12047 16543 12053
rect 16942 12044 16948 12056
rect 17000 12044 17006 12096
rect 184 11994 18860 12016
rect 184 11942 1556 11994
rect 1608 11942 1620 11994
rect 1672 11942 1684 11994
rect 1736 11942 1748 11994
rect 1800 11942 1812 11994
rect 1864 11942 4656 11994
rect 4708 11942 4720 11994
rect 4772 11942 4784 11994
rect 4836 11942 4848 11994
rect 4900 11942 4912 11994
rect 4964 11942 7756 11994
rect 7808 11942 7820 11994
rect 7872 11942 7884 11994
rect 7936 11942 7948 11994
rect 8000 11942 8012 11994
rect 8064 11942 10856 11994
rect 10908 11942 10920 11994
rect 10972 11942 10984 11994
rect 11036 11942 11048 11994
rect 11100 11942 11112 11994
rect 11164 11942 13956 11994
rect 14008 11942 14020 11994
rect 14072 11942 14084 11994
rect 14136 11942 14148 11994
rect 14200 11942 14212 11994
rect 14264 11942 17056 11994
rect 17108 11942 17120 11994
rect 17172 11942 17184 11994
rect 17236 11942 17248 11994
rect 17300 11942 17312 11994
rect 17364 11942 18860 11994
rect 184 11920 18860 11942
rect 4154 11840 4160 11892
rect 4212 11880 4218 11892
rect 4249 11883 4307 11889
rect 4249 11880 4261 11883
rect 4212 11852 4261 11880
rect 4212 11840 4218 11852
rect 4249 11849 4261 11852
rect 4295 11849 4307 11883
rect 4249 11843 4307 11849
rect 4709 11883 4767 11889
rect 4709 11849 4721 11883
rect 4755 11880 4767 11883
rect 5534 11880 5540 11892
rect 4755 11852 5540 11880
rect 4755 11849 4767 11852
rect 4709 11843 4767 11849
rect 2593 11815 2651 11821
rect 2593 11781 2605 11815
rect 2639 11812 2651 11815
rect 3510 11812 3516 11824
rect 2639 11784 3516 11812
rect 2639 11781 2651 11784
rect 2593 11775 2651 11781
rect 3510 11772 3516 11784
rect 3568 11772 3574 11824
rect 4264 11744 4292 11843
rect 5534 11840 5540 11852
rect 5592 11880 5598 11892
rect 5718 11880 5724 11892
rect 5592 11852 5724 11880
rect 5592 11840 5598 11852
rect 5718 11840 5724 11852
rect 5776 11840 5782 11892
rect 7098 11880 7104 11892
rect 7059 11852 7104 11880
rect 7098 11840 7104 11852
rect 7156 11840 7162 11892
rect 7190 11840 7196 11892
rect 7248 11880 7254 11892
rect 8205 11883 8263 11889
rect 8205 11880 8217 11883
rect 7248 11852 8217 11880
rect 7248 11840 7254 11852
rect 8205 11849 8217 11852
rect 8251 11880 8263 11883
rect 15378 11880 15384 11892
rect 8251 11852 15384 11880
rect 8251 11849 8263 11852
rect 8205 11843 8263 11849
rect 15378 11840 15384 11852
rect 15436 11840 15442 11892
rect 18230 11880 18236 11892
rect 15488 11852 18236 11880
rect 4522 11772 4528 11824
rect 4580 11812 4586 11824
rect 4580 11784 7604 11812
rect 4580 11772 4586 11784
rect 5258 11744 5264 11756
rect 4264 11716 5264 11744
rect 5258 11704 5264 11716
rect 5316 11744 5322 11756
rect 6546 11744 6552 11756
rect 5316 11716 5764 11744
rect 5316 11704 5322 11716
rect 2222 11676 2228 11688
rect 2183 11648 2228 11676
rect 2222 11636 2228 11648
rect 2280 11636 2286 11688
rect 2406 11685 2412 11688
rect 2379 11679 2412 11685
rect 2379 11645 2391 11679
rect 2379 11639 2412 11645
rect 2406 11636 2412 11639
rect 2464 11636 2470 11688
rect 4338 11636 4344 11688
rect 4396 11676 4402 11688
rect 4617 11679 4675 11685
rect 4617 11676 4629 11679
rect 4396 11648 4629 11676
rect 4396 11636 4402 11648
rect 4617 11645 4629 11648
rect 4663 11645 4675 11679
rect 4617 11639 4675 11645
rect 4893 11679 4951 11685
rect 4893 11645 4905 11679
rect 4939 11645 4951 11679
rect 4893 11639 4951 11645
rect 4985 11679 5043 11685
rect 4985 11645 4997 11679
rect 5031 11676 5043 11679
rect 5626 11676 5632 11688
rect 5031 11648 5632 11676
rect 5031 11645 5043 11648
rect 4985 11639 5043 11645
rect 3694 11568 3700 11620
rect 3752 11608 3758 11620
rect 4908 11608 4936 11639
rect 5626 11636 5632 11648
rect 5684 11636 5690 11688
rect 5736 11685 5764 11716
rect 5920 11716 6552 11744
rect 5920 11685 5948 11716
rect 6546 11704 6552 11716
rect 6604 11704 6610 11756
rect 7576 11753 7604 11784
rect 10778 11772 10784 11824
rect 10836 11812 10842 11824
rect 11149 11815 11207 11821
rect 11149 11812 11161 11815
rect 10836 11784 11161 11812
rect 10836 11772 10842 11784
rect 11149 11781 11161 11784
rect 11195 11781 11207 11815
rect 11698 11812 11704 11824
rect 11149 11775 11207 11781
rect 11440 11784 11704 11812
rect 7561 11747 7619 11753
rect 7561 11713 7573 11747
rect 7607 11713 7619 11747
rect 7561 11707 7619 11713
rect 7650 11704 7656 11756
rect 7708 11744 7714 11756
rect 7708 11716 7753 11744
rect 7708 11704 7714 11716
rect 8294 11704 8300 11756
rect 8352 11744 8358 11756
rect 9214 11744 9220 11756
rect 8352 11716 9220 11744
rect 8352 11704 8358 11716
rect 9214 11704 9220 11716
rect 9272 11744 9278 11756
rect 10505 11747 10563 11753
rect 10505 11744 10517 11747
rect 9272 11716 10517 11744
rect 9272 11704 9278 11716
rect 10505 11713 10517 11716
rect 10551 11713 10563 11747
rect 10505 11707 10563 11713
rect 5721 11679 5779 11685
rect 5721 11645 5733 11679
rect 5767 11645 5779 11679
rect 5721 11639 5779 11645
rect 5905 11679 5963 11685
rect 5905 11645 5917 11679
rect 5951 11645 5963 11679
rect 5905 11639 5963 11645
rect 5920 11608 5948 11639
rect 5994 11636 6000 11688
rect 6052 11676 6058 11688
rect 6825 11679 6883 11685
rect 6825 11676 6837 11679
rect 6052 11648 6592 11676
rect 6052 11636 6058 11648
rect 6564 11620 6592 11648
rect 6656 11648 6837 11676
rect 6546 11608 6552 11620
rect 3752 11580 4936 11608
rect 5000 11580 5948 11608
rect 6507 11580 6552 11608
rect 3752 11568 3758 11580
rect 5000 11552 5028 11580
rect 6546 11568 6552 11580
rect 6604 11568 6610 11620
rect 6656 11608 6684 11648
rect 6825 11645 6837 11648
rect 6871 11645 6883 11679
rect 6825 11639 6883 11645
rect 7374 11636 7380 11688
rect 7432 11676 7438 11688
rect 7469 11679 7527 11685
rect 7469 11676 7481 11679
rect 7432 11648 7481 11676
rect 7432 11636 7438 11648
rect 7469 11645 7481 11648
rect 7515 11645 7527 11679
rect 11330 11676 11336 11688
rect 11291 11648 11336 11676
rect 7469 11639 7527 11645
rect 11330 11636 11336 11648
rect 11388 11636 11394 11688
rect 11440 11685 11468 11784
rect 11698 11772 11704 11784
rect 11756 11772 11762 11824
rect 11517 11747 11575 11753
rect 11517 11713 11529 11747
rect 11563 11744 11575 11747
rect 11790 11744 11796 11756
rect 11563 11716 11796 11744
rect 11563 11713 11575 11716
rect 11517 11707 11575 11713
rect 11790 11704 11796 11716
rect 11848 11744 11854 11756
rect 11848 11716 12434 11744
rect 11848 11704 11854 11716
rect 11425 11679 11483 11685
rect 11425 11645 11437 11679
rect 11471 11645 11483 11679
rect 11606 11676 11612 11688
rect 11567 11648 11612 11676
rect 11425 11639 11483 11645
rect 11606 11636 11612 11648
rect 11664 11636 11670 11688
rect 12406 11676 12434 11716
rect 15102 11676 15108 11688
rect 12406 11648 15108 11676
rect 15102 11636 15108 11648
rect 15160 11636 15166 11688
rect 8662 11608 8668 11620
rect 6656 11580 8668 11608
rect 4982 11500 4988 11552
rect 5040 11500 5046 11552
rect 5169 11543 5227 11549
rect 5169 11509 5181 11543
rect 5215 11540 5227 11543
rect 5442 11540 5448 11552
rect 5215 11512 5448 11540
rect 5215 11509 5227 11512
rect 5169 11503 5227 11509
rect 5442 11500 5448 11512
rect 5500 11500 5506 11552
rect 6086 11500 6092 11552
rect 6144 11540 6150 11552
rect 6656 11540 6684 11580
rect 8662 11568 8668 11580
rect 8720 11568 8726 11620
rect 8938 11568 8944 11620
rect 8996 11608 9002 11620
rect 10229 11611 10287 11617
rect 8996 11580 9062 11608
rect 8996 11568 9002 11580
rect 10229 11577 10241 11611
rect 10275 11608 10287 11611
rect 15488 11608 15516 11852
rect 18230 11840 18236 11852
rect 18288 11840 18294 11892
rect 16114 11744 16120 11756
rect 16075 11716 16120 11744
rect 16114 11704 16120 11716
rect 16172 11704 16178 11756
rect 17954 11744 17960 11756
rect 16408 11716 17960 11744
rect 15565 11679 15623 11685
rect 15565 11645 15577 11679
rect 15611 11676 15623 11679
rect 16408 11676 16436 11716
rect 17954 11704 17960 11716
rect 18012 11704 18018 11756
rect 15611 11648 16436 11676
rect 15611 11645 15623 11648
rect 15565 11639 15623 11645
rect 16482 11636 16488 11688
rect 16540 11676 16546 11688
rect 16540 11648 16585 11676
rect 16540 11636 16546 11648
rect 10275 11580 15516 11608
rect 10275 11577 10287 11580
rect 10229 11571 10287 11577
rect 16850 11568 16856 11620
rect 16908 11568 16914 11620
rect 6144 11512 6684 11540
rect 8757 11543 8815 11549
rect 6144 11500 6150 11512
rect 8757 11509 8769 11543
rect 8803 11540 8815 11543
rect 9950 11540 9956 11552
rect 8803 11512 9956 11540
rect 8803 11509 8815 11512
rect 8757 11503 8815 11509
rect 9950 11500 9956 11512
rect 10008 11500 10014 11552
rect 14277 11543 14335 11549
rect 14277 11509 14289 11543
rect 14323 11540 14335 11543
rect 14366 11540 14372 11552
rect 14323 11512 14372 11540
rect 14323 11509 14335 11512
rect 14277 11503 14335 11509
rect 14366 11500 14372 11512
rect 14424 11500 14430 11552
rect 17310 11500 17316 11552
rect 17368 11540 17374 11552
rect 17911 11543 17969 11549
rect 17911 11540 17923 11543
rect 17368 11512 17923 11540
rect 17368 11500 17374 11512
rect 17911 11509 17923 11512
rect 17957 11509 17969 11543
rect 17911 11503 17969 11509
rect 184 11450 18920 11472
rect 184 11398 3106 11450
rect 3158 11398 3170 11450
rect 3222 11398 3234 11450
rect 3286 11398 3298 11450
rect 3350 11398 3362 11450
rect 3414 11398 6206 11450
rect 6258 11398 6270 11450
rect 6322 11398 6334 11450
rect 6386 11398 6398 11450
rect 6450 11398 6462 11450
rect 6514 11398 9306 11450
rect 9358 11398 9370 11450
rect 9422 11398 9434 11450
rect 9486 11398 9498 11450
rect 9550 11398 9562 11450
rect 9614 11398 12406 11450
rect 12458 11398 12470 11450
rect 12522 11398 12534 11450
rect 12586 11398 12598 11450
rect 12650 11398 12662 11450
rect 12714 11398 15506 11450
rect 15558 11398 15570 11450
rect 15622 11398 15634 11450
rect 15686 11398 15698 11450
rect 15750 11398 15762 11450
rect 15814 11398 18606 11450
rect 18658 11398 18670 11450
rect 18722 11398 18734 11450
rect 18786 11398 18798 11450
rect 18850 11398 18862 11450
rect 18914 11398 18920 11450
rect 184 11376 18920 11398
rect 1949 11339 2007 11345
rect 1949 11305 1961 11339
rect 1995 11336 2007 11339
rect 2958 11336 2964 11348
rect 1995 11308 2964 11336
rect 1995 11305 2007 11308
rect 1949 11299 2007 11305
rect 2958 11296 2964 11308
rect 3016 11296 3022 11348
rect 6914 11336 6920 11348
rect 6875 11308 6920 11336
rect 6914 11296 6920 11308
rect 6972 11296 6978 11348
rect 8294 11336 8300 11348
rect 8255 11308 8300 11336
rect 8294 11296 8300 11308
rect 8352 11296 8358 11348
rect 10594 11296 10600 11348
rect 10652 11336 10658 11348
rect 10873 11339 10931 11345
rect 10873 11336 10885 11339
rect 10652 11308 10885 11336
rect 10652 11296 10658 11308
rect 10873 11305 10885 11308
rect 10919 11305 10931 11339
rect 10873 11299 10931 11305
rect 13725 11339 13783 11345
rect 13725 11305 13737 11339
rect 13771 11336 13783 11339
rect 14737 11339 14795 11345
rect 14737 11336 14749 11339
rect 13771 11308 14749 11336
rect 13771 11305 13783 11308
rect 13725 11299 13783 11305
rect 14737 11305 14749 11308
rect 14783 11305 14795 11339
rect 15194 11336 15200 11348
rect 15107 11308 15200 11336
rect 14737 11299 14795 11305
rect 15194 11296 15200 11308
rect 15252 11336 15258 11348
rect 16022 11336 16028 11348
rect 15252 11308 16028 11336
rect 15252 11296 15258 11308
rect 16022 11296 16028 11308
rect 16080 11296 16086 11348
rect 16117 11339 16175 11345
rect 16117 11305 16129 11339
rect 16163 11336 16175 11339
rect 16482 11336 16488 11348
rect 16163 11308 16488 11336
rect 16163 11305 16175 11308
rect 16117 11299 16175 11305
rect 16482 11296 16488 11308
rect 16540 11296 16546 11348
rect 16577 11339 16635 11345
rect 16577 11305 16589 11339
rect 16623 11336 16635 11339
rect 16666 11336 16672 11348
rect 16623 11308 16672 11336
rect 16623 11305 16635 11308
rect 16577 11299 16635 11305
rect 16666 11296 16672 11308
rect 16724 11296 16730 11348
rect 18046 11296 18052 11348
rect 18104 11336 18110 11348
rect 18233 11339 18291 11345
rect 18233 11336 18245 11339
rect 18104 11308 18245 11336
rect 18104 11296 18110 11308
rect 18233 11305 18245 11308
rect 18279 11305 18291 11339
rect 18233 11299 18291 11305
rect 1118 11268 1124 11280
rect 584 11240 1124 11268
rect 584 11209 612 11240
rect 1118 11228 1124 11240
rect 1176 11228 1182 11280
rect 5442 11268 5448 11280
rect 5403 11240 5448 11268
rect 5442 11228 5448 11240
rect 5500 11228 5506 11280
rect 6730 11268 6736 11280
rect 6670 11240 6736 11268
rect 6730 11228 6736 11240
rect 6788 11228 6794 11280
rect 9585 11271 9643 11277
rect 9585 11237 9597 11271
rect 9631 11268 9643 11271
rect 10318 11268 10324 11280
rect 9631 11240 10324 11268
rect 9631 11237 9643 11240
rect 9585 11231 9643 11237
rect 10318 11228 10324 11240
rect 10376 11228 10382 11280
rect 11606 11268 11612 11280
rect 11072 11240 11612 11268
rect 569 11203 627 11209
rect 569 11169 581 11203
rect 615 11169 627 11203
rect 569 11163 627 11169
rect 836 11203 894 11209
rect 836 11169 848 11203
rect 882 11200 894 11203
rect 2130 11200 2136 11212
rect 882 11172 2136 11200
rect 882 11169 894 11172
rect 836 11163 894 11169
rect 2130 11160 2136 11172
rect 2188 11160 2194 11212
rect 2774 11160 2780 11212
rect 2832 11200 2838 11212
rect 2961 11203 3019 11209
rect 2961 11200 2973 11203
rect 2832 11172 2973 11200
rect 2832 11160 2838 11172
rect 2961 11169 2973 11172
rect 3007 11169 3019 11203
rect 2961 11163 3019 11169
rect 4522 11160 4528 11212
rect 4580 11200 4586 11212
rect 11072 11209 11100 11240
rect 11606 11228 11612 11240
rect 11664 11228 11670 11280
rect 16393 11271 16451 11277
rect 13740 11240 15884 11268
rect 13740 11212 13768 11240
rect 5169 11203 5227 11209
rect 5169 11200 5181 11203
rect 4580 11172 5181 11200
rect 4580 11160 4586 11172
rect 5169 11169 5181 11172
rect 5215 11169 5227 11203
rect 5169 11163 5227 11169
rect 11057 11203 11115 11209
rect 11057 11169 11069 11203
rect 11103 11169 11115 11203
rect 11057 11163 11115 11169
rect 11149 11203 11207 11209
rect 11149 11169 11161 11203
rect 11195 11200 11207 11203
rect 11330 11200 11336 11212
rect 11195 11172 11336 11200
rect 11195 11169 11207 11172
rect 11149 11163 11207 11169
rect 11330 11160 11336 11172
rect 11388 11160 11394 11212
rect 11425 11203 11483 11209
rect 11425 11169 11437 11203
rect 11471 11200 11483 11203
rect 11790 11200 11796 11212
rect 11471 11172 11796 11200
rect 11471 11169 11483 11172
rect 11425 11163 11483 11169
rect 11790 11160 11796 11172
rect 11848 11160 11854 11212
rect 13722 11160 13728 11212
rect 13780 11160 13786 11212
rect 13817 11203 13875 11209
rect 13817 11169 13829 11203
rect 13863 11200 13875 11203
rect 13863 11172 14780 11200
rect 13863 11169 13875 11172
rect 13817 11163 13875 11169
rect 2869 11135 2927 11141
rect 2869 11101 2881 11135
rect 2915 11132 2927 11135
rect 10965 11135 11023 11141
rect 2915 11104 3004 11132
rect 2915 11101 2927 11104
rect 2869 11095 2927 11101
rect 2976 11076 3004 11104
rect 10965 11101 10977 11135
rect 11011 11101 11023 11135
rect 10965 11095 11023 11101
rect 11241 11135 11299 11141
rect 11241 11101 11253 11135
rect 11287 11132 11299 11135
rect 11698 11132 11704 11144
rect 11287 11104 11704 11132
rect 11287 11101 11299 11104
rect 11241 11095 11299 11101
rect 2958 11024 2964 11076
rect 3016 11024 3022 11076
rect 3329 11067 3387 11073
rect 3329 11033 3341 11067
rect 3375 11064 3387 11067
rect 3510 11064 3516 11076
rect 3375 11036 3516 11064
rect 3375 11033 3387 11036
rect 3329 11027 3387 11033
rect 3510 11024 3516 11036
rect 3568 11024 3574 11076
rect 10980 11064 11008 11095
rect 11698 11092 11704 11104
rect 11756 11092 11762 11144
rect 14001 11135 14059 11141
rect 14001 11101 14013 11135
rect 14047 11132 14059 11135
rect 14752 11132 14780 11172
rect 14826 11160 14832 11212
rect 14884 11200 14890 11212
rect 15856 11209 15884 11240
rect 16393 11237 16405 11271
rect 16439 11268 16451 11271
rect 16758 11268 16764 11280
rect 16439 11240 16764 11268
rect 16439 11237 16451 11240
rect 16393 11231 16451 11237
rect 16758 11228 16764 11240
rect 16816 11268 16822 11280
rect 17129 11271 17187 11277
rect 17129 11268 17141 11271
rect 16816 11240 17141 11268
rect 16816 11228 16822 11240
rect 17129 11237 17141 11240
rect 17175 11237 17187 11271
rect 17129 11231 17187 11237
rect 15105 11203 15163 11209
rect 15105 11200 15117 11203
rect 14884 11172 15117 11200
rect 14884 11160 14890 11172
rect 15105 11169 15117 11172
rect 15151 11169 15163 11203
rect 15105 11163 15163 11169
rect 15841 11203 15899 11209
rect 15841 11169 15853 11203
rect 15887 11200 15899 11203
rect 16669 11203 16727 11209
rect 16669 11200 16681 11203
rect 15887 11172 16681 11200
rect 15887 11169 15899 11172
rect 15841 11163 15899 11169
rect 16669 11169 16681 11172
rect 16715 11200 16727 11203
rect 17310 11200 17316 11212
rect 16715 11172 17316 11200
rect 16715 11169 16727 11172
rect 16669 11163 16727 11169
rect 17310 11160 17316 11172
rect 17368 11160 17374 11212
rect 17494 11200 17500 11212
rect 17455 11172 17500 11200
rect 17494 11160 17500 11172
rect 17552 11160 17558 11212
rect 17957 11203 18015 11209
rect 17957 11169 17969 11203
rect 18003 11200 18015 11203
rect 18414 11200 18420 11212
rect 18003 11172 18420 11200
rect 18003 11169 18015 11172
rect 17957 11163 18015 11169
rect 18414 11160 18420 11172
rect 18472 11160 18478 11212
rect 15194 11132 15200 11144
rect 14047 11104 14136 11132
rect 14752 11104 15200 11132
rect 14047 11101 14059 11104
rect 14001 11095 14059 11101
rect 12802 11064 12808 11076
rect 4540 11036 5304 11064
rect 10980 11036 12808 11064
rect 2222 10956 2228 11008
rect 2280 10996 2286 11008
rect 4540 10996 4568 11036
rect 2280 10968 4568 10996
rect 4617 10999 4675 11005
rect 2280 10956 2286 10968
rect 4617 10965 4629 10999
rect 4663 10996 4675 10999
rect 4982 10996 4988 11008
rect 4663 10968 4988 10996
rect 4663 10965 4675 10968
rect 4617 10959 4675 10965
rect 4982 10956 4988 10968
rect 5040 10956 5046 11008
rect 5276 10996 5304 11036
rect 12802 11024 12808 11036
rect 12860 11024 12866 11076
rect 5626 10996 5632 11008
rect 5276 10968 5632 10996
rect 5626 10956 5632 10968
rect 5684 10956 5690 11008
rect 12434 10956 12440 11008
rect 12492 10996 12498 11008
rect 13357 10999 13415 11005
rect 13357 10996 13369 10999
rect 12492 10968 13369 10996
rect 12492 10956 12498 10968
rect 13357 10965 13369 10968
rect 13403 10965 13415 10999
rect 13357 10959 13415 10965
rect 13446 10956 13452 11008
rect 13504 10996 13510 11008
rect 14108 10996 14136 11104
rect 15194 11092 15200 11104
rect 15252 11092 15258 11144
rect 15289 11135 15347 11141
rect 15289 11101 15301 11135
rect 15335 11101 15347 11135
rect 15289 11095 15347 11101
rect 16117 11135 16175 11141
rect 16117 11101 16129 11135
rect 16163 11101 16175 11135
rect 16117 11095 16175 11101
rect 15102 11024 15108 11076
rect 15160 11064 15166 11076
rect 15304 11064 15332 11095
rect 15930 11064 15936 11076
rect 15160 11036 15332 11064
rect 15891 11036 15936 11064
rect 15160 11024 15166 11036
rect 15930 11024 15936 11036
rect 15988 11024 15994 11076
rect 16132 11064 16160 11095
rect 16393 11067 16451 11073
rect 16393 11064 16405 11067
rect 16132 11036 16405 11064
rect 16393 11033 16405 11036
rect 16439 11033 16451 11067
rect 16393 11027 16451 11033
rect 16758 10996 16764 11008
rect 13504 10968 16764 10996
rect 13504 10956 13510 10968
rect 16758 10956 16764 10968
rect 16816 10956 16822 11008
rect 184 10906 18860 10928
rect 184 10854 1556 10906
rect 1608 10854 1620 10906
rect 1672 10854 1684 10906
rect 1736 10854 1748 10906
rect 1800 10854 1812 10906
rect 1864 10854 4656 10906
rect 4708 10854 4720 10906
rect 4772 10854 4784 10906
rect 4836 10854 4848 10906
rect 4900 10854 4912 10906
rect 4964 10854 7756 10906
rect 7808 10854 7820 10906
rect 7872 10854 7884 10906
rect 7936 10854 7948 10906
rect 8000 10854 8012 10906
rect 8064 10854 10856 10906
rect 10908 10854 10920 10906
rect 10972 10854 10984 10906
rect 11036 10854 11048 10906
rect 11100 10854 11112 10906
rect 11164 10854 13956 10906
rect 14008 10854 14020 10906
rect 14072 10854 14084 10906
rect 14136 10854 14148 10906
rect 14200 10854 14212 10906
rect 14264 10854 17056 10906
rect 17108 10854 17120 10906
rect 17172 10854 17184 10906
rect 17236 10854 17248 10906
rect 17300 10854 17312 10906
rect 17364 10854 18860 10906
rect 184 10832 18860 10854
rect 4338 10752 4344 10804
rect 4396 10792 4402 10804
rect 6546 10792 6552 10804
rect 4396 10764 6552 10792
rect 4396 10752 4402 10764
rect 6546 10752 6552 10764
rect 6604 10752 6610 10804
rect 12802 10752 12808 10804
rect 12860 10792 12866 10804
rect 12897 10795 12955 10801
rect 12897 10792 12909 10795
rect 12860 10764 12909 10792
rect 12860 10752 12866 10764
rect 12897 10761 12909 10764
rect 12943 10792 12955 10795
rect 13446 10792 13452 10804
rect 12943 10764 13452 10792
rect 12943 10761 12955 10764
rect 12897 10755 12955 10761
rect 13446 10752 13452 10764
rect 13504 10752 13510 10804
rect 15930 10752 15936 10804
rect 15988 10792 15994 10804
rect 16666 10792 16672 10804
rect 15988 10764 16672 10792
rect 15988 10752 15994 10764
rect 16666 10752 16672 10764
rect 16724 10752 16730 10804
rect 17494 10752 17500 10804
rect 17552 10792 17558 10804
rect 17678 10792 17684 10804
rect 17552 10764 17684 10792
rect 17552 10752 17558 10764
rect 17678 10752 17684 10764
rect 17736 10792 17742 10804
rect 17957 10795 18015 10801
rect 17957 10792 17969 10795
rect 17736 10764 17969 10792
rect 17736 10752 17742 10764
rect 17957 10761 17969 10764
rect 18003 10761 18015 10795
rect 17957 10755 18015 10761
rect 4154 10684 4160 10736
rect 4212 10724 4218 10736
rect 4709 10727 4767 10733
rect 4709 10724 4721 10727
rect 4212 10696 4721 10724
rect 4212 10684 4218 10696
rect 4709 10693 4721 10696
rect 4755 10693 4767 10727
rect 5258 10724 5264 10736
rect 5219 10696 5264 10724
rect 4709 10687 4767 10693
rect 5258 10684 5264 10696
rect 5316 10684 5322 10736
rect 14826 10724 14832 10736
rect 14787 10696 14832 10724
rect 14826 10684 14832 10696
rect 14884 10684 14890 10736
rect 4341 10659 4399 10665
rect 4341 10625 4353 10659
rect 4387 10656 4399 10659
rect 4387 10628 5028 10656
rect 4387 10625 4399 10628
rect 4341 10619 4399 10625
rect 1118 10588 1124 10600
rect 1079 10560 1124 10588
rect 1118 10548 1124 10560
rect 1176 10548 1182 10600
rect 1213 10591 1271 10597
rect 1213 10557 1225 10591
rect 1259 10588 1271 10591
rect 1581 10591 1639 10597
rect 1581 10588 1593 10591
rect 1259 10560 1593 10588
rect 1259 10557 1271 10560
rect 1213 10551 1271 10557
rect 1581 10557 1593 10560
rect 1627 10557 1639 10591
rect 1946 10588 1952 10600
rect 1907 10560 1952 10588
rect 1581 10551 1639 10557
rect 1946 10548 1952 10560
rect 2004 10548 2010 10600
rect 4062 10548 4068 10600
rect 4120 10588 4126 10600
rect 4433 10591 4491 10597
rect 4433 10588 4445 10591
rect 4120 10560 4445 10588
rect 4120 10548 4126 10560
rect 4433 10557 4445 10560
rect 4479 10557 4491 10591
rect 4433 10551 4491 10557
rect 4614 10548 4620 10600
rect 4672 10588 4678 10600
rect 4709 10591 4767 10597
rect 4709 10588 4721 10591
rect 4672 10560 4721 10588
rect 4672 10548 4678 10560
rect 4709 10557 4721 10560
rect 4755 10557 4767 10591
rect 4709 10551 4767 10557
rect 4893 10591 4951 10597
rect 4893 10557 4905 10591
rect 4939 10557 4951 10591
rect 4893 10551 4951 10557
rect 2314 10480 2320 10532
rect 2372 10480 2378 10532
rect 4157 10523 4215 10529
rect 4157 10489 4169 10523
rect 4203 10520 4215 10523
rect 4338 10520 4344 10532
rect 4203 10492 4344 10520
rect 4203 10489 4215 10492
rect 4157 10483 4215 10489
rect 4338 10480 4344 10492
rect 4396 10480 4402 10532
rect 4908 10520 4936 10551
rect 5000 10532 5028 10628
rect 14274 10616 14280 10668
rect 14332 10656 14338 10668
rect 14369 10659 14427 10665
rect 14369 10656 14381 10659
rect 14332 10628 14381 10656
rect 14332 10616 14338 10628
rect 14369 10625 14381 10628
rect 14415 10625 14427 10659
rect 14369 10619 14427 10625
rect 16114 10616 16120 10668
rect 16172 10656 16178 10668
rect 16209 10659 16267 10665
rect 16209 10656 16221 10659
rect 16172 10628 16221 10656
rect 16172 10616 16178 10628
rect 16209 10625 16221 10628
rect 16255 10625 16267 10659
rect 16209 10619 16267 10625
rect 10042 10548 10048 10600
rect 10100 10588 10106 10600
rect 10321 10591 10379 10597
rect 10321 10588 10333 10591
rect 10100 10560 10333 10588
rect 10100 10548 10106 10560
rect 10321 10557 10333 10560
rect 10367 10557 10379 10591
rect 10321 10551 10379 10557
rect 12434 10548 12440 10600
rect 12492 10588 12498 10600
rect 12989 10591 13047 10597
rect 12492 10560 12537 10588
rect 12492 10548 12498 10560
rect 12989 10557 13001 10591
rect 13035 10588 13047 10591
rect 13078 10588 13084 10600
rect 13035 10560 13084 10588
rect 13035 10557 13047 10560
rect 12989 10551 13047 10557
rect 13078 10548 13084 10560
rect 13136 10548 13142 10600
rect 14458 10588 14464 10600
rect 14419 10560 14464 10588
rect 14458 10548 14464 10560
rect 14516 10548 14522 10600
rect 4632 10492 4936 10520
rect 2774 10412 2780 10464
rect 2832 10452 2838 10464
rect 3375 10455 3433 10461
rect 3375 10452 3387 10455
rect 2832 10424 3387 10452
rect 2832 10412 2838 10424
rect 3375 10421 3387 10424
rect 3421 10421 3433 10455
rect 3375 10415 3433 10421
rect 4433 10455 4491 10461
rect 4433 10421 4445 10455
rect 4479 10452 4491 10455
rect 4632 10452 4660 10492
rect 4982 10480 4988 10532
rect 5040 10520 5046 10532
rect 6365 10523 6423 10529
rect 6365 10520 6377 10523
rect 5040 10492 6377 10520
rect 5040 10480 5046 10492
rect 6365 10489 6377 10492
rect 6411 10489 6423 10523
rect 6365 10483 6423 10489
rect 10502 10480 10508 10532
rect 10560 10520 10566 10532
rect 16482 10520 16488 10532
rect 10560 10492 12756 10520
rect 16443 10492 16488 10520
rect 10560 10480 10566 10492
rect 4479 10424 4660 10452
rect 4479 10421 4491 10424
rect 4433 10415 4491 10421
rect 10134 10412 10140 10464
rect 10192 10452 10198 10464
rect 10321 10455 10379 10461
rect 10321 10452 10333 10455
rect 10192 10424 10333 10452
rect 10192 10412 10198 10424
rect 10321 10421 10333 10424
rect 10367 10421 10379 10455
rect 10321 10415 10379 10421
rect 12250 10412 12256 10464
rect 12308 10452 12314 10464
rect 12728 10461 12756 10492
rect 16482 10480 16488 10492
rect 16540 10480 16546 10532
rect 16592 10492 16974 10520
rect 12529 10455 12587 10461
rect 12529 10452 12541 10455
rect 12308 10424 12541 10452
rect 12308 10412 12314 10424
rect 12529 10421 12541 10424
rect 12575 10421 12587 10455
rect 12529 10415 12587 10421
rect 12713 10455 12771 10461
rect 12713 10421 12725 10455
rect 12759 10421 12771 10455
rect 12713 10415 12771 10421
rect 16022 10412 16028 10464
rect 16080 10452 16086 10464
rect 16206 10452 16212 10464
rect 16080 10424 16212 10452
rect 16080 10412 16086 10424
rect 16206 10412 16212 10424
rect 16264 10452 16270 10464
rect 16592 10452 16620 10492
rect 16264 10424 16620 10452
rect 16264 10412 16270 10424
rect 184 10362 18920 10384
rect 184 10310 3106 10362
rect 3158 10310 3170 10362
rect 3222 10310 3234 10362
rect 3286 10310 3298 10362
rect 3350 10310 3362 10362
rect 3414 10310 6206 10362
rect 6258 10310 6270 10362
rect 6322 10310 6334 10362
rect 6386 10310 6398 10362
rect 6450 10310 6462 10362
rect 6514 10310 9306 10362
rect 9358 10310 9370 10362
rect 9422 10310 9434 10362
rect 9486 10310 9498 10362
rect 9550 10310 9562 10362
rect 9614 10310 12406 10362
rect 12458 10310 12470 10362
rect 12522 10310 12534 10362
rect 12586 10310 12598 10362
rect 12650 10310 12662 10362
rect 12714 10310 15506 10362
rect 15558 10310 15570 10362
rect 15622 10310 15634 10362
rect 15686 10310 15698 10362
rect 15750 10310 15762 10362
rect 15814 10310 18606 10362
rect 18658 10310 18670 10362
rect 18722 10310 18734 10362
rect 18786 10310 18798 10362
rect 18850 10310 18862 10362
rect 18914 10310 18920 10362
rect 184 10288 18920 10310
rect 1581 10251 1639 10257
rect 1581 10217 1593 10251
rect 1627 10248 1639 10251
rect 1946 10248 1952 10260
rect 1627 10220 1952 10248
rect 1627 10217 1639 10220
rect 1581 10211 1639 10217
rect 1946 10208 1952 10220
rect 2004 10208 2010 10260
rect 6457 10251 6515 10257
rect 6457 10217 6469 10251
rect 6503 10248 6515 10251
rect 6638 10248 6644 10260
rect 6503 10220 6644 10248
rect 6503 10217 6515 10220
rect 6457 10211 6515 10217
rect 6638 10208 6644 10220
rect 6696 10208 6702 10260
rect 7006 10208 7012 10260
rect 7064 10248 7070 10260
rect 7193 10251 7251 10257
rect 7193 10248 7205 10251
rect 7064 10220 7205 10248
rect 7064 10208 7070 10220
rect 7193 10217 7205 10220
rect 7239 10217 7251 10251
rect 7193 10211 7251 10217
rect 12250 10208 12256 10260
rect 12308 10248 12314 10260
rect 12437 10251 12495 10257
rect 12437 10248 12449 10251
rect 12308 10220 12449 10248
rect 12308 10208 12314 10220
rect 12437 10217 12449 10220
rect 12483 10217 12495 10251
rect 13078 10248 13084 10260
rect 13039 10220 13084 10248
rect 12437 10211 12495 10217
rect 13078 10208 13084 10220
rect 13136 10208 13142 10260
rect 16482 10208 16488 10260
rect 16540 10248 16546 10260
rect 17129 10251 17187 10257
rect 17129 10248 17141 10251
rect 16540 10220 17141 10248
rect 16540 10208 16546 10220
rect 17129 10217 17141 10220
rect 17175 10217 17187 10251
rect 17129 10211 17187 10217
rect 1118 10140 1124 10192
rect 1176 10180 1182 10192
rect 2777 10183 2835 10189
rect 2777 10180 2789 10183
rect 1176 10152 2789 10180
rect 1176 10140 1182 10152
rect 2777 10149 2789 10152
rect 2823 10149 2835 10183
rect 4522 10180 4528 10192
rect 4435 10152 4528 10180
rect 2777 10143 2835 10149
rect 4522 10140 4528 10152
rect 4580 10180 4586 10192
rect 5166 10180 5172 10192
rect 4580 10152 5172 10180
rect 4580 10140 4586 10152
rect 5166 10140 5172 10152
rect 5224 10140 5230 10192
rect 8478 10140 8484 10192
rect 8536 10140 8542 10192
rect 11422 10140 11428 10192
rect 11480 10140 11486 10192
rect 12894 10180 12900 10192
rect 12728 10152 12900 10180
rect 1949 10115 2007 10121
rect 1949 10081 1961 10115
rect 1995 10081 2007 10115
rect 1949 10075 2007 10081
rect 2041 10115 2099 10121
rect 2041 10081 2053 10115
rect 2087 10112 2099 10115
rect 2866 10112 2872 10124
rect 2087 10084 2872 10112
rect 2087 10081 2099 10084
rect 2041 10075 2099 10081
rect 1964 9976 1992 10075
rect 2866 10072 2872 10084
rect 2924 10072 2930 10124
rect 6365 10115 6423 10121
rect 6365 10081 6377 10115
rect 6411 10081 6423 10115
rect 6365 10075 6423 10081
rect 6549 10115 6607 10121
rect 6549 10081 6561 10115
rect 6595 10112 6607 10115
rect 7006 10112 7012 10124
rect 6595 10084 7012 10112
rect 6595 10081 6607 10084
rect 6549 10075 6607 10081
rect 2222 10044 2228 10056
rect 2183 10016 2228 10044
rect 2222 10004 2228 10016
rect 2280 10004 2286 10056
rect 6380 10044 6408 10075
rect 7006 10072 7012 10084
rect 7064 10072 7070 10124
rect 7558 10112 7564 10124
rect 7519 10084 7564 10112
rect 7558 10072 7564 10084
rect 7616 10072 7622 10124
rect 10134 10112 10140 10124
rect 10095 10084 10140 10112
rect 10134 10072 10140 10084
rect 10192 10072 10198 10124
rect 10502 10112 10508 10124
rect 10463 10084 10508 10112
rect 10502 10072 10508 10084
rect 10560 10072 10566 10124
rect 12728 10121 12756 10152
rect 12894 10140 12900 10152
rect 12952 10180 12958 10192
rect 12952 10152 13124 10180
rect 12952 10140 12958 10152
rect 12712 10115 12770 10121
rect 12712 10081 12724 10115
rect 12758 10081 12770 10115
rect 12712 10075 12770 10081
rect 12802 10072 12808 10124
rect 12860 10112 12866 10124
rect 13096 10121 13124 10152
rect 16942 10140 16948 10192
rect 17000 10180 17006 10192
rect 17000 10152 17494 10180
rect 17000 10140 17006 10152
rect 13081 10115 13139 10121
rect 12860 10084 12905 10112
rect 12860 10072 12866 10084
rect 13081 10081 13093 10115
rect 13127 10081 13139 10115
rect 13081 10075 13139 10081
rect 13265 10115 13323 10121
rect 13265 10081 13277 10115
rect 13311 10112 13323 10115
rect 14458 10112 14464 10124
rect 13311 10084 14464 10112
rect 13311 10081 13323 10084
rect 13265 10075 13323 10081
rect 6822 10044 6828 10056
rect 6380 10016 6828 10044
rect 6822 10004 6828 10016
rect 6880 10004 6886 10056
rect 7929 10047 7987 10053
rect 7929 10013 7941 10047
rect 7975 10044 7987 10047
rect 8294 10044 8300 10056
rect 7975 10016 8300 10044
rect 7975 10013 7987 10016
rect 7929 10007 7987 10013
rect 8294 10004 8300 10016
rect 8352 10004 8358 10056
rect 11931 10047 11989 10053
rect 11931 10013 11943 10047
rect 11977 10044 11989 10047
rect 13280 10044 13308 10075
rect 14458 10072 14464 10084
rect 14516 10072 14522 10124
rect 17310 10072 17316 10124
rect 17368 10121 17374 10124
rect 17466 10121 17494 10152
rect 17368 10115 17391 10121
rect 17379 10081 17391 10115
rect 17368 10075 17391 10081
rect 17451 10115 17509 10121
rect 17451 10081 17463 10115
rect 17497 10081 17509 10115
rect 17678 10112 17684 10124
rect 17639 10084 17684 10112
rect 17451 10075 17509 10081
rect 17368 10072 17374 10075
rect 17678 10072 17684 10084
rect 17736 10072 17742 10124
rect 11977 10016 13308 10044
rect 11977 10013 11989 10016
rect 11931 10007 11989 10013
rect 2774 9976 2780 9988
rect 1964 9948 2780 9976
rect 2774 9936 2780 9948
rect 2832 9936 2838 9988
rect 11330 9936 11336 9988
rect 11388 9976 11394 9988
rect 16574 9976 16580 9988
rect 11388 9948 16580 9976
rect 11388 9936 11394 9948
rect 16574 9936 16580 9948
rect 16632 9976 16638 9988
rect 17586 9976 17592 9988
rect 16632 9948 17592 9976
rect 16632 9936 16638 9948
rect 17586 9936 17592 9948
rect 17644 9936 17650 9988
rect 9030 9868 9036 9920
rect 9088 9908 9094 9920
rect 9355 9911 9413 9917
rect 9355 9908 9367 9911
rect 9088 9880 9367 9908
rect 9088 9868 9094 9880
rect 9355 9877 9367 9880
rect 9401 9877 9413 9911
rect 9355 9871 9413 9877
rect 12342 9868 12348 9920
rect 12400 9908 12406 9920
rect 16022 9908 16028 9920
rect 12400 9880 16028 9908
rect 12400 9868 12406 9880
rect 16022 9868 16028 9880
rect 16080 9868 16086 9920
rect 184 9818 18860 9840
rect 184 9766 1556 9818
rect 1608 9766 1620 9818
rect 1672 9766 1684 9818
rect 1736 9766 1748 9818
rect 1800 9766 1812 9818
rect 1864 9766 4656 9818
rect 4708 9766 4720 9818
rect 4772 9766 4784 9818
rect 4836 9766 4848 9818
rect 4900 9766 4912 9818
rect 4964 9766 7756 9818
rect 7808 9766 7820 9818
rect 7872 9766 7884 9818
rect 7936 9766 7948 9818
rect 8000 9766 8012 9818
rect 8064 9766 10856 9818
rect 10908 9766 10920 9818
rect 10972 9766 10984 9818
rect 11036 9766 11048 9818
rect 11100 9766 11112 9818
rect 11164 9766 13956 9818
rect 14008 9766 14020 9818
rect 14072 9766 14084 9818
rect 14136 9766 14148 9818
rect 14200 9766 14212 9818
rect 14264 9766 17056 9818
rect 17108 9766 17120 9818
rect 17172 9766 17184 9818
rect 17236 9766 17248 9818
rect 17300 9766 17312 9818
rect 17364 9766 18860 9818
rect 184 9744 18860 9766
rect 2866 9636 2872 9648
rect 2827 9608 2872 9636
rect 2866 9596 2872 9608
rect 2924 9596 2930 9648
rect 8294 9636 8300 9648
rect 8255 9608 8300 9636
rect 8294 9596 8300 9608
rect 8352 9596 8358 9648
rect 8757 9639 8815 9645
rect 8757 9636 8769 9639
rect 8404 9608 8769 9636
rect 3421 9571 3479 9577
rect 3421 9537 3433 9571
rect 3467 9568 3479 9571
rect 4246 9568 4252 9580
rect 3467 9540 4252 9568
rect 3467 9537 3479 9540
rect 3421 9531 3479 9537
rect 4246 9528 4252 9540
rect 4304 9528 4310 9580
rect 7006 9528 7012 9580
rect 7064 9568 7070 9580
rect 8404 9577 8432 9608
rect 8757 9605 8769 9608
rect 8803 9605 8815 9639
rect 8757 9599 8815 9605
rect 8389 9571 8447 9577
rect 7064 9540 8340 9568
rect 7064 9528 7070 9540
rect 2406 9460 2412 9512
rect 2464 9500 2470 9512
rect 2501 9503 2559 9509
rect 2501 9500 2513 9503
rect 2464 9472 2513 9500
rect 2464 9460 2470 9472
rect 2501 9469 2513 9472
rect 2547 9469 2559 9503
rect 2501 9463 2559 9469
rect 3237 9503 3295 9509
rect 3237 9469 3249 9503
rect 3283 9500 3295 9503
rect 3510 9500 3516 9512
rect 3283 9472 3516 9500
rect 3283 9469 3295 9472
rect 3237 9463 3295 9469
rect 3510 9460 3516 9472
rect 3568 9460 3574 9512
rect 5721 9503 5779 9509
rect 5721 9469 5733 9503
rect 5767 9500 5779 9503
rect 7558 9500 7564 9512
rect 5767 9472 7564 9500
rect 5767 9469 5779 9472
rect 5721 9463 5779 9469
rect 7558 9460 7564 9472
rect 7616 9460 7622 9512
rect 8128 9509 8156 9540
rect 8113 9503 8171 9509
rect 8113 9469 8125 9503
rect 8159 9469 8171 9503
rect 8113 9463 8171 9469
rect 8205 9503 8263 9509
rect 8205 9469 8217 9503
rect 8251 9469 8263 9503
rect 8312 9500 8340 9540
rect 8389 9537 8401 9571
rect 8435 9537 8447 9571
rect 8389 9531 8447 9537
rect 9030 9500 9036 9512
rect 8312 9472 9036 9500
rect 8205 9463 8263 9469
rect 2225 9435 2283 9441
rect 2225 9401 2237 9435
rect 2271 9432 2283 9435
rect 3329 9435 3387 9441
rect 2271 9404 2305 9432
rect 2271 9401 2283 9404
rect 2225 9395 2283 9401
rect 3329 9401 3341 9435
rect 3375 9432 3387 9435
rect 4154 9432 4160 9444
rect 3375 9404 4160 9432
rect 3375 9401 3387 9404
rect 3329 9395 3387 9401
rect 2130 9324 2136 9376
rect 2188 9364 2194 9376
rect 2240 9364 2268 9395
rect 4154 9392 4160 9404
rect 4212 9392 4218 9444
rect 2314 9364 2320 9376
rect 2188 9336 2320 9364
rect 2188 9324 2194 9336
rect 2314 9324 2320 9336
rect 2372 9324 2378 9376
rect 4801 9367 4859 9373
rect 4801 9333 4813 9367
rect 4847 9364 4859 9367
rect 4982 9364 4988 9376
rect 4847 9336 4988 9364
rect 4847 9333 4859 9336
rect 4801 9327 4859 9333
rect 4982 9324 4988 9336
rect 5040 9324 5046 9376
rect 5258 9324 5264 9376
rect 5316 9364 5322 9376
rect 5445 9367 5503 9373
rect 5445 9364 5457 9367
rect 5316 9336 5457 9364
rect 5316 9324 5322 9336
rect 5445 9333 5457 9336
rect 5491 9333 5503 9367
rect 8220 9364 8248 9463
rect 9030 9460 9036 9472
rect 9088 9460 9094 9512
rect 14274 9500 14280 9512
rect 14235 9472 14280 9500
rect 14274 9460 14280 9472
rect 14332 9460 14338 9512
rect 14642 9500 14648 9512
rect 14603 9472 14648 9500
rect 14642 9460 14648 9472
rect 14700 9460 14706 9512
rect 15013 9503 15071 9509
rect 15013 9469 15025 9503
rect 15059 9469 15071 9503
rect 15013 9463 15071 9469
rect 8294 9392 8300 9444
rect 8352 9432 8358 9444
rect 8757 9435 8815 9441
rect 8757 9432 8769 9435
rect 8352 9404 8769 9432
rect 8352 9392 8358 9404
rect 8757 9401 8769 9404
rect 8803 9401 8815 9435
rect 8757 9395 8815 9401
rect 14458 9392 14464 9444
rect 14516 9432 14522 9444
rect 15028 9432 15056 9463
rect 14516 9404 15056 9432
rect 14516 9392 14522 9404
rect 8941 9367 8999 9373
rect 8941 9364 8953 9367
rect 8220 9336 8953 9364
rect 5445 9327 5503 9333
rect 8941 9333 8953 9336
rect 8987 9364 8999 9367
rect 9030 9364 9036 9376
rect 8987 9336 9036 9364
rect 8987 9333 8999 9336
rect 8941 9327 8999 9333
rect 9030 9324 9036 9336
rect 9088 9324 9094 9376
rect 11422 9324 11428 9376
rect 11480 9364 11486 9376
rect 11790 9364 11796 9376
rect 11480 9336 11796 9364
rect 11480 9324 11486 9336
rect 11790 9324 11796 9336
rect 11848 9364 11854 9376
rect 12069 9367 12127 9373
rect 12069 9364 12081 9367
rect 11848 9336 12081 9364
rect 11848 9324 11854 9336
rect 12069 9333 12081 9336
rect 12115 9364 12127 9367
rect 12342 9364 12348 9376
rect 12115 9336 12348 9364
rect 12115 9333 12127 9336
rect 12069 9327 12127 9333
rect 12342 9324 12348 9336
rect 12400 9364 12406 9376
rect 12437 9367 12495 9373
rect 12437 9364 12449 9367
rect 12400 9336 12449 9364
rect 12400 9324 12406 9336
rect 12437 9333 12449 9336
rect 12483 9333 12495 9367
rect 12437 9327 12495 9333
rect 15013 9367 15071 9373
rect 15013 9333 15025 9367
rect 15059 9364 15071 9367
rect 15102 9364 15108 9376
rect 15059 9336 15108 9364
rect 15059 9333 15071 9336
rect 15013 9327 15071 9333
rect 15102 9324 15108 9336
rect 15160 9324 15166 9376
rect 184 9274 18920 9296
rect 184 9222 3106 9274
rect 3158 9222 3170 9274
rect 3222 9222 3234 9274
rect 3286 9222 3298 9274
rect 3350 9222 3362 9274
rect 3414 9222 6206 9274
rect 6258 9222 6270 9274
rect 6322 9222 6334 9274
rect 6386 9222 6398 9274
rect 6450 9222 6462 9274
rect 6514 9222 9306 9274
rect 9358 9222 9370 9274
rect 9422 9222 9434 9274
rect 9486 9222 9498 9274
rect 9550 9222 9562 9274
rect 9614 9222 12406 9274
rect 12458 9222 12470 9274
rect 12522 9222 12534 9274
rect 12586 9222 12598 9274
rect 12650 9222 12662 9274
rect 12714 9222 15506 9274
rect 15558 9222 15570 9274
rect 15622 9222 15634 9274
rect 15686 9222 15698 9274
rect 15750 9222 15762 9274
rect 15814 9222 18606 9274
rect 18658 9222 18670 9274
rect 18722 9222 18734 9274
rect 18786 9222 18798 9274
rect 18850 9222 18862 9274
rect 18914 9222 18920 9274
rect 184 9200 18920 9222
rect 1765 9163 1823 9169
rect 1765 9129 1777 9163
rect 1811 9160 1823 9163
rect 3145 9163 3203 9169
rect 3145 9160 3157 9163
rect 1811 9132 3157 9160
rect 1811 9129 1823 9132
rect 1765 9123 1823 9129
rect 3145 9129 3157 9132
rect 3191 9129 3203 9163
rect 3145 9123 3203 9129
rect 3605 9163 3663 9169
rect 3605 9129 3617 9163
rect 3651 9160 3663 9163
rect 4157 9163 4215 9169
rect 4157 9160 4169 9163
rect 3651 9132 4169 9160
rect 3651 9129 3663 9132
rect 3605 9123 3663 9129
rect 4157 9129 4169 9132
rect 4203 9160 4215 9163
rect 4430 9160 4436 9172
rect 4203 9132 4436 9160
rect 4203 9129 4215 9132
rect 4157 9123 4215 9129
rect 4430 9120 4436 9132
rect 4488 9120 4494 9172
rect 5626 9120 5632 9172
rect 5684 9160 5690 9172
rect 5684 9132 6775 9160
rect 5684 9120 5690 9132
rect 6747 9092 6775 9132
rect 14642 9120 14648 9172
rect 14700 9160 14706 9172
rect 17313 9163 17371 9169
rect 14700 9132 15516 9160
rect 14700 9120 14706 9132
rect 8478 9092 8484 9104
rect 6670 9064 8484 9092
rect 8478 9052 8484 9064
rect 8536 9052 8542 9104
rect 11790 9092 11796 9104
rect 11730 9064 11796 9092
rect 11790 9052 11796 9064
rect 11848 9052 11854 9104
rect 12894 9092 12900 9104
rect 12544 9064 12900 9092
rect 1673 9027 1731 9033
rect 1673 8993 1685 9027
rect 1719 9024 1731 9027
rect 2314 9024 2320 9036
rect 1719 8996 2320 9024
rect 1719 8993 1731 8996
rect 1673 8987 1731 8993
rect 2314 8984 2320 8996
rect 2372 8984 2378 9036
rect 3513 9027 3571 9033
rect 3513 8993 3525 9027
rect 3559 9024 3571 9027
rect 3970 9024 3976 9036
rect 3559 8996 3976 9024
rect 3559 8993 3571 8996
rect 3513 8987 3571 8993
rect 3970 8984 3976 8996
rect 4028 8984 4034 9036
rect 4338 9024 4344 9036
rect 4251 8996 4344 9024
rect 4338 8984 4344 8996
rect 4396 9024 4402 9036
rect 5074 9024 5080 9036
rect 4396 8996 5080 9024
rect 4396 8984 4402 8996
rect 5074 8984 5080 8996
rect 5132 8984 5138 9036
rect 5258 9024 5264 9036
rect 5219 8996 5264 9024
rect 5258 8984 5264 8996
rect 5316 8984 5322 9036
rect 12544 9033 12572 9064
rect 12894 9052 12900 9064
rect 12952 9052 12958 9104
rect 14093 9095 14151 9101
rect 14093 9061 14105 9095
rect 14139 9092 14151 9095
rect 14458 9092 14464 9104
rect 14139 9064 14464 9092
rect 14139 9061 14151 9064
rect 14093 9055 14151 9061
rect 14458 9052 14464 9064
rect 14516 9052 14522 9104
rect 15381 9095 15439 9101
rect 15381 9061 15393 9095
rect 15427 9061 15439 9095
rect 15381 9055 15439 9061
rect 12529 9027 12587 9033
rect 12529 8993 12541 9027
rect 12575 8993 12587 9027
rect 12529 8987 12587 8993
rect 12621 9027 12679 9033
rect 12621 8993 12633 9027
rect 12667 8993 12679 9027
rect 12621 8987 12679 8993
rect 12713 9027 12771 9033
rect 12713 8993 12725 9027
rect 12759 9024 12771 9027
rect 12802 9024 12808 9036
rect 12759 8996 12808 9024
rect 12759 8993 12771 8996
rect 12713 8987 12771 8993
rect 1949 8959 2007 8965
rect 1949 8925 1961 8959
rect 1995 8956 2007 8959
rect 2222 8956 2228 8968
rect 1995 8928 2228 8956
rect 1995 8925 2007 8928
rect 1949 8919 2007 8925
rect 2222 8916 2228 8928
rect 2280 8956 2286 8968
rect 2406 8956 2412 8968
rect 2280 8928 2412 8956
rect 2280 8916 2286 8928
rect 2406 8916 2412 8928
rect 2464 8916 2470 8968
rect 3789 8959 3847 8965
rect 3789 8925 3801 8959
rect 3835 8956 3847 8959
rect 4246 8956 4252 8968
rect 3835 8928 4252 8956
rect 3835 8925 3847 8928
rect 3789 8919 3847 8925
rect 4246 8916 4252 8928
rect 4304 8916 4310 8968
rect 4617 8959 4675 8965
rect 4617 8925 4629 8959
rect 4663 8956 4675 8959
rect 4982 8956 4988 8968
rect 4663 8928 4988 8956
rect 4663 8925 4675 8928
rect 4617 8919 4675 8925
rect 4982 8916 4988 8928
rect 5040 8916 5046 8968
rect 5626 8956 5632 8968
rect 5587 8928 5632 8956
rect 5626 8916 5632 8928
rect 5684 8916 5690 8968
rect 10229 8959 10287 8965
rect 10229 8925 10241 8959
rect 10275 8925 10287 8959
rect 10229 8919 10287 8925
rect 10505 8959 10563 8965
rect 10505 8925 10517 8959
rect 10551 8956 10563 8959
rect 11238 8956 11244 8968
rect 10551 8928 11244 8956
rect 10551 8925 10563 8928
rect 10505 8919 10563 8925
rect 4264 8888 4292 8916
rect 4264 8860 5304 8888
rect 842 8780 848 8832
rect 900 8820 906 8832
rect 1305 8823 1363 8829
rect 1305 8820 1317 8823
rect 900 8792 1317 8820
rect 900 8780 906 8792
rect 1305 8789 1317 8792
rect 1351 8789 1363 8823
rect 1305 8783 1363 8789
rect 4525 8823 4583 8829
rect 4525 8789 4537 8823
rect 4571 8820 4583 8823
rect 5166 8820 5172 8832
rect 4571 8792 5172 8820
rect 4571 8789 4583 8792
rect 4525 8783 4583 8789
rect 5166 8780 5172 8792
rect 5224 8780 5230 8832
rect 5276 8820 5304 8860
rect 5902 8820 5908 8832
rect 5276 8792 5908 8820
rect 5902 8780 5908 8792
rect 5960 8780 5966 8832
rect 6822 8780 6828 8832
rect 6880 8820 6886 8832
rect 7055 8823 7113 8829
rect 7055 8820 7067 8823
rect 6880 8792 7067 8820
rect 6880 8780 6886 8792
rect 7055 8789 7067 8792
rect 7101 8789 7113 8823
rect 7055 8783 7113 8789
rect 10042 8780 10048 8832
rect 10100 8820 10106 8832
rect 10244 8820 10272 8919
rect 11238 8916 11244 8928
rect 11296 8916 11302 8968
rect 11977 8959 12035 8965
rect 11977 8925 11989 8959
rect 12023 8956 12035 8959
rect 12636 8956 12664 8987
rect 12802 8984 12808 8996
rect 12860 9024 12866 9036
rect 13722 9024 13728 9036
rect 12860 8996 13728 9024
rect 12860 8984 12866 8996
rect 13722 8984 13728 8996
rect 13780 8984 13786 9036
rect 14369 9027 14427 9033
rect 14369 9024 14381 9027
rect 13924 8996 14381 9024
rect 13924 8956 13952 8996
rect 14369 8993 14381 8996
rect 14415 9024 14427 9027
rect 14642 9024 14648 9036
rect 14415 8996 14648 9024
rect 14415 8993 14427 8996
rect 14369 8987 14427 8993
rect 14642 8984 14648 8996
rect 14700 8984 14706 9036
rect 14737 9027 14795 9033
rect 14737 8993 14749 9027
rect 14783 8993 14795 9027
rect 14737 8987 14795 8993
rect 14891 9027 14949 9033
rect 14891 8993 14903 9027
rect 14937 9024 14949 9027
rect 15396 9024 15424 9055
rect 14937 8996 15424 9024
rect 14937 8993 14949 8996
rect 14891 8987 14949 8993
rect 12023 8928 13952 8956
rect 12023 8925 12035 8928
rect 11977 8919 12035 8925
rect 12802 8888 12808 8900
rect 11532 8860 12808 8888
rect 11532 8820 11560 8860
rect 12802 8848 12808 8860
rect 12860 8848 12866 8900
rect 14274 8888 14280 8900
rect 14235 8860 14280 8888
rect 14274 8848 14280 8860
rect 14332 8848 14338 8900
rect 14369 8891 14427 8897
rect 14369 8857 14381 8891
rect 14415 8888 14427 8891
rect 14752 8888 14780 8987
rect 15381 8959 15439 8965
rect 15381 8925 15393 8959
rect 15427 8956 15439 8959
rect 15488 8956 15516 9132
rect 17313 9129 17325 9163
rect 17359 9160 17371 9163
rect 17402 9160 17408 9172
rect 17359 9132 17408 9160
rect 17359 9129 17371 9132
rect 17313 9123 17371 9129
rect 17402 9120 17408 9132
rect 17460 9120 17466 9172
rect 18230 9160 18236 9172
rect 18191 9132 18236 9160
rect 18230 9120 18236 9132
rect 18288 9120 18294 9172
rect 17221 9095 17279 9101
rect 17221 9061 17233 9095
rect 17267 9092 17279 9095
rect 17494 9092 17500 9104
rect 17267 9064 17500 9092
rect 17267 9061 17279 9064
rect 17221 9055 17279 9061
rect 17494 9052 17500 9064
rect 17552 9052 17558 9104
rect 15657 9027 15715 9033
rect 15657 8993 15669 9027
rect 15703 8993 15715 9027
rect 15657 8987 15715 8993
rect 15427 8928 15516 8956
rect 15427 8925 15439 8928
rect 15381 8919 15439 8925
rect 15102 8888 15108 8900
rect 14415 8860 14780 8888
rect 15063 8860 15108 8888
rect 14415 8857 14427 8860
rect 14369 8851 14427 8857
rect 15102 8848 15108 8860
rect 15160 8848 15166 8900
rect 15672 8888 15700 8987
rect 16298 8984 16304 9036
rect 16356 9024 16362 9036
rect 17129 9027 17187 9033
rect 17129 9024 17141 9027
rect 16356 8996 17141 9024
rect 16356 8984 16362 8996
rect 17129 8993 17141 8996
rect 17175 8993 17187 9027
rect 17129 8987 17187 8993
rect 17405 9027 17463 9033
rect 17405 8993 17417 9027
rect 17451 9024 17463 9027
rect 17954 9024 17960 9036
rect 17451 8996 17960 9024
rect 17451 8993 17463 8996
rect 17405 8987 17463 8993
rect 17954 8984 17960 8996
rect 18012 8984 18018 9036
rect 18414 9024 18420 9036
rect 18375 8996 18420 9024
rect 18414 8984 18420 8996
rect 18472 8984 18478 9036
rect 15488 8860 15700 8888
rect 17957 8891 18015 8897
rect 10100 8792 11560 8820
rect 10100 8780 10106 8792
rect 12066 8780 12072 8832
rect 12124 8820 12130 8832
rect 12345 8823 12403 8829
rect 12345 8820 12357 8823
rect 12124 8792 12357 8820
rect 12124 8780 12130 8792
rect 12345 8789 12357 8792
rect 12391 8789 12403 8823
rect 12345 8783 12403 8789
rect 14458 8780 14464 8832
rect 14516 8820 14522 8832
rect 15488 8820 15516 8860
rect 17957 8857 17969 8891
rect 18003 8888 18015 8891
rect 18414 8888 18420 8900
rect 18003 8860 18420 8888
rect 18003 8857 18015 8860
rect 17957 8851 18015 8857
rect 18414 8848 18420 8860
rect 18472 8848 18478 8900
rect 14516 8792 15516 8820
rect 14516 8780 14522 8792
rect 15562 8780 15568 8832
rect 15620 8820 15626 8832
rect 15620 8792 15665 8820
rect 15620 8780 15626 8792
rect 184 8730 18860 8752
rect 184 8678 1556 8730
rect 1608 8678 1620 8730
rect 1672 8678 1684 8730
rect 1736 8678 1748 8730
rect 1800 8678 1812 8730
rect 1864 8678 4656 8730
rect 4708 8678 4720 8730
rect 4772 8678 4784 8730
rect 4836 8678 4848 8730
rect 4900 8678 4912 8730
rect 4964 8678 7756 8730
rect 7808 8678 7820 8730
rect 7872 8678 7884 8730
rect 7936 8678 7948 8730
rect 8000 8678 8012 8730
rect 8064 8678 10856 8730
rect 10908 8678 10920 8730
rect 10972 8678 10984 8730
rect 11036 8678 11048 8730
rect 11100 8678 11112 8730
rect 11164 8678 13956 8730
rect 14008 8678 14020 8730
rect 14072 8678 14084 8730
rect 14136 8678 14148 8730
rect 14200 8678 14212 8730
rect 14264 8678 17056 8730
rect 17108 8678 17120 8730
rect 17172 8678 17184 8730
rect 17236 8678 17248 8730
rect 17300 8678 17312 8730
rect 17364 8678 18860 8730
rect 184 8656 18860 8678
rect 2958 8576 2964 8628
rect 3016 8616 3022 8628
rect 3053 8619 3111 8625
rect 3053 8616 3065 8619
rect 3016 8588 3065 8616
rect 3016 8576 3022 8588
rect 3053 8585 3065 8588
rect 3099 8585 3111 8619
rect 3970 8616 3976 8628
rect 3931 8588 3976 8616
rect 3053 8579 3111 8585
rect 3970 8576 3976 8588
rect 4028 8576 4034 8628
rect 4985 8619 5043 8625
rect 4985 8585 4997 8619
rect 5031 8616 5043 8619
rect 5166 8616 5172 8628
rect 5031 8588 5172 8616
rect 5031 8585 5043 8588
rect 4985 8579 5043 8585
rect 5166 8576 5172 8588
rect 5224 8576 5230 8628
rect 5353 8619 5411 8625
rect 5353 8585 5365 8619
rect 5399 8616 5411 8619
rect 5626 8616 5632 8628
rect 5399 8588 5632 8616
rect 5399 8585 5411 8588
rect 5353 8579 5411 8585
rect 5626 8576 5632 8588
rect 5684 8576 5690 8628
rect 11238 8616 11244 8628
rect 11199 8588 11244 8616
rect 11238 8576 11244 8588
rect 11296 8576 11302 8628
rect 14274 8576 14280 8628
rect 14332 8616 14338 8628
rect 15562 8616 15568 8628
rect 14332 8588 15568 8616
rect 14332 8576 14338 8588
rect 15562 8576 15568 8588
rect 15620 8576 15626 8628
rect 17954 8616 17960 8628
rect 17915 8588 17960 8616
rect 17954 8576 17960 8588
rect 18012 8576 18018 8628
rect 13541 8551 13599 8557
rect 13541 8517 13553 8551
rect 13587 8517 13599 8551
rect 14550 8548 14556 8560
rect 14511 8520 14556 8548
rect 13541 8511 13599 8517
rect 2774 8440 2780 8492
rect 2832 8480 2838 8492
rect 2961 8483 3019 8489
rect 2961 8480 2973 8483
rect 2832 8452 2973 8480
rect 2832 8440 2838 8452
rect 2961 8449 2973 8452
rect 3007 8480 3019 8483
rect 3970 8480 3976 8492
rect 3007 8452 3976 8480
rect 3007 8449 3019 8452
rect 2961 8443 3019 8449
rect 3970 8440 3976 8452
rect 4028 8440 4034 8492
rect 11149 8483 11207 8489
rect 11149 8449 11161 8483
rect 11195 8480 11207 8483
rect 12066 8480 12072 8492
rect 11195 8452 12072 8480
rect 11195 8449 11207 8452
rect 11149 8443 11207 8449
rect 12066 8440 12072 8452
rect 12124 8440 12130 8492
rect 3237 8415 3295 8421
rect 3237 8381 3249 8415
rect 3283 8381 3295 8415
rect 3237 8375 3295 8381
rect 3421 8415 3479 8421
rect 3421 8381 3433 8415
rect 3467 8412 3479 8415
rect 4157 8415 4215 8421
rect 4157 8412 4169 8415
rect 3467 8384 4169 8412
rect 3467 8381 3479 8384
rect 3421 8375 3479 8381
rect 4157 8381 4169 8384
rect 4203 8381 4215 8415
rect 4430 8412 4436 8424
rect 4391 8384 4436 8412
rect 4157 8375 4215 8381
rect 2314 8304 2320 8356
rect 2372 8344 2378 8356
rect 3252 8344 3280 8375
rect 4430 8372 4436 8384
rect 4488 8372 4494 8424
rect 5258 8412 5264 8424
rect 5219 8384 5264 8412
rect 5258 8372 5264 8384
rect 5316 8372 5322 8424
rect 5445 8415 5503 8421
rect 5445 8381 5457 8415
rect 5491 8412 5503 8415
rect 5626 8412 5632 8424
rect 5491 8384 5632 8412
rect 5491 8381 5503 8384
rect 5445 8375 5503 8381
rect 5626 8372 5632 8384
rect 5684 8372 5690 8424
rect 6822 8412 6828 8424
rect 6783 8384 6828 8412
rect 6822 8372 6828 8384
rect 6880 8372 6886 8424
rect 11330 8412 11336 8424
rect 11291 8384 11336 8412
rect 11330 8372 11336 8384
rect 11388 8372 11394 8424
rect 11425 8415 11483 8421
rect 11425 8381 11437 8415
rect 11471 8412 11483 8415
rect 12345 8415 12403 8421
rect 12345 8412 12357 8415
rect 11471 8384 12357 8412
rect 11471 8381 11483 8384
rect 11425 8375 11483 8381
rect 12345 8381 12357 8384
rect 12391 8381 12403 8415
rect 12345 8375 12403 8381
rect 12437 8415 12495 8421
rect 12437 8381 12449 8415
rect 12483 8412 12495 8415
rect 13556 8412 13584 8511
rect 14550 8508 14556 8520
rect 14608 8508 14614 8560
rect 16298 8548 16304 8560
rect 16259 8520 16304 8548
rect 16298 8508 16304 8520
rect 16356 8508 16362 8560
rect 13722 8440 13728 8492
rect 13780 8480 13786 8492
rect 14093 8483 14151 8489
rect 14093 8480 14105 8483
rect 13780 8452 14105 8480
rect 13780 8440 13786 8452
rect 14093 8449 14105 8452
rect 14139 8449 14151 8483
rect 14093 8443 14151 8449
rect 12483 8384 13584 8412
rect 14001 8415 14059 8421
rect 12483 8381 12495 8384
rect 12437 8375 12495 8381
rect 14001 8381 14013 8415
rect 14047 8412 14059 8415
rect 14568 8412 14596 8508
rect 16206 8480 16212 8492
rect 15948 8452 16212 8480
rect 15948 8421 15976 8452
rect 16206 8440 16212 8452
rect 16264 8480 16270 8492
rect 16264 8452 16712 8480
rect 16264 8440 16270 8452
rect 14047 8384 14596 8412
rect 15933 8415 15991 8421
rect 14047 8381 14059 8384
rect 14001 8375 14059 8381
rect 15933 8381 15945 8415
rect 15979 8381 15991 8415
rect 15933 8375 15991 8381
rect 16087 8415 16145 8421
rect 16087 8381 16099 8415
rect 16133 8412 16145 8415
rect 16133 8384 16344 8412
rect 16133 8381 16145 8384
rect 16087 8375 16145 8381
rect 2372 8316 3280 8344
rect 2372 8304 2378 8316
rect 5810 8304 5816 8356
rect 5868 8344 5874 8356
rect 6365 8347 6423 8353
rect 6365 8344 6377 8347
rect 5868 8316 6377 8344
rect 5868 8304 5874 8316
rect 6365 8313 6377 8316
rect 6411 8313 6423 8347
rect 6365 8307 6423 8313
rect 15286 8304 15292 8356
rect 15344 8344 15350 8356
rect 16316 8344 16344 8384
rect 16390 8372 16396 8424
rect 16448 8412 16454 8424
rect 16577 8415 16635 8421
rect 16577 8412 16589 8415
rect 16448 8384 16589 8412
rect 16448 8372 16454 8384
rect 16577 8381 16589 8384
rect 16623 8381 16635 8415
rect 16684 8412 16712 8452
rect 17218 8412 17224 8424
rect 16684 8384 17224 8412
rect 16577 8375 16635 8381
rect 17218 8372 17224 8384
rect 17276 8372 17282 8424
rect 16666 8344 16672 8356
rect 15344 8316 16252 8344
rect 16316 8316 16672 8344
rect 15344 8304 15350 8316
rect 4338 8276 4344 8288
rect 4299 8248 4344 8276
rect 4338 8236 4344 8248
rect 4396 8236 4402 8288
rect 13906 8276 13912 8288
rect 13867 8248 13912 8276
rect 13906 8236 13912 8248
rect 13964 8236 13970 8288
rect 16224 8276 16252 8316
rect 16666 8304 16672 8316
rect 16724 8304 16730 8356
rect 16833 8347 16891 8353
rect 16833 8344 16845 8347
rect 16776 8316 16845 8344
rect 16776 8276 16804 8316
rect 16833 8313 16845 8316
rect 16879 8313 16891 8347
rect 16833 8307 16891 8313
rect 16224 8248 16804 8276
rect 184 8186 18920 8208
rect 184 8134 3106 8186
rect 3158 8134 3170 8186
rect 3222 8134 3234 8186
rect 3286 8134 3298 8186
rect 3350 8134 3362 8186
rect 3414 8134 6206 8186
rect 6258 8134 6270 8186
rect 6322 8134 6334 8186
rect 6386 8134 6398 8186
rect 6450 8134 6462 8186
rect 6514 8134 9306 8186
rect 9358 8134 9370 8186
rect 9422 8134 9434 8186
rect 9486 8134 9498 8186
rect 9550 8134 9562 8186
rect 9614 8134 12406 8186
rect 12458 8134 12470 8186
rect 12522 8134 12534 8186
rect 12586 8134 12598 8186
rect 12650 8134 12662 8186
rect 12714 8134 15506 8186
rect 15558 8134 15570 8186
rect 15622 8134 15634 8186
rect 15686 8134 15698 8186
rect 15750 8134 15762 8186
rect 15814 8134 18606 8186
rect 18658 8134 18670 8186
rect 18722 8134 18734 8186
rect 18786 8134 18798 8186
rect 18850 8134 18862 8186
rect 18914 8134 18920 8186
rect 184 8112 18920 8134
rect 584 8044 2774 8072
rect 584 7948 612 8044
rect 842 8004 848 8016
rect 803 7976 848 8004
rect 842 7964 848 7976
rect 900 7964 906 8016
rect 2130 8004 2136 8016
rect 2070 7976 2136 8004
rect 2130 7964 2136 7976
rect 2188 7964 2194 8016
rect 566 7936 572 7948
rect 479 7908 572 7936
rect 566 7896 572 7908
rect 624 7896 630 7948
rect 2746 7936 2774 8044
rect 5258 8032 5264 8084
rect 5316 8072 5322 8084
rect 5353 8075 5411 8081
rect 5353 8072 5365 8075
rect 5316 8044 5365 8072
rect 5316 8032 5322 8044
rect 5353 8041 5365 8044
rect 5399 8041 5411 8075
rect 5353 8035 5411 8041
rect 13906 8032 13912 8084
rect 13964 8072 13970 8084
rect 14737 8075 14795 8081
rect 14737 8072 14749 8075
rect 13964 8044 14749 8072
rect 13964 8032 13970 8044
rect 14737 8041 14749 8044
rect 14783 8041 14795 8075
rect 15102 8072 15108 8084
rect 15063 8044 15108 8072
rect 14737 8035 14795 8041
rect 15102 8032 15108 8044
rect 15160 8032 15166 8084
rect 17494 8072 17500 8084
rect 17455 8044 17500 8072
rect 17494 8032 17500 8044
rect 17552 8032 17558 8084
rect 4522 8004 4528 8016
rect 4483 7976 4528 8004
rect 4522 7964 4528 7976
rect 4580 7964 4586 8016
rect 8478 7964 8484 8016
rect 8536 7964 8542 8016
rect 11238 8004 11244 8016
rect 10704 7976 11244 8004
rect 2961 7939 3019 7945
rect 2961 7936 2973 7939
rect 2746 7908 2973 7936
rect 2961 7905 2973 7908
rect 3007 7936 3019 7939
rect 7558 7936 7564 7948
rect 3007 7908 7564 7936
rect 3007 7905 3019 7908
rect 2961 7899 3019 7905
rect 7558 7896 7564 7908
rect 7616 7896 7622 7948
rect 10704 7945 10732 7976
rect 11238 7964 11244 7976
rect 11296 7964 11302 8016
rect 12802 8004 12808 8016
rect 12763 7976 12808 8004
rect 12802 7964 12808 7976
rect 12860 7964 12866 8016
rect 14366 8004 14372 8016
rect 14327 7976 14372 8004
rect 14366 7964 14372 7976
rect 14424 7964 14430 8016
rect 14550 7964 14556 8016
rect 14608 8004 14614 8016
rect 15197 8007 15255 8013
rect 15197 8004 15209 8007
rect 14608 7976 15209 8004
rect 14608 7964 14614 7976
rect 15197 7973 15209 7976
rect 15243 8004 15255 8007
rect 15749 8007 15807 8013
rect 15749 8004 15761 8007
rect 15243 7976 15761 8004
rect 15243 7973 15255 7976
rect 15197 7967 15255 7973
rect 15749 7973 15761 7976
rect 15795 7973 15807 8007
rect 15749 7967 15807 7973
rect 10689 7939 10747 7945
rect 10689 7905 10701 7939
rect 10735 7905 10747 7939
rect 10689 7899 10747 7905
rect 10778 7896 10784 7948
rect 10836 7936 10842 7948
rect 10965 7939 11023 7945
rect 10836 7908 10881 7936
rect 10836 7896 10842 7908
rect 10965 7905 10977 7939
rect 11011 7936 11023 7939
rect 12434 7936 12440 7948
rect 11011 7908 12440 7936
rect 11011 7905 11023 7908
rect 10965 7899 11023 7905
rect 12434 7896 12440 7908
rect 12492 7936 12498 7948
rect 13722 7936 13728 7948
rect 12492 7908 13728 7936
rect 12492 7896 12498 7908
rect 13722 7896 13728 7908
rect 13780 7896 13786 7948
rect 16666 7896 16672 7948
rect 16724 7936 16730 7948
rect 17129 7939 17187 7945
rect 17129 7936 17141 7939
rect 16724 7908 17141 7936
rect 16724 7896 16730 7908
rect 17129 7905 17141 7908
rect 17175 7905 17187 7939
rect 17129 7899 17187 7905
rect 17218 7896 17224 7948
rect 17276 7936 17282 7948
rect 17276 7908 17321 7936
rect 17276 7896 17282 7908
rect 2314 7868 2320 7880
rect 2275 7840 2320 7868
rect 2314 7828 2320 7840
rect 2372 7828 2378 7880
rect 5534 7868 5540 7880
rect 5495 7840 5540 7868
rect 5534 7828 5540 7840
rect 5592 7828 5598 7880
rect 5629 7871 5687 7877
rect 5629 7837 5641 7871
rect 5675 7837 5687 7871
rect 5629 7831 5687 7837
rect 5721 7871 5779 7877
rect 5721 7837 5733 7871
rect 5767 7837 5779 7871
rect 5721 7831 5779 7837
rect 5258 7760 5264 7812
rect 5316 7800 5322 7812
rect 5644 7800 5672 7831
rect 5316 7772 5672 7800
rect 5316 7760 5322 7772
rect 4062 7692 4068 7744
rect 4120 7732 4126 7744
rect 5736 7732 5764 7831
rect 5810 7828 5816 7880
rect 5868 7868 5874 7880
rect 7929 7871 7987 7877
rect 5868 7840 5913 7868
rect 5868 7828 5874 7840
rect 7929 7837 7941 7871
rect 7975 7868 7987 7871
rect 8202 7868 8208 7880
rect 7975 7840 8208 7868
rect 7975 7837 7987 7840
rect 7929 7831 7987 7837
rect 8202 7828 8208 7840
rect 8260 7828 8266 7880
rect 15010 7828 15016 7880
rect 15068 7868 15074 7880
rect 15289 7871 15347 7877
rect 15289 7868 15301 7871
rect 15068 7840 15301 7868
rect 15068 7828 15074 7840
rect 15289 7837 15301 7840
rect 15335 7837 15347 7871
rect 15289 7831 15347 7837
rect 10965 7803 11023 7809
rect 10965 7769 10977 7803
rect 11011 7800 11023 7803
rect 11330 7800 11336 7812
rect 11011 7772 11336 7800
rect 11011 7769 11023 7772
rect 10965 7763 11023 7769
rect 11330 7760 11336 7772
rect 11388 7760 11394 7812
rect 4120 7704 5764 7732
rect 4120 7692 4126 7704
rect 8662 7692 8668 7744
rect 8720 7732 8726 7744
rect 9306 7732 9312 7744
rect 8720 7704 9312 7732
rect 8720 7692 8726 7704
rect 9306 7692 9312 7704
rect 9364 7692 9370 7744
rect 184 7642 18860 7664
rect 184 7590 1556 7642
rect 1608 7590 1620 7642
rect 1672 7590 1684 7642
rect 1736 7590 1748 7642
rect 1800 7590 1812 7642
rect 1864 7590 4656 7642
rect 4708 7590 4720 7642
rect 4772 7590 4784 7642
rect 4836 7590 4848 7642
rect 4900 7590 4912 7642
rect 4964 7590 7756 7642
rect 7808 7590 7820 7642
rect 7872 7590 7884 7642
rect 7936 7590 7948 7642
rect 8000 7590 8012 7642
rect 8064 7590 10856 7642
rect 10908 7590 10920 7642
rect 10972 7590 10984 7642
rect 11036 7590 11048 7642
rect 11100 7590 11112 7642
rect 11164 7590 13956 7642
rect 14008 7590 14020 7642
rect 14072 7590 14084 7642
rect 14136 7590 14148 7642
rect 14200 7590 14212 7642
rect 14264 7590 17056 7642
rect 17108 7590 17120 7642
rect 17172 7590 17184 7642
rect 17236 7590 17248 7642
rect 17300 7590 17312 7642
rect 17364 7590 18860 7642
rect 184 7568 18860 7590
rect 3237 7531 3295 7537
rect 3237 7497 3249 7531
rect 3283 7528 3295 7531
rect 4338 7528 4344 7540
rect 3283 7500 4344 7528
rect 3283 7497 3295 7500
rect 3237 7491 3295 7497
rect 4338 7488 4344 7500
rect 4396 7488 4402 7540
rect 5626 7528 5632 7540
rect 5587 7500 5632 7528
rect 5626 7488 5632 7500
rect 5684 7488 5690 7540
rect 11330 7528 11336 7540
rect 11291 7500 11336 7528
rect 11330 7488 11336 7500
rect 11388 7488 11394 7540
rect 13722 7488 13728 7540
rect 13780 7528 13786 7540
rect 13780 7500 14228 7528
rect 13780 7488 13786 7500
rect 9030 7460 9036 7472
rect 8991 7432 9036 7460
rect 9030 7420 9036 7432
rect 9088 7420 9094 7472
rect 9585 7463 9643 7469
rect 9585 7460 9597 7463
rect 9232 7432 9597 7460
rect 2225 7395 2283 7401
rect 2225 7361 2237 7395
rect 2271 7392 2283 7395
rect 2406 7392 2412 7404
rect 2271 7364 2412 7392
rect 2271 7361 2283 7364
rect 2225 7355 2283 7361
rect 2406 7352 2412 7364
rect 2464 7352 2470 7404
rect 4062 7352 4068 7404
rect 4120 7392 4126 7404
rect 5077 7395 5135 7401
rect 5077 7392 5089 7395
rect 4120 7364 5089 7392
rect 4120 7352 4126 7364
rect 5077 7361 5089 7364
rect 5123 7361 5135 7395
rect 5077 7355 5135 7361
rect 5445 7395 5503 7401
rect 5445 7361 5457 7395
rect 5491 7392 5503 7395
rect 5810 7392 5816 7404
rect 5491 7364 5816 7392
rect 5491 7361 5503 7364
rect 5445 7355 5503 7361
rect 5810 7352 5816 7364
rect 5868 7352 5874 7404
rect 8662 7392 8668 7404
rect 6932 7364 8668 7392
rect 1949 7327 2007 7333
rect 1949 7293 1961 7327
rect 1995 7324 2007 7327
rect 2958 7324 2964 7336
rect 1995 7296 2964 7324
rect 1995 7293 2007 7296
rect 1949 7287 2007 7293
rect 2958 7284 2964 7296
rect 3016 7324 3022 7336
rect 3145 7327 3203 7333
rect 3145 7324 3157 7327
rect 3016 7296 3157 7324
rect 3016 7284 3022 7296
rect 3145 7293 3157 7296
rect 3191 7293 3203 7327
rect 3970 7324 3976 7336
rect 3931 7296 3976 7324
rect 3145 7287 3203 7293
rect 3970 7284 3976 7296
rect 4028 7284 4034 7336
rect 4157 7327 4215 7333
rect 4157 7293 4169 7327
rect 4203 7293 4215 7327
rect 4157 7287 4215 7293
rect 5537 7327 5595 7333
rect 5537 7293 5549 7327
rect 5583 7324 5595 7327
rect 5902 7324 5908 7336
rect 5583 7296 5908 7324
rect 5583 7293 5595 7296
rect 5537 7287 5595 7293
rect 2314 7216 2320 7268
rect 2372 7256 2378 7268
rect 4172 7256 4200 7287
rect 5902 7284 5908 7296
rect 5960 7324 5966 7336
rect 6822 7324 6828 7336
rect 5960 7296 6828 7324
rect 5960 7284 5966 7296
rect 6822 7284 6828 7296
rect 6880 7284 6886 7336
rect 6932 7333 6960 7364
rect 8662 7352 8668 7364
rect 8720 7352 8726 7404
rect 9232 7401 9260 7432
rect 9585 7429 9597 7432
rect 9631 7429 9643 7463
rect 13633 7463 13691 7469
rect 13633 7460 13645 7463
rect 9585 7423 9643 7429
rect 11992 7432 13645 7460
rect 8757 7395 8815 7401
rect 8757 7361 8769 7395
rect 8803 7392 8815 7395
rect 9217 7395 9275 7401
rect 8803 7364 8984 7392
rect 8803 7361 8815 7364
rect 8757 7355 8815 7361
rect 8956 7336 8984 7364
rect 9217 7361 9229 7395
rect 9263 7361 9275 7395
rect 9217 7355 9275 7361
rect 9306 7352 9312 7404
rect 9364 7392 9370 7404
rect 11149 7395 11207 7401
rect 9364 7364 9812 7392
rect 9364 7352 9370 7364
rect 6917 7327 6975 7333
rect 6917 7293 6929 7327
rect 6963 7293 6975 7327
rect 6917 7287 6975 7293
rect 7101 7327 7159 7333
rect 7101 7293 7113 7327
rect 7147 7324 7159 7327
rect 7282 7324 7288 7336
rect 7147 7296 7288 7324
rect 7147 7293 7159 7296
rect 7101 7287 7159 7293
rect 7282 7284 7288 7296
rect 7340 7284 7346 7336
rect 8110 7324 8116 7336
rect 7760 7296 8116 7324
rect 2372 7228 4200 7256
rect 4341 7259 4399 7265
rect 2372 7216 2378 7228
rect 4341 7225 4353 7259
rect 4387 7256 4399 7259
rect 4430 7256 4436 7268
rect 4387 7228 4436 7256
rect 4387 7225 4399 7228
rect 4341 7219 4399 7225
rect 4430 7216 4436 7228
rect 4488 7256 4494 7268
rect 5258 7256 5264 7268
rect 4488 7228 5264 7256
rect 4488 7216 4494 7228
rect 5258 7216 5264 7228
rect 5316 7216 5322 7268
rect 5353 7259 5411 7265
rect 5353 7225 5365 7259
rect 5399 7256 5411 7259
rect 5442 7256 5448 7268
rect 5399 7228 5448 7256
rect 5399 7225 5411 7228
rect 5353 7219 5411 7225
rect 5442 7216 5448 7228
rect 5500 7216 5506 7268
rect 6840 7256 6868 7284
rect 7760 7265 7788 7296
rect 8110 7284 8116 7296
rect 8168 7324 8174 7336
rect 8294 7324 8300 7336
rect 8168 7296 8300 7324
rect 8168 7284 8174 7296
rect 8294 7284 8300 7296
rect 8352 7284 8358 7336
rect 8849 7327 8907 7333
rect 8849 7293 8861 7327
rect 8895 7293 8907 7327
rect 8849 7287 8907 7293
rect 7745 7259 7803 7265
rect 7745 7256 7757 7259
rect 6840 7228 7757 7256
rect 7745 7225 7757 7228
rect 7791 7225 7803 7259
rect 8864 7256 8892 7287
rect 8938 7284 8944 7336
rect 8996 7284 9002 7336
rect 9784 7333 9812 7364
rect 11149 7361 11161 7395
rect 11195 7392 11207 7395
rect 11885 7395 11943 7401
rect 11885 7392 11897 7395
rect 11195 7364 11897 7392
rect 11195 7361 11207 7364
rect 11149 7355 11207 7361
rect 11885 7361 11897 7364
rect 11931 7361 11943 7395
rect 11885 7355 11943 7361
rect 9033 7327 9091 7333
rect 9033 7293 9045 7327
rect 9079 7293 9091 7327
rect 9585 7327 9643 7333
rect 9585 7324 9597 7327
rect 9033 7287 9091 7293
rect 9232 7296 9597 7324
rect 9048 7256 9076 7287
rect 9232 7268 9260 7296
rect 9585 7293 9597 7296
rect 9631 7293 9643 7327
rect 9585 7287 9643 7293
rect 9769 7327 9827 7333
rect 9769 7293 9781 7327
rect 9815 7293 9827 7327
rect 9769 7287 9827 7293
rect 11425 7327 11483 7333
rect 11425 7293 11437 7327
rect 11471 7324 11483 7327
rect 11992 7324 12020 7432
rect 13633 7429 13645 7432
rect 13679 7429 13691 7463
rect 13633 7423 13691 7429
rect 14093 7463 14151 7469
rect 14093 7429 14105 7463
rect 14139 7429 14151 7463
rect 14093 7423 14151 7429
rect 12894 7392 12900 7404
rect 12084 7364 12900 7392
rect 12084 7333 12112 7364
rect 12894 7352 12900 7364
rect 12952 7352 12958 7404
rect 11471 7296 12020 7324
rect 12069 7327 12127 7333
rect 11471 7293 11483 7296
rect 11425 7287 11483 7293
rect 12069 7293 12081 7327
rect 12115 7293 12127 7327
rect 12069 7287 12127 7293
rect 12158 7284 12164 7336
rect 12216 7324 12222 7336
rect 12289 7327 12347 7333
rect 12216 7296 12261 7324
rect 12216 7284 12222 7296
rect 12289 7293 12301 7327
rect 12335 7324 12347 7327
rect 12434 7324 12440 7336
rect 12335 7296 12440 7324
rect 12335 7293 12347 7296
rect 12289 7287 12347 7293
rect 12434 7284 12440 7296
rect 12492 7284 12498 7336
rect 13725 7327 13783 7333
rect 13725 7293 13737 7327
rect 13771 7324 13783 7327
rect 14108 7324 14136 7423
rect 14200 7392 14228 7500
rect 16666 7488 16672 7540
rect 16724 7528 16730 7540
rect 17773 7531 17831 7537
rect 17773 7528 17785 7531
rect 16724 7500 17785 7528
rect 16724 7488 16730 7500
rect 17773 7497 17785 7500
rect 17819 7497 17831 7531
rect 17773 7491 17831 7497
rect 14366 7392 14372 7404
rect 14200 7364 14372 7392
rect 14366 7352 14372 7364
rect 14424 7392 14430 7404
rect 14645 7395 14703 7401
rect 14645 7392 14657 7395
rect 14424 7364 14657 7392
rect 14424 7352 14430 7364
rect 14645 7361 14657 7364
rect 14691 7392 14703 7395
rect 15378 7392 15384 7404
rect 14691 7364 15384 7392
rect 14691 7361 14703 7364
rect 14645 7355 14703 7361
rect 15378 7352 15384 7364
rect 15436 7352 15442 7404
rect 16390 7392 16396 7404
rect 16351 7364 16396 7392
rect 16390 7352 16396 7364
rect 16448 7352 16454 7404
rect 13771 7296 14136 7324
rect 14553 7327 14611 7333
rect 13771 7293 13783 7296
rect 13725 7287 13783 7293
rect 14553 7293 14565 7327
rect 14599 7324 14611 7327
rect 15286 7324 15292 7336
rect 14599 7296 15292 7324
rect 14599 7293 14611 7296
rect 14553 7287 14611 7293
rect 15286 7284 15292 7296
rect 15344 7284 15350 7336
rect 7745 7219 7803 7225
rect 8312 7228 8892 7256
rect 8956 7228 9076 7256
rect 8312 7200 8340 7228
rect 8956 7200 8984 7228
rect 9214 7216 9220 7268
rect 9272 7216 9278 7268
rect 15194 7216 15200 7268
rect 15252 7256 15258 7268
rect 16298 7256 16304 7268
rect 15252 7228 16304 7256
rect 15252 7216 15258 7228
rect 16298 7216 16304 7228
rect 16356 7256 16362 7268
rect 16638 7259 16696 7265
rect 16638 7256 16650 7259
rect 16356 7228 16650 7256
rect 16356 7216 16362 7228
rect 16638 7225 16650 7228
rect 16684 7225 16696 7259
rect 16638 7219 16696 7225
rect 842 7148 848 7200
rect 900 7188 906 7200
rect 1581 7191 1639 7197
rect 1581 7188 1593 7191
rect 900 7160 1593 7188
rect 900 7148 906 7160
rect 1581 7157 1593 7160
rect 1627 7157 1639 7191
rect 1581 7151 1639 7157
rect 2041 7191 2099 7197
rect 2041 7157 2053 7191
rect 2087 7188 2099 7191
rect 2774 7188 2780 7200
rect 2087 7160 2780 7188
rect 2087 7157 2099 7160
rect 2041 7151 2099 7157
rect 2774 7148 2780 7160
rect 2832 7148 2838 7200
rect 7098 7188 7104 7200
rect 7059 7160 7104 7188
rect 7098 7148 7104 7160
rect 7156 7148 7162 7200
rect 7650 7188 7656 7200
rect 7611 7160 7656 7188
rect 7650 7148 7656 7160
rect 7708 7148 7714 7200
rect 8294 7188 8300 7200
rect 8255 7160 8300 7188
rect 8294 7148 8300 7160
rect 8352 7148 8358 7200
rect 8938 7148 8944 7200
rect 8996 7148 9002 7200
rect 9122 7188 9128 7200
rect 9083 7160 9128 7188
rect 9122 7148 9128 7160
rect 9180 7148 9186 7200
rect 11146 7188 11152 7200
rect 11107 7160 11152 7188
rect 11146 7148 11152 7160
rect 11204 7148 11210 7200
rect 14458 7188 14464 7200
rect 14419 7160 14464 7188
rect 14458 7148 14464 7160
rect 14516 7148 14522 7200
rect 184 7098 18920 7120
rect 184 7046 3106 7098
rect 3158 7046 3170 7098
rect 3222 7046 3234 7098
rect 3286 7046 3298 7098
rect 3350 7046 3362 7098
rect 3414 7046 6206 7098
rect 6258 7046 6270 7098
rect 6322 7046 6334 7098
rect 6386 7046 6398 7098
rect 6450 7046 6462 7098
rect 6514 7046 9306 7098
rect 9358 7046 9370 7098
rect 9422 7046 9434 7098
rect 9486 7046 9498 7098
rect 9550 7046 9562 7098
rect 9614 7046 12406 7098
rect 12458 7046 12470 7098
rect 12522 7046 12534 7098
rect 12586 7046 12598 7098
rect 12650 7046 12662 7098
rect 12714 7046 15506 7098
rect 15558 7046 15570 7098
rect 15622 7046 15634 7098
rect 15686 7046 15698 7098
rect 15750 7046 15762 7098
rect 15814 7046 18606 7098
rect 18658 7046 18670 7098
rect 18722 7046 18734 7098
rect 18786 7046 18798 7098
rect 18850 7046 18862 7098
rect 18914 7046 18920 7098
rect 184 7024 18920 7046
rect 2317 6987 2375 6993
rect 2317 6953 2329 6987
rect 2363 6953 2375 6987
rect 2317 6947 2375 6953
rect 2130 6916 2136 6928
rect 2070 6888 2136 6916
rect 2130 6876 2136 6888
rect 2188 6876 2194 6928
rect 2332 6916 2360 6947
rect 2774 6944 2780 6996
rect 2832 6984 2838 6996
rect 3145 6987 3203 6993
rect 2832 6956 2877 6984
rect 2832 6944 2838 6956
rect 3145 6953 3157 6987
rect 3191 6984 3203 6987
rect 4338 6984 4344 6996
rect 3191 6956 4344 6984
rect 3191 6953 3203 6956
rect 3145 6947 3203 6953
rect 4338 6944 4344 6956
rect 4396 6944 4402 6996
rect 8202 6984 8208 6996
rect 8163 6956 8208 6984
rect 8202 6944 8208 6956
rect 8260 6944 8266 6996
rect 10778 6944 10784 6996
rect 10836 6984 10842 6996
rect 11698 6984 11704 6996
rect 10836 6956 11704 6984
rect 10836 6944 10842 6956
rect 11698 6944 11704 6956
rect 11756 6984 11762 6996
rect 11756 6956 12434 6984
rect 11756 6944 11762 6956
rect 2958 6916 2964 6928
rect 2332 6888 2964 6916
rect 2958 6876 2964 6888
rect 3016 6876 3022 6928
rect 4157 6919 4215 6925
rect 4157 6885 4169 6919
rect 4203 6916 4215 6919
rect 6638 6916 6644 6928
rect 4203 6888 6644 6916
rect 4203 6885 4215 6888
rect 4157 6879 4215 6885
rect 566 6848 572 6860
rect 527 6820 572 6848
rect 566 6808 572 6820
rect 624 6808 630 6860
rect 6472 6857 6500 6888
rect 6638 6876 6644 6888
rect 6696 6916 6702 6928
rect 6696 6888 7052 6916
rect 6696 6876 6702 6888
rect 6457 6851 6515 6857
rect 6457 6817 6469 6851
rect 6503 6817 6515 6851
rect 6457 6811 6515 6817
rect 6732 6851 6790 6857
rect 6732 6817 6744 6851
rect 6778 6817 6790 6851
rect 6732 6811 6790 6817
rect 842 6780 848 6792
rect 803 6752 848 6780
rect 842 6740 848 6752
rect 900 6740 906 6792
rect 2222 6740 2228 6792
rect 2280 6780 2286 6792
rect 3237 6783 3295 6789
rect 3237 6780 3249 6783
rect 2280 6752 3249 6780
rect 2280 6740 2286 6752
rect 3237 6749 3249 6752
rect 3283 6749 3295 6783
rect 3237 6743 3295 6749
rect 3421 6783 3479 6789
rect 3421 6749 3433 6783
rect 3467 6780 3479 6783
rect 3510 6780 3516 6792
rect 3467 6752 3516 6780
rect 3467 6749 3479 6752
rect 3421 6743 3479 6749
rect 3510 6740 3516 6752
rect 3568 6780 3574 6792
rect 4249 6783 4307 6789
rect 4249 6780 4261 6783
rect 3568 6752 4261 6780
rect 3568 6740 3574 6752
rect 4249 6749 4261 6752
rect 4295 6749 4307 6783
rect 4249 6743 4307 6749
rect 4338 6740 4344 6792
rect 4396 6780 4402 6792
rect 6748 6780 6776 6811
rect 6822 6808 6828 6860
rect 6880 6848 6886 6860
rect 7024 6848 7052 6888
rect 7098 6876 7104 6928
rect 7156 6916 7162 6928
rect 11790 6916 11796 6928
rect 7156 6888 7972 6916
rect 11638 6888 11796 6916
rect 7156 6876 7162 6888
rect 6880 6820 6925 6848
rect 7024 6820 7420 6848
rect 6880 6808 6886 6820
rect 7282 6780 7288 6792
rect 4396 6752 4441 6780
rect 6748 6752 7288 6780
rect 4396 6740 4402 6752
rect 7282 6740 7288 6752
rect 7340 6740 7346 6792
rect 7392 6780 7420 6820
rect 7466 6808 7472 6860
rect 7524 6848 7530 6860
rect 7944 6857 7972 6888
rect 11790 6876 11796 6888
rect 11848 6916 11854 6928
rect 12066 6916 12072 6928
rect 11848 6888 12072 6916
rect 11848 6876 11854 6888
rect 12066 6876 12072 6888
rect 12124 6876 12130 6928
rect 7653 6851 7711 6857
rect 7653 6848 7665 6851
rect 7524 6820 7665 6848
rect 7524 6808 7530 6820
rect 7653 6817 7665 6820
rect 7699 6817 7711 6851
rect 7653 6811 7711 6817
rect 7929 6851 7987 6857
rect 7929 6817 7941 6851
rect 7975 6817 7987 6851
rect 8481 6851 8539 6857
rect 8481 6848 8493 6851
rect 7929 6811 7987 6817
rect 8128 6820 8493 6848
rect 7561 6783 7619 6789
rect 7561 6780 7573 6783
rect 7392 6752 7573 6780
rect 7561 6749 7573 6752
rect 7607 6749 7619 6783
rect 7561 6743 7619 6749
rect 7742 6740 7748 6792
rect 7800 6780 7806 6792
rect 8021 6783 8079 6789
rect 8021 6780 8033 6783
rect 7800 6752 8033 6780
rect 7800 6740 7806 6752
rect 8021 6749 8033 6752
rect 8067 6749 8079 6783
rect 8021 6743 8079 6749
rect 2406 6672 2412 6724
rect 2464 6712 2470 6724
rect 3789 6715 3847 6721
rect 3789 6712 3801 6715
rect 2464 6684 3801 6712
rect 2464 6672 2470 6684
rect 3789 6681 3801 6684
rect 3835 6681 3847 6715
rect 7300 6712 7328 6740
rect 8128 6712 8156 6820
rect 8481 6817 8493 6820
rect 8527 6817 8539 6851
rect 8481 6811 8539 6817
rect 8665 6851 8723 6857
rect 8665 6817 8677 6851
rect 8711 6848 8723 6851
rect 9214 6848 9220 6860
rect 8711 6820 9220 6848
rect 8711 6817 8723 6820
rect 8665 6811 8723 6817
rect 9214 6808 9220 6820
rect 9272 6808 9278 6860
rect 12406 6848 12434 6956
rect 14458 6944 14464 6996
rect 14516 6984 14522 6996
rect 14737 6987 14795 6993
rect 14737 6984 14749 6987
rect 14516 6956 14749 6984
rect 14516 6944 14522 6956
rect 14737 6953 14749 6956
rect 14783 6953 14795 6987
rect 15194 6984 15200 6996
rect 14737 6947 14795 6953
rect 14936 6956 15200 6984
rect 12897 6851 12955 6857
rect 12897 6848 12909 6851
rect 12406 6820 12909 6848
rect 12897 6817 12909 6820
rect 12943 6817 12955 6851
rect 12897 6811 12955 6817
rect 13357 6851 13415 6857
rect 13357 6817 13369 6851
rect 13403 6848 13415 6851
rect 13725 6851 13783 6857
rect 13403 6820 13676 6848
rect 13403 6817 13415 6820
rect 13357 6811 13415 6817
rect 10042 6740 10048 6792
rect 10100 6780 10106 6792
rect 10137 6783 10195 6789
rect 10137 6780 10149 6783
rect 10100 6752 10149 6780
rect 10100 6740 10106 6752
rect 10137 6749 10149 6752
rect 10183 6749 10195 6783
rect 10137 6743 10195 6749
rect 10413 6783 10471 6789
rect 10413 6749 10425 6783
rect 10459 6780 10471 6783
rect 11146 6780 11152 6792
rect 10459 6752 11152 6780
rect 10459 6749 10471 6752
rect 10413 6743 10471 6749
rect 11146 6740 11152 6752
rect 11204 6740 11210 6792
rect 11885 6783 11943 6789
rect 11885 6749 11897 6783
rect 11931 6780 11943 6783
rect 12158 6780 12164 6792
rect 11931 6752 12164 6780
rect 11931 6749 11943 6752
rect 11885 6743 11943 6749
rect 12158 6740 12164 6752
rect 12216 6740 12222 6792
rect 13446 6780 13452 6792
rect 12406 6752 13124 6780
rect 13407 6752 13452 6780
rect 7300 6684 8156 6712
rect 3789 6675 3847 6681
rect 8846 6672 8852 6724
rect 8904 6712 8910 6724
rect 12406 6712 12434 6752
rect 8904 6684 9076 6712
rect 8904 6672 8910 6684
rect 8570 6644 8576 6656
rect 8531 6616 8576 6644
rect 8570 6604 8576 6616
rect 8628 6604 8634 6656
rect 8938 6644 8944 6656
rect 8899 6616 8944 6644
rect 8938 6604 8944 6616
rect 8996 6604 9002 6656
rect 9048 6644 9076 6684
rect 11440 6684 12434 6712
rect 12621 6715 12679 6721
rect 11440 6644 11468 6684
rect 12621 6681 12633 6715
rect 12667 6712 12679 6715
rect 12894 6712 12900 6724
rect 12667 6684 12900 6712
rect 12667 6681 12679 6684
rect 12621 6675 12679 6681
rect 12894 6672 12900 6684
rect 12952 6672 12958 6724
rect 13096 6712 13124 6752
rect 13446 6740 13452 6752
rect 13504 6740 13510 6792
rect 13648 6780 13676 6820
rect 13725 6817 13737 6851
rect 13771 6848 13783 6851
rect 14936 6848 14964 6956
rect 15194 6944 15200 6956
rect 15252 6944 15258 6996
rect 15010 6876 15016 6928
rect 15068 6916 15074 6928
rect 15068 6888 15332 6916
rect 15068 6876 15074 6888
rect 15102 6848 15108 6860
rect 13771 6820 14964 6848
rect 15063 6820 15108 6848
rect 13771 6817 13783 6820
rect 13725 6811 13783 6817
rect 15102 6808 15108 6820
rect 15160 6808 15166 6860
rect 15194 6780 15200 6792
rect 13648 6752 15200 6780
rect 15194 6740 15200 6752
rect 15252 6740 15258 6792
rect 15304 6789 15332 6888
rect 15378 6808 15384 6860
rect 15436 6848 15442 6860
rect 17221 6851 17279 6857
rect 17221 6848 17233 6851
rect 15436 6820 17233 6848
rect 15436 6808 15442 6820
rect 17221 6817 17233 6820
rect 17267 6817 17279 6851
rect 17221 6811 17279 6817
rect 17957 6851 18015 6857
rect 17957 6817 17969 6851
rect 18003 6848 18015 6851
rect 18414 6848 18420 6860
rect 18003 6820 18420 6848
rect 18003 6817 18015 6820
rect 17957 6811 18015 6817
rect 18414 6808 18420 6820
rect 18472 6808 18478 6860
rect 15289 6783 15347 6789
rect 15289 6749 15301 6783
rect 15335 6749 15347 6783
rect 15289 6743 15347 6749
rect 18233 6715 18291 6721
rect 18233 6712 18245 6715
rect 13096 6684 18245 6712
rect 18233 6681 18245 6684
rect 18279 6681 18291 6715
rect 18233 6675 18291 6681
rect 9048 6616 11468 6644
rect 16758 6604 16764 6656
rect 16816 6644 16822 6656
rect 17313 6647 17371 6653
rect 17313 6644 17325 6647
rect 16816 6616 17325 6644
rect 16816 6604 16822 6616
rect 17313 6613 17325 6616
rect 17359 6613 17371 6647
rect 17313 6607 17371 6613
rect 184 6554 18860 6576
rect 184 6502 1556 6554
rect 1608 6502 1620 6554
rect 1672 6502 1684 6554
rect 1736 6502 1748 6554
rect 1800 6502 1812 6554
rect 1864 6502 4656 6554
rect 4708 6502 4720 6554
rect 4772 6502 4784 6554
rect 4836 6502 4848 6554
rect 4900 6502 4912 6554
rect 4964 6502 7756 6554
rect 7808 6502 7820 6554
rect 7872 6502 7884 6554
rect 7936 6502 7948 6554
rect 8000 6502 8012 6554
rect 8064 6502 10856 6554
rect 10908 6502 10920 6554
rect 10972 6502 10984 6554
rect 11036 6502 11048 6554
rect 11100 6502 11112 6554
rect 11164 6502 13956 6554
rect 14008 6502 14020 6554
rect 14072 6502 14084 6554
rect 14136 6502 14148 6554
rect 14200 6502 14212 6554
rect 14264 6502 17056 6554
rect 17108 6502 17120 6554
rect 17172 6502 17184 6554
rect 17236 6502 17248 6554
rect 17300 6502 17312 6554
rect 17364 6502 18860 6554
rect 184 6480 18860 6502
rect 2222 6440 2228 6452
rect 2183 6412 2228 6440
rect 2222 6400 2228 6412
rect 2280 6400 2286 6452
rect 2685 6443 2743 6449
rect 2685 6409 2697 6443
rect 2731 6440 2743 6443
rect 2731 6412 4752 6440
rect 2731 6409 2743 6412
rect 2685 6403 2743 6409
rect 2041 6307 2099 6313
rect 2041 6273 2053 6307
rect 2087 6304 2099 6307
rect 2700 6304 2728 6403
rect 2087 6276 2728 6304
rect 4065 6307 4123 6313
rect 2087 6273 2099 6276
rect 2041 6267 2099 6273
rect 4065 6273 4077 6307
rect 4111 6304 4123 6307
rect 4246 6304 4252 6316
rect 4111 6276 4252 6304
rect 4111 6273 4123 6276
rect 4065 6267 4123 6273
rect 4246 6264 4252 6276
rect 4304 6264 4310 6316
rect 4724 6313 4752 6412
rect 5166 6400 5172 6452
rect 5224 6440 5230 6452
rect 5813 6443 5871 6449
rect 5813 6440 5825 6443
rect 5224 6412 5825 6440
rect 5224 6400 5230 6412
rect 5813 6409 5825 6412
rect 5859 6440 5871 6443
rect 6086 6440 6092 6452
rect 5859 6412 6092 6440
rect 5859 6409 5871 6412
rect 5813 6403 5871 6409
rect 6086 6400 6092 6412
rect 6144 6440 6150 6452
rect 8938 6440 8944 6452
rect 6144 6412 8944 6440
rect 6144 6400 6150 6412
rect 8938 6400 8944 6412
rect 8996 6400 9002 6452
rect 13446 6400 13452 6452
rect 13504 6440 13510 6452
rect 14277 6443 14335 6449
rect 14277 6440 14289 6443
rect 13504 6412 14289 6440
rect 13504 6400 13510 6412
rect 14277 6409 14289 6412
rect 14323 6440 14335 6443
rect 14550 6440 14556 6452
rect 14323 6412 14556 6440
rect 14323 6409 14335 6412
rect 14277 6403 14335 6409
rect 14550 6400 14556 6412
rect 14608 6400 14614 6452
rect 14921 6443 14979 6449
rect 14921 6409 14933 6443
rect 14967 6440 14979 6443
rect 15102 6440 15108 6452
rect 14967 6412 15108 6440
rect 14967 6409 14979 6412
rect 14921 6403 14979 6409
rect 15102 6400 15108 6412
rect 15160 6400 15166 6452
rect 4709 6307 4767 6313
rect 4709 6273 4721 6307
rect 4755 6304 4767 6307
rect 5184 6304 5212 6400
rect 8294 6372 8300 6384
rect 4755 6276 5212 6304
rect 6380 6344 8300 6372
rect 4755 6273 4767 6276
rect 4709 6267 4767 6273
rect 1949 6239 2007 6245
rect 1949 6205 1961 6239
rect 1995 6236 2007 6239
rect 2222 6236 2228 6248
rect 1995 6208 2228 6236
rect 1995 6205 2007 6208
rect 1949 6199 2007 6205
rect 2222 6196 2228 6208
rect 2280 6236 2286 6248
rect 2961 6239 3019 6245
rect 2961 6236 2973 6239
rect 2280 6208 2973 6236
rect 2280 6196 2286 6208
rect 2961 6205 2973 6208
rect 3007 6205 3019 6239
rect 4430 6236 4436 6248
rect 4391 6208 4436 6236
rect 2961 6199 3019 6205
rect 2976 6168 3004 6199
rect 4430 6196 4436 6208
rect 4488 6196 4494 6248
rect 4982 6236 4988 6248
rect 4895 6208 4988 6236
rect 4982 6196 4988 6208
rect 5040 6196 5046 6248
rect 5074 6196 5080 6248
rect 5132 6236 5138 6248
rect 5442 6236 5448 6248
rect 5132 6208 5448 6236
rect 5132 6196 5138 6208
rect 5442 6196 5448 6208
rect 5500 6196 5506 6248
rect 5000 6168 5028 6196
rect 6380 6177 6408 6344
rect 8294 6332 8300 6344
rect 8352 6332 8358 6384
rect 8113 6307 8171 6313
rect 8113 6273 8125 6307
rect 8159 6304 8171 6307
rect 8754 6304 8760 6316
rect 8159 6276 8760 6304
rect 8159 6273 8171 6276
rect 8113 6267 8171 6273
rect 8754 6264 8760 6276
rect 8812 6264 8818 6316
rect 12158 6264 12164 6316
rect 12216 6304 12222 6316
rect 14274 6304 14280 6316
rect 12216 6276 14280 6304
rect 12216 6264 12222 6276
rect 14274 6264 14280 6276
rect 14332 6304 14338 6316
rect 16117 6307 16175 6313
rect 14332 6276 14780 6304
rect 14332 6264 14338 6276
rect 7650 6196 7656 6248
rect 7708 6236 7714 6248
rect 7745 6239 7803 6245
rect 7745 6236 7757 6239
rect 7708 6208 7757 6236
rect 7708 6196 7714 6208
rect 7745 6205 7757 6208
rect 7791 6205 7803 6239
rect 7745 6199 7803 6205
rect 7837 6239 7895 6245
rect 7837 6205 7849 6239
rect 7883 6236 7895 6239
rect 8570 6236 8576 6248
rect 7883 6208 8576 6236
rect 7883 6205 7895 6208
rect 7837 6199 7895 6205
rect 8570 6196 8576 6208
rect 8628 6196 8634 6248
rect 12805 6239 12863 6245
rect 12805 6205 12817 6239
rect 12851 6236 12863 6239
rect 12894 6236 12900 6248
rect 12851 6208 12900 6236
rect 12851 6205 12863 6208
rect 12805 6199 12863 6205
rect 12894 6196 12900 6208
rect 12952 6196 12958 6248
rect 14752 6245 14780 6276
rect 16117 6273 16129 6307
rect 16163 6304 16175 6307
rect 16390 6304 16396 6316
rect 16163 6276 16396 6304
rect 16163 6273 16175 6276
rect 16117 6267 16175 6273
rect 16390 6264 16396 6276
rect 16448 6264 16454 6316
rect 14737 6239 14795 6245
rect 14737 6205 14749 6239
rect 14783 6205 14795 6239
rect 16482 6236 16488 6248
rect 16443 6208 16488 6236
rect 14737 6199 14795 6205
rect 16482 6196 16488 6208
rect 16540 6196 16546 6248
rect 17500 6180 17552 6186
rect 6365 6171 6423 6177
rect 6365 6168 6377 6171
rect 2976 6140 6377 6168
rect 6365 6137 6377 6140
rect 6411 6137 6423 6171
rect 6365 6131 6423 6137
rect 6638 6128 6644 6180
rect 6696 6168 6702 6180
rect 6822 6168 6828 6180
rect 6696 6140 6828 6168
rect 6696 6128 6702 6140
rect 6822 6128 6828 6140
rect 6880 6168 6886 6180
rect 8205 6171 8263 6177
rect 8205 6168 8217 6171
rect 6880 6140 8217 6168
rect 6880 6128 6886 6140
rect 8205 6137 8217 6140
rect 8251 6137 8263 6171
rect 8205 6131 8263 6137
rect 15565 6171 15623 6177
rect 15565 6137 15577 6171
rect 15611 6168 15623 6171
rect 16022 6168 16028 6180
rect 15611 6140 16028 6168
rect 15611 6137 15623 6140
rect 15565 6131 15623 6137
rect 16022 6128 16028 6140
rect 16080 6128 16086 6180
rect 17954 6168 17960 6180
rect 17915 6140 17960 6168
rect 17954 6128 17960 6140
rect 18012 6128 18018 6180
rect 17500 6122 17552 6128
rect 7561 6103 7619 6109
rect 7561 6069 7573 6103
rect 7607 6100 7619 6103
rect 8018 6100 8024 6112
rect 7607 6072 8024 6100
rect 7607 6069 7619 6072
rect 7561 6063 7619 6069
rect 8018 6060 8024 6072
rect 8076 6060 8082 6112
rect 12066 6100 12072 6112
rect 12027 6072 12072 6100
rect 12066 6060 12072 6072
rect 12124 6060 12130 6112
rect 12897 6103 12955 6109
rect 12897 6069 12909 6103
rect 12943 6100 12955 6103
rect 13262 6100 13268 6112
rect 12943 6072 13268 6100
rect 12943 6069 12955 6072
rect 12897 6063 12955 6069
rect 13262 6060 13268 6072
rect 13320 6060 13326 6112
rect 14550 6060 14556 6112
rect 14608 6100 14614 6112
rect 16942 6100 16948 6112
rect 14608 6072 16948 6100
rect 14608 6060 14614 6072
rect 16942 6060 16948 6072
rect 17000 6060 17006 6112
rect 184 6010 18920 6032
rect 184 5958 3106 6010
rect 3158 5958 3170 6010
rect 3222 5958 3234 6010
rect 3286 5958 3298 6010
rect 3350 5958 3362 6010
rect 3414 5958 6206 6010
rect 6258 5958 6270 6010
rect 6322 5958 6334 6010
rect 6386 5958 6398 6010
rect 6450 5958 6462 6010
rect 6514 5958 9306 6010
rect 9358 5958 9370 6010
rect 9422 5958 9434 6010
rect 9486 5958 9498 6010
rect 9550 5958 9562 6010
rect 9614 5958 12406 6010
rect 12458 5958 12470 6010
rect 12522 5958 12534 6010
rect 12586 5958 12598 6010
rect 12650 5958 12662 6010
rect 12714 5958 15506 6010
rect 15558 5958 15570 6010
rect 15622 5958 15634 6010
rect 15686 5958 15698 6010
rect 15750 5958 15762 6010
rect 15814 5958 18606 6010
rect 18658 5958 18670 6010
rect 18722 5958 18734 6010
rect 18786 5958 18798 6010
rect 18850 5958 18862 6010
rect 18914 5958 18920 6010
rect 184 5936 18920 5958
rect 4157 5899 4215 5905
rect 4157 5865 4169 5899
rect 4203 5896 4215 5899
rect 4338 5896 4344 5908
rect 4203 5868 4344 5896
rect 4203 5865 4215 5868
rect 4157 5859 4215 5865
rect 4338 5856 4344 5868
rect 4396 5856 4402 5908
rect 4430 5856 4436 5908
rect 4488 5896 4494 5908
rect 5258 5896 5264 5908
rect 4488 5868 5264 5896
rect 4488 5856 4494 5868
rect 5258 5856 5264 5868
rect 5316 5896 5322 5908
rect 5353 5899 5411 5905
rect 5353 5896 5365 5899
rect 5316 5868 5365 5896
rect 5316 5856 5322 5868
rect 5353 5865 5365 5868
rect 5399 5865 5411 5899
rect 5353 5859 5411 5865
rect 16482 5856 16488 5908
rect 16540 5896 16546 5908
rect 17129 5899 17187 5905
rect 17129 5896 17141 5899
rect 16540 5868 17141 5896
rect 16540 5856 16546 5868
rect 17129 5865 17141 5868
rect 17175 5865 17187 5899
rect 17129 5859 17187 5865
rect 3510 5788 3516 5840
rect 3568 5828 3574 5840
rect 5169 5831 5227 5837
rect 5169 5828 5181 5831
rect 3568 5800 5181 5828
rect 3568 5788 3574 5800
rect 5169 5797 5181 5800
rect 5215 5828 5227 5831
rect 7650 5828 7656 5840
rect 5215 5800 7656 5828
rect 5215 5797 5227 5800
rect 5169 5791 5227 5797
rect 7650 5788 7656 5800
rect 7708 5788 7714 5840
rect 8018 5828 8024 5840
rect 7979 5800 8024 5828
rect 8018 5788 8024 5800
rect 8076 5788 8082 5840
rect 8478 5788 8484 5840
rect 8536 5788 8542 5840
rect 12066 5828 12072 5840
rect 11546 5800 12072 5828
rect 12066 5788 12072 5800
rect 12124 5788 12130 5840
rect 15194 5788 15200 5840
rect 15252 5828 15258 5840
rect 16942 5828 16948 5840
rect 15252 5800 16252 5828
rect 15252 5788 15258 5800
rect 566 5720 572 5772
rect 624 5760 630 5772
rect 1857 5763 1915 5769
rect 1857 5760 1869 5763
rect 624 5732 1869 5760
rect 624 5720 630 5732
rect 1857 5729 1869 5732
rect 1903 5729 1915 5763
rect 4246 5760 4252 5772
rect 4207 5732 4252 5760
rect 1857 5723 1915 5729
rect 4246 5720 4252 5732
rect 4304 5720 4310 5772
rect 5445 5763 5503 5769
rect 5445 5729 5457 5763
rect 5491 5760 5503 5763
rect 5534 5760 5540 5772
rect 5491 5732 5540 5760
rect 5491 5729 5503 5732
rect 5445 5723 5503 5729
rect 5534 5720 5540 5732
rect 5592 5720 5598 5772
rect 5902 5720 5908 5772
rect 5960 5760 5966 5772
rect 6181 5763 6239 5769
rect 6181 5760 6193 5763
rect 5960 5732 6193 5760
rect 5960 5720 5966 5732
rect 6181 5729 6193 5732
rect 6227 5729 6239 5763
rect 6181 5723 6239 5729
rect 7558 5720 7564 5772
rect 7616 5760 7622 5772
rect 7745 5763 7803 5769
rect 7745 5760 7757 5763
rect 7616 5732 7757 5760
rect 7616 5720 7622 5732
rect 7745 5729 7757 5732
rect 7791 5729 7803 5763
rect 13081 5763 13139 5769
rect 13081 5760 13093 5763
rect 7745 5723 7803 5729
rect 13004 5732 13093 5760
rect 5552 5692 5580 5720
rect 6273 5695 6331 5701
rect 6273 5692 6285 5695
rect 5552 5664 6285 5692
rect 6273 5661 6285 5664
rect 6319 5661 6331 5695
rect 6273 5655 6331 5661
rect 6457 5695 6515 5701
rect 6457 5661 6469 5695
rect 6503 5692 6515 5695
rect 6546 5692 6552 5704
rect 6503 5664 6552 5692
rect 6503 5661 6515 5664
rect 6457 5655 6515 5661
rect 6546 5652 6552 5664
rect 6604 5652 6610 5704
rect 10042 5692 10048 5704
rect 10003 5664 10048 5692
rect 10042 5652 10048 5664
rect 10100 5652 10106 5704
rect 10321 5695 10379 5701
rect 10321 5661 10333 5695
rect 10367 5692 10379 5695
rect 11330 5692 11336 5704
rect 10367 5664 11336 5692
rect 10367 5661 10379 5664
rect 10321 5655 10379 5661
rect 11330 5652 11336 5664
rect 11388 5652 11394 5704
rect 13004 5624 13032 5732
rect 13081 5729 13093 5732
rect 13127 5729 13139 5763
rect 13725 5763 13783 5769
rect 13725 5760 13737 5763
rect 13081 5723 13139 5729
rect 13188 5732 13737 5760
rect 13188 5704 13216 5732
rect 13725 5729 13737 5732
rect 13771 5729 13783 5763
rect 13725 5723 13783 5729
rect 13814 5720 13820 5772
rect 13872 5760 13878 5772
rect 15289 5763 15347 5769
rect 13872 5732 13917 5760
rect 13872 5720 13878 5732
rect 15289 5729 15301 5763
rect 15335 5729 15347 5763
rect 15289 5723 15347 5729
rect 15473 5763 15531 5769
rect 15473 5729 15485 5763
rect 15519 5760 15531 5763
rect 15654 5760 15660 5772
rect 15519 5732 15660 5760
rect 15519 5729 15531 5732
rect 15473 5723 15531 5729
rect 13170 5692 13176 5704
rect 13131 5664 13176 5692
rect 13170 5652 13176 5664
rect 13228 5652 13234 5704
rect 13262 5652 13268 5704
rect 13320 5692 13326 5704
rect 13320 5664 13365 5692
rect 13320 5652 13326 5664
rect 14093 5627 14151 5633
rect 14093 5624 14105 5627
rect 13004 5596 14105 5624
rect 14093 5593 14105 5596
rect 14139 5624 14151 5627
rect 14918 5624 14924 5636
rect 14139 5596 14924 5624
rect 14139 5593 14151 5596
rect 14093 5587 14151 5593
rect 14918 5584 14924 5596
rect 14976 5584 14982 5636
rect 1946 5516 1952 5568
rect 2004 5556 2010 5568
rect 2041 5559 2099 5565
rect 2041 5556 2053 5559
rect 2004 5528 2053 5556
rect 2004 5516 2010 5528
rect 2041 5525 2053 5528
rect 2087 5525 2099 5559
rect 2041 5519 2099 5525
rect 5074 5516 5080 5568
rect 5132 5556 5138 5568
rect 5169 5559 5227 5565
rect 5169 5556 5181 5559
rect 5132 5528 5181 5556
rect 5132 5516 5138 5528
rect 5169 5525 5181 5528
rect 5215 5525 5227 5559
rect 5169 5519 5227 5525
rect 6365 5559 6423 5565
rect 6365 5525 6377 5559
rect 6411 5556 6423 5559
rect 6730 5556 6736 5568
rect 6411 5528 6736 5556
rect 6411 5525 6423 5528
rect 6365 5519 6423 5525
rect 6730 5516 6736 5528
rect 6788 5516 6794 5568
rect 9214 5516 9220 5568
rect 9272 5556 9278 5568
rect 9493 5559 9551 5565
rect 9493 5556 9505 5559
rect 9272 5528 9505 5556
rect 9272 5516 9278 5528
rect 9493 5525 9505 5528
rect 9539 5525 9551 5559
rect 9493 5519 9551 5525
rect 11514 5516 11520 5568
rect 11572 5556 11578 5568
rect 11793 5559 11851 5565
rect 11793 5556 11805 5559
rect 11572 5528 11805 5556
rect 11572 5516 11578 5528
rect 11793 5525 11805 5528
rect 11839 5525 11851 5559
rect 11793 5519 11851 5525
rect 12066 5516 12072 5568
rect 12124 5556 12130 5568
rect 12434 5556 12440 5568
rect 12124 5528 12440 5556
rect 12124 5516 12130 5528
rect 12434 5516 12440 5528
rect 12492 5516 12498 5568
rect 12710 5556 12716 5568
rect 12671 5528 12716 5556
rect 12710 5516 12716 5528
rect 12768 5516 12774 5568
rect 15304 5556 15332 5723
rect 15654 5720 15660 5732
rect 15712 5720 15718 5772
rect 15749 5763 15807 5769
rect 15749 5729 15761 5763
rect 15795 5729 15807 5763
rect 15749 5723 15807 5729
rect 15381 5695 15439 5701
rect 15381 5661 15393 5695
rect 15427 5692 15439 5695
rect 15764 5692 15792 5723
rect 15838 5720 15844 5772
rect 15896 5760 15902 5772
rect 16224 5769 16252 5800
rect 16684 5800 16948 5828
rect 15933 5763 15991 5769
rect 15933 5760 15945 5763
rect 15896 5732 15945 5760
rect 15896 5720 15902 5732
rect 15933 5729 15945 5732
rect 15979 5729 15991 5763
rect 15933 5723 15991 5729
rect 16209 5763 16267 5769
rect 16209 5729 16221 5763
rect 16255 5729 16267 5763
rect 16209 5723 16267 5729
rect 16298 5720 16304 5772
rect 16356 5760 16362 5772
rect 16684 5769 16712 5800
rect 16942 5788 16948 5800
rect 17000 5828 17006 5840
rect 18049 5831 18107 5837
rect 18049 5828 18061 5831
rect 17000 5800 18061 5828
rect 17000 5788 17006 5800
rect 18049 5797 18061 5800
rect 18095 5797 18107 5831
rect 18049 5791 18107 5797
rect 16393 5763 16451 5769
rect 16393 5760 16405 5763
rect 16356 5732 16405 5760
rect 16356 5720 16362 5732
rect 16393 5729 16405 5732
rect 16439 5729 16451 5763
rect 16393 5723 16451 5729
rect 16669 5763 16727 5769
rect 16669 5729 16681 5763
rect 16715 5729 16727 5763
rect 16669 5723 16727 5729
rect 16758 5720 16764 5772
rect 16816 5760 16822 5772
rect 17313 5763 17371 5769
rect 17313 5760 17325 5763
rect 16816 5732 17325 5760
rect 16816 5720 16822 5732
rect 17313 5729 17325 5732
rect 17359 5729 17371 5763
rect 17313 5723 17371 5729
rect 17402 5720 17408 5772
rect 17460 5760 17466 5772
rect 17497 5763 17555 5769
rect 17497 5760 17509 5763
rect 17460 5732 17509 5760
rect 17460 5720 17466 5732
rect 17497 5729 17509 5732
rect 17543 5729 17555 5763
rect 17497 5723 17555 5729
rect 17589 5763 17647 5769
rect 17589 5729 17601 5763
rect 17635 5729 17647 5763
rect 17589 5723 17647 5729
rect 17604 5692 17632 5723
rect 15427 5664 15792 5692
rect 16776 5664 17632 5692
rect 15427 5661 15439 5664
rect 15381 5655 15439 5661
rect 15841 5627 15899 5633
rect 15841 5593 15853 5627
rect 15887 5624 15899 5627
rect 15930 5624 15936 5636
rect 15887 5596 15936 5624
rect 15887 5593 15899 5596
rect 15841 5587 15899 5593
rect 15930 5584 15936 5596
rect 15988 5584 15994 5636
rect 16298 5584 16304 5636
rect 16356 5624 16362 5636
rect 16776 5624 16804 5664
rect 17954 5652 17960 5704
rect 18012 5652 18018 5704
rect 16356 5596 16804 5624
rect 17405 5627 17463 5633
rect 16356 5584 16362 5596
rect 17405 5593 17417 5627
rect 17451 5593 17463 5627
rect 17972 5624 18000 5652
rect 17405 5587 17463 5593
rect 17604 5596 18000 5624
rect 17420 5556 17448 5587
rect 17604 5556 17632 5596
rect 15304 5528 17632 5556
rect 184 5466 18860 5488
rect 184 5414 1556 5466
rect 1608 5414 1620 5466
rect 1672 5414 1684 5466
rect 1736 5414 1748 5466
rect 1800 5414 1812 5466
rect 1864 5414 4656 5466
rect 4708 5414 4720 5466
rect 4772 5414 4784 5466
rect 4836 5414 4848 5466
rect 4900 5414 4912 5466
rect 4964 5414 7756 5466
rect 7808 5414 7820 5466
rect 7872 5414 7884 5466
rect 7936 5414 7948 5466
rect 8000 5414 8012 5466
rect 8064 5414 10856 5466
rect 10908 5414 10920 5466
rect 10972 5414 10984 5466
rect 11036 5414 11048 5466
rect 11100 5414 11112 5466
rect 11164 5414 13956 5466
rect 14008 5414 14020 5466
rect 14072 5414 14084 5466
rect 14136 5414 14148 5466
rect 14200 5414 14212 5466
rect 14264 5414 17056 5466
rect 17108 5414 17120 5466
rect 17172 5414 17184 5466
rect 17236 5414 17248 5466
rect 17300 5414 17312 5466
rect 17364 5414 18860 5466
rect 184 5392 18860 5414
rect 5810 5352 5816 5364
rect 3804 5324 5816 5352
rect 1673 5219 1731 5225
rect 1673 5185 1685 5219
rect 1719 5216 1731 5219
rect 1946 5216 1952 5228
rect 1719 5188 1952 5216
rect 1719 5185 1731 5188
rect 1673 5179 1731 5185
rect 1946 5176 1952 5188
rect 2004 5176 2010 5228
rect 2038 5148 2044 5160
rect 1999 5120 2044 5148
rect 2038 5108 2044 5120
rect 2096 5108 2102 5160
rect 3050 5040 3056 5092
rect 3108 5080 3114 5092
rect 3804 5080 3832 5324
rect 5810 5312 5816 5324
rect 5868 5312 5874 5364
rect 11149 5355 11207 5361
rect 11149 5321 11161 5355
rect 11195 5352 11207 5355
rect 11330 5352 11336 5364
rect 11195 5324 11336 5352
rect 11195 5321 11207 5324
rect 11149 5315 11207 5321
rect 11330 5312 11336 5324
rect 11388 5312 11394 5364
rect 15654 5312 15660 5364
rect 15712 5352 15718 5364
rect 17586 5352 17592 5364
rect 15712 5324 17592 5352
rect 15712 5312 15718 5324
rect 17586 5312 17592 5324
rect 17644 5352 17650 5364
rect 17865 5355 17923 5361
rect 17865 5352 17877 5355
rect 17644 5324 17877 5352
rect 17644 5312 17650 5324
rect 17865 5321 17877 5324
rect 17911 5321 17923 5355
rect 17865 5315 17923 5321
rect 12253 5287 12311 5293
rect 12253 5253 12265 5287
rect 12299 5284 12311 5287
rect 12434 5284 12440 5296
rect 12299 5256 12440 5284
rect 12299 5253 12311 5256
rect 12253 5247 12311 5253
rect 12434 5244 12440 5256
rect 12492 5284 12498 5296
rect 12621 5287 12679 5293
rect 12621 5284 12633 5287
rect 12492 5256 12633 5284
rect 12492 5244 12498 5256
rect 12621 5253 12633 5256
rect 12667 5284 12679 5287
rect 12667 5256 13216 5284
rect 12667 5253 12679 5256
rect 12621 5247 12679 5253
rect 4249 5219 4307 5225
rect 4249 5185 4261 5219
rect 4295 5216 4307 5219
rect 6365 5219 6423 5225
rect 6365 5216 6377 5219
rect 4295 5188 6377 5216
rect 4295 5185 4307 5188
rect 4249 5179 4307 5185
rect 6365 5185 6377 5188
rect 6411 5216 6423 5219
rect 7650 5216 7656 5228
rect 6411 5188 7656 5216
rect 6411 5185 6423 5188
rect 6365 5179 6423 5185
rect 7650 5176 7656 5188
rect 7708 5176 7714 5228
rect 8110 5176 8116 5228
rect 8168 5216 8174 5228
rect 8389 5219 8447 5225
rect 8389 5216 8401 5219
rect 8168 5188 8401 5216
rect 8168 5176 8174 5188
rect 8389 5185 8401 5188
rect 8435 5216 8447 5219
rect 9122 5216 9128 5228
rect 8435 5188 9128 5216
rect 8435 5185 8447 5188
rect 8389 5179 8447 5185
rect 9122 5176 9128 5188
rect 9180 5176 9186 5228
rect 11793 5219 11851 5225
rect 11793 5185 11805 5219
rect 11839 5216 11851 5219
rect 12710 5216 12716 5228
rect 11839 5188 12716 5216
rect 11839 5185 11851 5188
rect 11793 5179 11851 5185
rect 12710 5176 12716 5188
rect 12768 5176 12774 5228
rect 13188 5225 13216 5256
rect 13173 5219 13231 5225
rect 13173 5185 13185 5219
rect 13219 5216 13231 5219
rect 13262 5216 13268 5228
rect 13219 5188 13268 5216
rect 13219 5185 13231 5188
rect 13173 5179 13231 5185
rect 13262 5176 13268 5188
rect 13320 5216 13326 5228
rect 16117 5219 16175 5225
rect 13320 5188 14964 5216
rect 13320 5176 13326 5188
rect 10042 5108 10048 5160
rect 10100 5148 10106 5160
rect 10413 5151 10471 5157
rect 10413 5148 10425 5151
rect 10100 5120 10425 5148
rect 10100 5108 10106 5120
rect 10413 5117 10425 5120
rect 10459 5148 10471 5151
rect 13538 5148 13544 5160
rect 10459 5120 13544 5148
rect 10459 5117 10471 5120
rect 10413 5111 10471 5117
rect 13538 5108 13544 5120
rect 13596 5108 13602 5160
rect 14936 5148 14964 5188
rect 16117 5185 16129 5219
rect 16163 5216 16175 5219
rect 16390 5216 16396 5228
rect 16163 5188 16396 5216
rect 16163 5185 16175 5188
rect 16117 5179 16175 5185
rect 16390 5176 16396 5188
rect 16448 5176 16454 5228
rect 16022 5148 16028 5160
rect 14936 5134 16028 5148
rect 14950 5120 16028 5134
rect 16022 5108 16028 5120
rect 16080 5108 16086 5160
rect 17494 5108 17500 5160
rect 17552 5108 17558 5160
rect 4522 5080 4528 5092
rect 3108 5052 3832 5080
rect 4483 5052 4528 5080
rect 3108 5040 3114 5052
rect 4522 5040 4528 5052
rect 4580 5040 4586 5092
rect 5810 5080 5816 5092
rect 5750 5052 5816 5080
rect 5810 5040 5816 5052
rect 5868 5080 5874 5092
rect 6638 5080 6644 5092
rect 5868 5052 6132 5080
rect 6599 5052 6644 5080
rect 5868 5040 5874 5052
rect 3467 5015 3525 5021
rect 3467 4981 3479 5015
rect 3513 5012 3525 5015
rect 3970 5012 3976 5024
rect 3513 4984 3976 5012
rect 3513 4981 3525 4984
rect 3467 4975 3525 4981
rect 3970 4972 3976 4984
rect 4028 4972 4034 5024
rect 5166 4972 5172 5024
rect 5224 5012 5230 5024
rect 5997 5015 6055 5021
rect 5997 5012 6009 5015
rect 5224 4984 6009 5012
rect 5224 4972 5230 4984
rect 5997 4981 6009 4984
rect 6043 4981 6055 5015
rect 6104 5012 6132 5052
rect 6638 5040 6644 5052
rect 6696 5040 6702 5092
rect 8478 5080 8484 5092
rect 7866 5052 8484 5080
rect 7944 5012 7972 5052
rect 8478 5040 8484 5052
rect 8536 5040 8542 5092
rect 11514 5080 11520 5092
rect 11475 5052 11520 5080
rect 11514 5040 11520 5052
rect 11572 5040 11578 5092
rect 13814 5080 13820 5092
rect 13775 5052 13820 5080
rect 13814 5040 13820 5052
rect 13872 5040 13878 5092
rect 15565 5083 15623 5089
rect 15565 5049 15577 5083
rect 15611 5080 15623 5083
rect 15838 5080 15844 5092
rect 15611 5052 15844 5080
rect 15611 5049 15623 5052
rect 15565 5043 15623 5049
rect 15838 5040 15844 5052
rect 15896 5040 15902 5092
rect 16393 5083 16451 5089
rect 16393 5049 16405 5083
rect 16439 5080 16451 5083
rect 16666 5080 16672 5092
rect 16439 5052 16672 5080
rect 16439 5049 16451 5052
rect 16393 5043 16451 5049
rect 16666 5040 16672 5052
rect 16724 5040 16730 5092
rect 6104 4984 7972 5012
rect 5997 4975 6055 4981
rect 9950 4972 9956 5024
rect 10008 5012 10014 5024
rect 10137 5015 10195 5021
rect 10137 5012 10149 5015
rect 10008 4984 10149 5012
rect 10008 4972 10014 4984
rect 10137 4981 10149 4984
rect 10183 4981 10195 5015
rect 10137 4975 10195 4981
rect 11609 5015 11667 5021
rect 11609 4981 11621 5015
rect 11655 5012 11667 5015
rect 11882 5012 11888 5024
rect 11655 4984 11888 5012
rect 11655 4981 11667 4984
rect 11609 4975 11667 4981
rect 11882 4972 11888 4984
rect 11940 4972 11946 5024
rect 184 4922 18920 4944
rect 184 4870 3106 4922
rect 3158 4870 3170 4922
rect 3222 4870 3234 4922
rect 3286 4870 3298 4922
rect 3350 4870 3362 4922
rect 3414 4870 6206 4922
rect 6258 4870 6270 4922
rect 6322 4870 6334 4922
rect 6386 4870 6398 4922
rect 6450 4870 6462 4922
rect 6514 4870 9306 4922
rect 9358 4870 9370 4922
rect 9422 4870 9434 4922
rect 9486 4870 9498 4922
rect 9550 4870 9562 4922
rect 9614 4870 12406 4922
rect 12458 4870 12470 4922
rect 12522 4870 12534 4922
rect 12586 4870 12598 4922
rect 12650 4870 12662 4922
rect 12714 4870 15506 4922
rect 15558 4870 15570 4922
rect 15622 4870 15634 4922
rect 15686 4870 15698 4922
rect 15750 4870 15762 4922
rect 15814 4870 18606 4922
rect 18658 4870 18670 4922
rect 18722 4870 18734 4922
rect 18786 4870 18798 4922
rect 18850 4870 18862 4922
rect 18914 4870 18920 4922
rect 184 4848 18920 4870
rect 4522 4808 4528 4820
rect 4483 4780 4528 4808
rect 4522 4768 4528 4780
rect 4580 4768 4586 4820
rect 6549 4811 6607 4817
rect 6549 4777 6561 4811
rect 6595 4808 6607 4811
rect 6638 4808 6644 4820
rect 6595 4780 6644 4808
rect 6595 4777 6607 4780
rect 6549 4771 6607 4777
rect 6638 4768 6644 4780
rect 6696 4768 6702 4820
rect 13814 4768 13820 4820
rect 13872 4808 13878 4820
rect 14737 4811 14795 4817
rect 14737 4808 14749 4811
rect 13872 4780 14749 4808
rect 13872 4768 13878 4780
rect 14737 4777 14749 4780
rect 14783 4777 14795 4811
rect 16022 4808 16028 4820
rect 15935 4780 16028 4808
rect 14737 4771 14795 4777
rect 16022 4768 16028 4780
rect 16080 4808 16086 4820
rect 17494 4808 17500 4820
rect 16080 4780 17500 4808
rect 16080 4768 16086 4780
rect 17494 4768 17500 4780
rect 17552 4768 17558 4820
rect 2130 4740 2136 4752
rect 2043 4712 2136 4740
rect 2130 4700 2136 4712
rect 2188 4740 2194 4752
rect 2958 4740 2964 4752
rect 2188 4712 2964 4740
rect 2188 4700 2194 4712
rect 2958 4700 2964 4712
rect 3016 4700 3022 4752
rect 4246 4740 4252 4752
rect 3344 4712 4252 4740
rect 566 4672 572 4684
rect 527 4644 572 4672
rect 566 4632 572 4644
rect 624 4632 630 4684
rect 3344 4681 3372 4712
rect 4246 4700 4252 4712
rect 4304 4700 4310 4752
rect 12066 4740 12072 4752
rect 11362 4712 12072 4740
rect 12066 4700 12072 4712
rect 12124 4700 12130 4752
rect 13262 4700 13268 4752
rect 13320 4700 13326 4752
rect 13538 4700 13544 4752
rect 13596 4740 13602 4752
rect 16390 4740 16396 4752
rect 13596 4712 16396 4740
rect 13596 4700 13602 4712
rect 3329 4675 3387 4681
rect 3329 4641 3341 4675
rect 3375 4641 3387 4675
rect 3329 4635 3387 4641
rect 3421 4675 3479 4681
rect 3421 4641 3433 4675
rect 3467 4641 3479 4675
rect 3421 4635 3479 4641
rect 842 4604 848 4616
rect 803 4576 848 4604
rect 842 4564 848 4576
rect 900 4564 906 4616
rect 2317 4607 2375 4613
rect 2317 4573 2329 4607
rect 2363 4604 2375 4607
rect 2774 4604 2780 4616
rect 2363 4576 2780 4604
rect 2363 4573 2375 4576
rect 2317 4567 2375 4573
rect 2774 4564 2780 4576
rect 2832 4604 2838 4616
rect 3436 4604 3464 4635
rect 3510 4632 3516 4684
rect 3568 4672 3574 4684
rect 4801 4675 4859 4681
rect 3568 4644 3613 4672
rect 3568 4632 3574 4644
rect 4801 4641 4813 4675
rect 4847 4672 4859 4675
rect 5258 4672 5264 4684
rect 4847 4644 5264 4672
rect 4847 4641 4859 4644
rect 4801 4635 4859 4641
rect 5258 4632 5264 4644
rect 5316 4632 5322 4684
rect 6825 4675 6883 4681
rect 6825 4641 6837 4675
rect 6871 4672 6883 4675
rect 7282 4672 7288 4684
rect 6871 4644 7288 4672
rect 6871 4641 6883 4644
rect 6825 4635 6883 4641
rect 7282 4632 7288 4644
rect 7340 4632 7346 4684
rect 9950 4672 9956 4684
rect 9911 4644 9956 4672
rect 9950 4632 9956 4644
rect 10008 4632 10014 4684
rect 14108 4681 14136 4712
rect 16390 4700 16396 4712
rect 16448 4700 16454 4752
rect 14093 4675 14151 4681
rect 14093 4641 14105 4675
rect 14139 4641 14151 4675
rect 14918 4672 14924 4684
rect 14879 4644 14924 4672
rect 14093 4635 14151 4641
rect 14918 4632 14924 4644
rect 14976 4632 14982 4684
rect 15013 4675 15071 4681
rect 15013 4641 15025 4675
rect 15059 4672 15071 4675
rect 15378 4672 15384 4684
rect 15059 4644 15384 4672
rect 15059 4641 15071 4644
rect 15013 4635 15071 4641
rect 15378 4632 15384 4644
rect 15436 4632 15442 4684
rect 4522 4604 4528 4616
rect 2832 4576 3464 4604
rect 4483 4576 4528 4604
rect 2832 4564 2838 4576
rect 4522 4564 4528 4576
rect 4580 4564 4586 4616
rect 4709 4607 4767 4613
rect 4709 4573 4721 4607
rect 4755 4604 4767 4607
rect 5074 4604 5080 4616
rect 4755 4576 5080 4604
rect 4755 4573 4767 4576
rect 4709 4567 4767 4573
rect 5074 4564 5080 4576
rect 5132 4564 5138 4616
rect 6549 4607 6607 4613
rect 6549 4573 6561 4607
rect 6595 4604 6607 4607
rect 6730 4604 6736 4616
rect 6595 4576 6736 4604
rect 6595 4573 6607 4576
rect 6549 4567 6607 4573
rect 6730 4564 6736 4576
rect 6788 4564 6794 4616
rect 10321 4607 10379 4613
rect 10321 4573 10333 4607
rect 10367 4604 10379 4607
rect 11238 4604 11244 4616
rect 10367 4576 11244 4604
rect 10367 4573 10379 4576
rect 10321 4567 10379 4573
rect 11238 4564 11244 4576
rect 11296 4564 11302 4616
rect 13814 4604 13820 4616
rect 13775 4576 13820 4604
rect 13814 4564 13820 4576
rect 13872 4564 13878 4616
rect 14734 4604 14740 4616
rect 14695 4576 14740 4604
rect 14734 4564 14740 4576
rect 14792 4564 14798 4616
rect 3142 4468 3148 4480
rect 3103 4440 3148 4468
rect 3142 4428 3148 4440
rect 3200 4428 3206 4480
rect 6733 4471 6791 4477
rect 6733 4437 6745 4471
rect 6779 4468 6791 4471
rect 6822 4468 6828 4480
rect 6779 4440 6828 4468
rect 6779 4437 6791 4440
rect 6733 4431 6791 4437
rect 6822 4428 6828 4440
rect 6880 4428 6886 4480
rect 11606 4428 11612 4480
rect 11664 4468 11670 4480
rect 11747 4471 11805 4477
rect 11747 4468 11759 4471
rect 11664 4440 11759 4468
rect 11664 4428 11670 4440
rect 11747 4437 11759 4440
rect 11793 4437 11805 4471
rect 11747 4431 11805 4437
rect 12250 4428 12256 4480
rect 12308 4468 12314 4480
rect 12345 4471 12403 4477
rect 12345 4468 12357 4471
rect 12308 4440 12357 4468
rect 12308 4428 12314 4440
rect 12345 4437 12357 4440
rect 12391 4437 12403 4471
rect 12345 4431 12403 4437
rect 184 4378 18860 4400
rect 184 4326 1556 4378
rect 1608 4326 1620 4378
rect 1672 4326 1684 4378
rect 1736 4326 1748 4378
rect 1800 4326 1812 4378
rect 1864 4326 4656 4378
rect 4708 4326 4720 4378
rect 4772 4326 4784 4378
rect 4836 4326 4848 4378
rect 4900 4326 4912 4378
rect 4964 4326 7756 4378
rect 7808 4326 7820 4378
rect 7872 4326 7884 4378
rect 7936 4326 7948 4378
rect 8000 4326 8012 4378
rect 8064 4326 10856 4378
rect 10908 4326 10920 4378
rect 10972 4326 10984 4378
rect 11036 4326 11048 4378
rect 11100 4326 11112 4378
rect 11164 4326 13956 4378
rect 14008 4326 14020 4378
rect 14072 4326 14084 4378
rect 14136 4326 14148 4378
rect 14200 4326 14212 4378
rect 14264 4326 17056 4378
rect 17108 4326 17120 4378
rect 17172 4326 17184 4378
rect 17236 4326 17248 4378
rect 17300 4326 17312 4378
rect 17364 4326 18860 4378
rect 184 4304 18860 4326
rect 842 4224 848 4276
rect 900 4264 906 4276
rect 937 4267 995 4273
rect 937 4264 949 4267
rect 900 4236 949 4264
rect 900 4224 906 4236
rect 937 4233 949 4236
rect 983 4233 995 4267
rect 937 4227 995 4233
rect 4522 4224 4528 4276
rect 4580 4264 4586 4276
rect 4801 4267 4859 4273
rect 4801 4264 4813 4267
rect 4580 4236 4813 4264
rect 4580 4224 4586 4236
rect 4801 4233 4813 4236
rect 4847 4233 4859 4267
rect 4801 4227 4859 4233
rect 11149 4267 11207 4273
rect 11149 4233 11161 4267
rect 11195 4264 11207 4267
rect 11238 4264 11244 4276
rect 11195 4236 11244 4264
rect 11195 4233 11207 4236
rect 11149 4227 11207 4233
rect 11238 4224 11244 4236
rect 11296 4224 11302 4276
rect 14645 4267 14703 4273
rect 14645 4233 14657 4267
rect 14691 4264 14703 4267
rect 14734 4264 14740 4276
rect 14691 4236 14740 4264
rect 14691 4233 14703 4236
rect 14645 4227 14703 4233
rect 14734 4224 14740 4236
rect 14792 4224 14798 4276
rect 5074 4196 5080 4208
rect 860 4168 5080 4196
rect 860 4137 888 4168
rect 5074 4156 5080 4168
rect 5132 4156 5138 4208
rect 8202 4156 8208 4208
rect 8260 4196 8266 4208
rect 12802 4196 12808 4208
rect 8260 4168 9352 4196
rect 8260 4156 8266 4168
rect 845 4131 903 4137
rect 845 4097 857 4131
rect 891 4097 903 4131
rect 845 4091 903 4097
rect 1029 4131 1087 4137
rect 1029 4097 1041 4131
rect 1075 4128 1087 4131
rect 3142 4128 3148 4140
rect 1075 4100 3148 4128
rect 1075 4097 1087 4100
rect 1029 4091 1087 4097
rect 3142 4088 3148 4100
rect 3200 4088 3206 4140
rect 4706 4128 4712 4140
rect 4540 4100 4712 4128
rect 750 4060 756 4072
rect 711 4032 756 4060
rect 750 4020 756 4032
rect 808 4020 814 4072
rect 3510 4020 3516 4072
rect 3568 4060 3574 4072
rect 4540 4069 4568 4100
rect 4706 4088 4712 4100
rect 4764 4128 4770 4140
rect 5166 4128 5172 4140
rect 4764 4100 5172 4128
rect 4764 4088 4770 4100
rect 5166 4088 5172 4100
rect 5224 4088 5230 4140
rect 8312 4137 8340 4168
rect 9324 4137 9352 4168
rect 11808 4168 12808 4196
rect 11808 4137 11836 4168
rect 12360 4137 12388 4168
rect 12802 4156 12808 4168
rect 12860 4156 12866 4208
rect 16850 4156 16856 4208
rect 16908 4196 16914 4208
rect 17313 4199 17371 4205
rect 17313 4196 17325 4199
rect 16908 4168 17325 4196
rect 16908 4156 16914 4168
rect 17313 4165 17325 4168
rect 17359 4196 17371 4199
rect 17586 4196 17592 4208
rect 17359 4168 17592 4196
rect 17359 4165 17371 4168
rect 17313 4159 17371 4165
rect 17586 4156 17592 4168
rect 17644 4156 17650 4208
rect 8297 4131 8355 4137
rect 8297 4097 8309 4131
rect 8343 4097 8355 4131
rect 8297 4091 8355 4097
rect 9309 4131 9367 4137
rect 9309 4097 9321 4131
rect 9355 4097 9367 4131
rect 9309 4091 9367 4097
rect 11793 4131 11851 4137
rect 11793 4097 11805 4131
rect 11839 4097 11851 4131
rect 11793 4091 11851 4097
rect 12345 4131 12403 4137
rect 12345 4097 12357 4131
rect 12391 4128 12403 4131
rect 14737 4131 14795 4137
rect 12391 4100 12425 4128
rect 12391 4097 12403 4100
rect 12345 4091 12403 4097
rect 14737 4097 14749 4131
rect 14783 4128 14795 4131
rect 14826 4128 14832 4140
rect 14783 4100 14832 4128
rect 14783 4097 14795 4100
rect 14737 4091 14795 4097
rect 14826 4088 14832 4100
rect 14884 4088 14890 4140
rect 16482 4128 16488 4140
rect 16443 4100 16488 4128
rect 16482 4088 16488 4100
rect 16540 4088 16546 4140
rect 16666 4088 16672 4140
rect 16724 4128 16730 4140
rect 17037 4131 17095 4137
rect 17037 4128 17049 4131
rect 16724 4100 17049 4128
rect 16724 4088 16730 4100
rect 17037 4097 17049 4100
rect 17083 4097 17095 4131
rect 17402 4128 17408 4140
rect 17363 4100 17408 4128
rect 17037 4091 17095 4097
rect 17402 4088 17408 4100
rect 17460 4088 17466 4140
rect 4433 4063 4491 4069
rect 4433 4060 4445 4063
rect 3568 4032 4445 4060
rect 3568 4020 3574 4032
rect 4433 4029 4445 4032
rect 4479 4029 4491 4063
rect 4433 4023 4491 4029
rect 4525 4063 4583 4069
rect 4525 4029 4537 4063
rect 4571 4029 4583 4063
rect 4525 4023 4583 4029
rect 4617 4063 4675 4069
rect 4617 4029 4629 4063
rect 4663 4029 4675 4063
rect 4617 4023 4675 4029
rect 4246 3952 4252 4004
rect 4304 3992 4310 4004
rect 4632 3992 4660 4023
rect 11238 4020 11244 4072
rect 11296 4060 11302 4072
rect 11517 4063 11575 4069
rect 11517 4060 11529 4063
rect 11296 4032 11529 4060
rect 11296 4020 11302 4032
rect 11517 4029 11529 4032
rect 11563 4060 11575 4063
rect 11606 4060 11612 4072
rect 11563 4032 11612 4060
rect 11563 4029 11575 4032
rect 11517 4023 11575 4029
rect 11606 4020 11612 4032
rect 11664 4020 11670 4072
rect 14366 4020 14372 4072
rect 14424 4060 14430 4072
rect 14461 4063 14519 4069
rect 14461 4060 14473 4063
rect 14424 4032 14473 4060
rect 14424 4020 14430 4032
rect 14461 4029 14473 4032
rect 14507 4029 14519 4063
rect 14461 4023 14519 4029
rect 14553 4063 14611 4069
rect 14553 4029 14565 4063
rect 14599 4029 14611 4063
rect 14553 4023 14611 4029
rect 4304 3964 4660 3992
rect 8021 3995 8079 4001
rect 4304 3952 4310 3964
rect 8021 3961 8033 3995
rect 8067 3992 8079 3995
rect 8202 3992 8208 4004
rect 8067 3964 8208 3992
rect 8067 3961 8079 3964
rect 8021 3955 8079 3961
rect 8202 3952 8208 3964
rect 8260 3952 8266 4004
rect 9030 3952 9036 4004
rect 9088 3992 9094 4004
rect 9217 3995 9275 4001
rect 9217 3992 9229 3995
rect 9088 3964 9229 3992
rect 9088 3952 9094 3964
rect 9217 3961 9229 3964
rect 9263 3961 9275 3995
rect 9217 3955 9275 3961
rect 12529 3995 12587 4001
rect 12529 3961 12541 3995
rect 12575 3992 12587 3995
rect 12802 3992 12808 4004
rect 12575 3964 12808 3992
rect 12575 3961 12587 3964
rect 12529 3955 12587 3961
rect 12802 3952 12808 3964
rect 12860 3952 12866 4004
rect 14182 3952 14188 4004
rect 14240 3992 14246 4004
rect 14568 3992 14596 4023
rect 16206 4020 16212 4072
rect 16264 4060 16270 4072
rect 16393 4063 16451 4069
rect 16393 4060 16405 4063
rect 16264 4032 16405 4060
rect 16264 4020 16270 4032
rect 16393 4029 16405 4032
rect 16439 4029 16451 4063
rect 16500 4060 16528 4088
rect 17221 4063 17279 4069
rect 17221 4060 17233 4063
rect 16500 4032 17233 4060
rect 16393 4023 16451 4029
rect 17221 4029 17233 4032
rect 17267 4029 17279 4063
rect 17221 4023 17279 4029
rect 17494 4020 17500 4072
rect 17552 4060 17558 4072
rect 17552 4032 17597 4060
rect 17552 4020 17558 4032
rect 16301 3995 16359 4001
rect 14240 3964 16252 3992
rect 14240 3952 14246 3964
rect 7466 3884 7472 3936
rect 7524 3924 7530 3936
rect 7653 3927 7711 3933
rect 7653 3924 7665 3927
rect 7524 3896 7665 3924
rect 7524 3884 7530 3896
rect 7653 3893 7665 3896
rect 7699 3893 7711 3927
rect 7653 3887 7711 3893
rect 8113 3927 8171 3933
rect 8113 3893 8125 3927
rect 8159 3924 8171 3927
rect 8478 3924 8484 3936
rect 8159 3896 8484 3924
rect 8159 3893 8171 3896
rect 8113 3887 8171 3893
rect 8478 3884 8484 3896
rect 8536 3884 8542 3936
rect 8754 3924 8760 3936
rect 8715 3896 8760 3924
rect 8754 3884 8760 3896
rect 8812 3884 8818 3936
rect 9122 3924 9128 3936
rect 9083 3896 9128 3924
rect 9122 3884 9128 3896
rect 9180 3884 9186 3936
rect 11606 3884 11612 3936
rect 11664 3924 11670 3936
rect 11664 3896 11709 3924
rect 11664 3884 11670 3896
rect 12250 3884 12256 3936
rect 12308 3924 12314 3936
rect 12621 3927 12679 3933
rect 12621 3924 12633 3927
rect 12308 3896 12633 3924
rect 12308 3884 12314 3896
rect 12621 3893 12633 3896
rect 12667 3893 12679 3927
rect 12621 3887 12679 3893
rect 12989 3927 13047 3933
rect 12989 3893 13001 3927
rect 13035 3924 13047 3927
rect 13814 3924 13820 3936
rect 13035 3896 13820 3924
rect 13035 3893 13047 3896
rect 12989 3887 13047 3893
rect 13814 3884 13820 3896
rect 13872 3884 13878 3936
rect 15933 3927 15991 3933
rect 15933 3893 15945 3927
rect 15979 3924 15991 3927
rect 16114 3924 16120 3936
rect 15979 3896 16120 3924
rect 15979 3893 15991 3896
rect 15933 3887 15991 3893
rect 16114 3884 16120 3896
rect 16172 3884 16178 3936
rect 16224 3924 16252 3964
rect 16301 3961 16313 3995
rect 16347 3992 16359 3995
rect 16666 3992 16672 4004
rect 16347 3964 16672 3992
rect 16347 3961 16359 3964
rect 16301 3955 16359 3961
rect 16666 3952 16672 3964
rect 16724 3952 16730 4004
rect 16574 3924 16580 3936
rect 16224 3896 16580 3924
rect 16574 3884 16580 3896
rect 16632 3924 16638 3936
rect 17402 3924 17408 3936
rect 16632 3896 17408 3924
rect 16632 3884 16638 3896
rect 17402 3884 17408 3896
rect 17460 3884 17466 3936
rect 184 3834 18920 3856
rect 184 3782 3106 3834
rect 3158 3782 3170 3834
rect 3222 3782 3234 3834
rect 3286 3782 3298 3834
rect 3350 3782 3362 3834
rect 3414 3782 6206 3834
rect 6258 3782 6270 3834
rect 6322 3782 6334 3834
rect 6386 3782 6398 3834
rect 6450 3782 6462 3834
rect 6514 3782 9306 3834
rect 9358 3782 9370 3834
rect 9422 3782 9434 3834
rect 9486 3782 9498 3834
rect 9550 3782 9562 3834
rect 9614 3782 12406 3834
rect 12458 3782 12470 3834
rect 12522 3782 12534 3834
rect 12586 3782 12598 3834
rect 12650 3782 12662 3834
rect 12714 3782 15506 3834
rect 15558 3782 15570 3834
rect 15622 3782 15634 3834
rect 15686 3782 15698 3834
rect 15750 3782 15762 3834
rect 15814 3782 18606 3834
rect 18658 3782 18670 3834
rect 18722 3782 18734 3834
rect 18786 3782 18798 3834
rect 18850 3782 18862 3834
rect 18914 3782 18920 3834
rect 184 3760 18920 3782
rect 1857 3723 1915 3729
rect 1857 3689 1869 3723
rect 1903 3720 1915 3723
rect 2038 3720 2044 3732
rect 1903 3692 2044 3720
rect 1903 3689 1915 3692
rect 1857 3683 1915 3689
rect 2038 3680 2044 3692
rect 2096 3680 2102 3732
rect 5258 3720 5264 3732
rect 5219 3692 5264 3720
rect 5258 3680 5264 3692
rect 5316 3680 5322 3732
rect 6086 3720 6092 3732
rect 6047 3692 6092 3720
rect 6086 3680 6092 3692
rect 6144 3680 6150 3732
rect 6457 3723 6515 3729
rect 6457 3689 6469 3723
rect 6503 3720 6515 3723
rect 6546 3720 6552 3732
rect 6503 3692 6552 3720
rect 6503 3689 6515 3692
rect 6457 3683 6515 3689
rect 6546 3680 6552 3692
rect 6604 3680 6610 3732
rect 8478 3720 8484 3732
rect 8439 3692 8484 3720
rect 8478 3680 8484 3692
rect 8536 3680 8542 3732
rect 14182 3720 14188 3732
rect 14143 3692 14188 3720
rect 14182 3680 14188 3692
rect 14240 3680 14246 3732
rect 14550 3680 14556 3732
rect 14608 3720 14614 3732
rect 14737 3723 14795 3729
rect 14737 3720 14749 3723
rect 14608 3692 14749 3720
rect 14608 3680 14614 3692
rect 14737 3689 14749 3692
rect 14783 3689 14795 3723
rect 16298 3720 16304 3732
rect 16259 3692 16304 3720
rect 14737 3683 14795 3689
rect 16298 3680 16304 3692
rect 16356 3680 16362 3732
rect 16574 3720 16580 3732
rect 16408 3692 16580 3720
rect 1673 3655 1731 3661
rect 1673 3621 1685 3655
rect 1719 3652 1731 3655
rect 3145 3655 3203 3661
rect 3145 3652 3157 3655
rect 1719 3624 3157 3652
rect 1719 3621 1731 3624
rect 1673 3615 1731 3621
rect 3145 3621 3157 3624
rect 3191 3621 3203 3655
rect 4246 3652 4252 3664
rect 3145 3615 3203 3621
rect 3436 3624 4252 3652
rect 1394 3544 1400 3596
rect 1452 3584 1458 3596
rect 3436 3593 3464 3624
rect 1581 3587 1639 3593
rect 1581 3584 1593 3587
rect 1452 3556 1593 3584
rect 1452 3544 1458 3556
rect 1581 3553 1593 3556
rect 1627 3553 1639 3587
rect 1581 3547 1639 3553
rect 2133 3587 2191 3593
rect 2133 3553 2145 3587
rect 2179 3584 2191 3587
rect 3420 3587 3478 3593
rect 2179 3556 2774 3584
rect 2179 3553 2191 3556
rect 2133 3547 2191 3553
rect 2746 3516 2774 3556
rect 3420 3553 3432 3587
rect 3466 3553 3478 3587
rect 3420 3547 3478 3553
rect 3510 3544 3516 3596
rect 3568 3584 3574 3596
rect 3804 3593 3832 3624
rect 4246 3612 4252 3624
rect 4304 3612 4310 3664
rect 6104 3652 6132 3680
rect 6638 3652 6644 3664
rect 6104 3624 6644 3652
rect 6638 3612 6644 3624
rect 6696 3652 6702 3664
rect 6917 3655 6975 3661
rect 6917 3652 6929 3655
rect 6696 3624 6929 3652
rect 6696 3612 6702 3624
rect 6917 3621 6929 3624
rect 6963 3621 6975 3655
rect 14366 3652 14372 3664
rect 6917 3615 6975 3621
rect 13740 3624 14372 3652
rect 3789 3587 3847 3593
rect 3568 3556 3613 3584
rect 3568 3544 3574 3556
rect 3789 3553 3801 3587
rect 3835 3553 3847 3587
rect 3970 3584 3976 3596
rect 3931 3556 3976 3584
rect 3789 3547 3847 3553
rect 3970 3544 3976 3556
rect 4028 3544 4034 3596
rect 4982 3544 4988 3596
rect 5040 3584 5046 3596
rect 5169 3587 5227 3593
rect 5169 3584 5181 3587
rect 5040 3556 5181 3584
rect 5040 3544 5046 3556
rect 5169 3553 5181 3556
rect 5215 3553 5227 3587
rect 6822 3584 6828 3596
rect 6783 3556 6828 3584
rect 5169 3547 5227 3553
rect 6822 3544 6828 3556
rect 6880 3544 6886 3596
rect 11238 3584 11244 3596
rect 11199 3556 11244 3584
rect 11238 3544 11244 3556
rect 11296 3544 11302 3596
rect 11330 3544 11336 3596
rect 11388 3584 11394 3596
rect 11425 3587 11483 3593
rect 11425 3584 11437 3587
rect 11388 3556 11437 3584
rect 11388 3544 11394 3556
rect 11425 3553 11437 3556
rect 11471 3584 11483 3587
rect 12250 3584 12256 3596
rect 11471 3556 12256 3584
rect 11471 3553 11483 3556
rect 11425 3547 11483 3553
rect 12250 3544 12256 3556
rect 12308 3544 12314 3596
rect 13740 3593 13768 3624
rect 14366 3612 14372 3624
rect 14424 3652 14430 3664
rect 14568 3652 14596 3680
rect 14424 3624 14596 3652
rect 14424 3612 14430 3624
rect 13725 3587 13783 3593
rect 13725 3553 13737 3587
rect 13771 3553 13783 3587
rect 13725 3547 13783 3553
rect 14001 3587 14059 3593
rect 14001 3553 14013 3587
rect 14047 3584 14059 3587
rect 14458 3584 14464 3596
rect 14047 3556 14464 3584
rect 14047 3553 14059 3556
rect 14001 3547 14059 3553
rect 14458 3544 14464 3556
rect 14516 3584 14522 3596
rect 15102 3584 15108 3596
rect 14516 3556 15108 3584
rect 14516 3544 14522 3556
rect 15102 3544 15108 3556
rect 15160 3544 15166 3596
rect 16114 3584 16120 3596
rect 16075 3556 16120 3584
rect 16114 3544 16120 3556
rect 16172 3544 16178 3596
rect 16408 3593 16436 3692
rect 16574 3680 16580 3692
rect 16632 3680 16638 3732
rect 17405 3723 17463 3729
rect 17405 3689 17417 3723
rect 17451 3720 17463 3723
rect 17494 3720 17500 3732
rect 17451 3692 17500 3720
rect 17451 3689 17463 3692
rect 17405 3683 17463 3689
rect 17494 3680 17500 3692
rect 17552 3680 17558 3732
rect 18138 3680 18144 3732
rect 18196 3720 18202 3732
rect 18233 3723 18291 3729
rect 18233 3720 18245 3723
rect 18196 3692 18245 3720
rect 18196 3680 18202 3692
rect 18233 3689 18245 3692
rect 18279 3689 18291 3723
rect 18233 3683 18291 3689
rect 16592 3624 17724 3652
rect 16393 3587 16451 3593
rect 16393 3553 16405 3587
rect 16439 3553 16451 3587
rect 16393 3547 16451 3553
rect 16482 3544 16488 3596
rect 16540 3584 16546 3596
rect 16592 3593 16620 3624
rect 16577 3587 16635 3593
rect 16577 3584 16589 3587
rect 16540 3556 16589 3584
rect 16540 3544 16546 3556
rect 16577 3553 16589 3556
rect 16623 3553 16635 3587
rect 16577 3547 16635 3553
rect 17402 3544 17408 3596
rect 17460 3584 17466 3596
rect 17696 3593 17724 3624
rect 17497 3587 17555 3593
rect 17497 3584 17509 3587
rect 17460 3556 17509 3584
rect 17460 3544 17466 3556
rect 17497 3553 17509 3556
rect 17543 3553 17555 3587
rect 17497 3547 17555 3553
rect 17681 3587 17739 3593
rect 17681 3553 17693 3587
rect 17727 3553 17739 3587
rect 18414 3584 18420 3596
rect 18327 3556 18420 3584
rect 17681 3547 17739 3553
rect 18414 3544 18420 3556
rect 18472 3584 18478 3596
rect 19058 3584 19064 3596
rect 18472 3556 19064 3584
rect 18472 3544 18478 3556
rect 19058 3544 19064 3556
rect 19116 3544 19122 3596
rect 3881 3519 3939 3525
rect 3881 3516 3893 3519
rect 2746 3488 3893 3516
rect 3881 3485 3893 3488
rect 3927 3485 3939 3519
rect 3881 3479 3939 3485
rect 7009 3519 7067 3525
rect 7009 3485 7021 3519
rect 7055 3485 7067 3519
rect 7009 3479 7067 3485
rect 7024 3448 7052 3479
rect 3528 3420 7052 3448
rect 3528 3392 3556 3420
rect 10778 3408 10784 3460
rect 10836 3448 10842 3460
rect 11425 3451 11483 3457
rect 11425 3448 11437 3451
rect 10836 3420 11437 3448
rect 10836 3408 10842 3420
rect 11425 3417 11437 3420
rect 11471 3417 11483 3451
rect 11425 3411 11483 3417
rect 13817 3451 13875 3457
rect 13817 3417 13829 3451
rect 13863 3448 13875 3451
rect 16206 3448 16212 3460
rect 13863 3420 16212 3448
rect 13863 3417 13875 3420
rect 13817 3411 13875 3417
rect 16206 3408 16212 3420
rect 16264 3408 16270 3460
rect 2041 3383 2099 3389
rect 2041 3349 2053 3383
rect 2087 3380 2099 3383
rect 2130 3380 2136 3392
rect 2087 3352 2136 3380
rect 2087 3349 2099 3352
rect 2041 3343 2099 3349
rect 2130 3340 2136 3352
rect 2188 3380 2194 3392
rect 3510 3380 3516 3392
rect 2188 3352 3516 3380
rect 2188 3340 2194 3352
rect 3510 3340 3516 3352
rect 3568 3340 3574 3392
rect 16942 3340 16948 3392
rect 17000 3380 17006 3392
rect 17221 3383 17279 3389
rect 17221 3380 17233 3383
rect 17000 3352 17233 3380
rect 17000 3340 17006 3352
rect 17221 3349 17233 3352
rect 17267 3349 17279 3383
rect 17221 3343 17279 3349
rect 184 3290 18860 3312
rect 184 3238 1556 3290
rect 1608 3238 1620 3290
rect 1672 3238 1684 3290
rect 1736 3238 1748 3290
rect 1800 3238 1812 3290
rect 1864 3238 4656 3290
rect 4708 3238 4720 3290
rect 4772 3238 4784 3290
rect 4836 3238 4848 3290
rect 4900 3238 4912 3290
rect 4964 3238 7756 3290
rect 7808 3238 7820 3290
rect 7872 3238 7884 3290
rect 7936 3238 7948 3290
rect 8000 3238 8012 3290
rect 8064 3238 10856 3290
rect 10908 3238 10920 3290
rect 10972 3238 10984 3290
rect 11036 3238 11048 3290
rect 11100 3238 11112 3290
rect 11164 3238 13956 3290
rect 14008 3238 14020 3290
rect 14072 3238 14084 3290
rect 14136 3238 14148 3290
rect 14200 3238 14212 3290
rect 14264 3238 17056 3290
rect 17108 3238 17120 3290
rect 17172 3238 17184 3290
rect 17236 3238 17248 3290
rect 17300 3238 17312 3290
rect 17364 3238 18860 3290
rect 184 3216 18860 3238
rect 750 3136 756 3188
rect 808 3176 814 3188
rect 845 3179 903 3185
rect 845 3176 857 3179
rect 808 3148 857 3176
rect 808 3136 814 3148
rect 845 3145 857 3148
rect 891 3145 903 3179
rect 4982 3176 4988 3188
rect 4943 3148 4988 3176
rect 845 3139 903 3145
rect 4982 3136 4988 3148
rect 5040 3136 5046 3188
rect 6638 3176 6644 3188
rect 6599 3148 6644 3176
rect 6638 3136 6644 3148
rect 6696 3136 6702 3188
rect 6822 3136 6828 3188
rect 6880 3176 6886 3188
rect 6917 3179 6975 3185
rect 6917 3176 6929 3179
rect 6880 3148 6929 3176
rect 6880 3136 6886 3148
rect 6917 3145 6929 3148
rect 6963 3145 6975 3179
rect 6917 3139 6975 3145
rect 8757 3179 8815 3185
rect 8757 3145 8769 3179
rect 8803 3176 8815 3179
rect 9122 3176 9128 3188
rect 8803 3148 9128 3176
rect 8803 3145 8815 3148
rect 8757 3139 8815 3145
rect 9122 3136 9128 3148
rect 9180 3136 9186 3188
rect 11514 3176 11520 3188
rect 11475 3148 11520 3176
rect 11514 3136 11520 3148
rect 11572 3176 11578 3188
rect 11790 3176 11796 3188
rect 11572 3148 11796 3176
rect 11572 3136 11578 3148
rect 11790 3136 11796 3148
rect 11848 3136 11854 3188
rect 12437 3179 12495 3185
rect 12437 3145 12449 3179
rect 12483 3176 12495 3179
rect 12802 3176 12808 3188
rect 12483 3148 12808 3176
rect 12483 3145 12495 3148
rect 12437 3139 12495 3145
rect 12802 3136 12808 3148
rect 12860 3136 12866 3188
rect 14826 3176 14832 3188
rect 14787 3148 14832 3176
rect 14826 3136 14832 3148
rect 14884 3136 14890 3188
rect 16942 3136 16948 3188
rect 17000 3176 17006 3188
rect 17129 3179 17187 3185
rect 17129 3176 17141 3179
rect 17000 3148 17141 3176
rect 17000 3136 17006 3148
rect 17129 3145 17141 3148
rect 17175 3145 17187 3179
rect 18414 3176 18420 3188
rect 18375 3148 18420 3176
rect 17129 3139 17187 3145
rect 18414 3136 18420 3148
rect 18472 3136 18478 3188
rect 10321 3111 10379 3117
rect 10321 3077 10333 3111
rect 10367 3108 10379 3111
rect 10367 3080 12434 3108
rect 10367 3077 10379 3080
rect 10321 3071 10379 3077
rect 5629 3043 5687 3049
rect 5629 3009 5641 3043
rect 5675 3040 5687 3043
rect 5902 3040 5908 3052
rect 5675 3012 5908 3040
rect 5675 3009 5687 3012
rect 5629 3003 5687 3009
rect 5902 3000 5908 3012
rect 5960 3000 5966 3052
rect 6638 3000 6644 3052
rect 6696 3040 6702 3052
rect 7377 3043 7435 3049
rect 7377 3040 7389 3043
rect 6696 3012 7389 3040
rect 6696 3000 6702 3012
rect 7377 3009 7389 3012
rect 7423 3009 7435 3043
rect 7558 3040 7564 3052
rect 7471 3012 7564 3040
rect 7377 3003 7435 3009
rect 7558 3000 7564 3012
rect 7616 3040 7622 3052
rect 9309 3043 9367 3049
rect 9309 3040 9321 3043
rect 7616 3012 9321 3040
rect 7616 3000 7622 3012
rect 9309 3009 9321 3012
rect 9355 3009 9367 3043
rect 11149 3043 11207 3049
rect 11149 3040 11161 3043
rect 9309 3003 9367 3009
rect 10520 3012 11161 3040
rect 750 2972 756 2984
rect 711 2944 756 2972
rect 750 2932 756 2944
rect 808 2932 814 2984
rect 7282 2972 7288 2984
rect 7243 2944 7288 2972
rect 7282 2932 7288 2944
rect 7340 2932 7346 2984
rect 9030 2932 9036 2984
rect 9088 2972 9094 2984
rect 10520 2981 10548 3012
rect 11149 3009 11161 3012
rect 11195 3009 11207 3043
rect 11149 3003 11207 3009
rect 11238 3000 11244 3052
rect 11296 3040 11302 3052
rect 11422 3040 11428 3052
rect 11296 3012 11428 3040
rect 11296 3000 11302 3012
rect 11422 3000 11428 3012
rect 11480 3040 11486 3052
rect 11609 3043 11667 3049
rect 11609 3040 11621 3043
rect 11480 3012 11621 3040
rect 11480 3000 11486 3012
rect 11609 3009 11621 3012
rect 11655 3009 11667 3043
rect 11609 3003 11667 3009
rect 9217 2975 9275 2981
rect 9217 2972 9229 2975
rect 9088 2944 9229 2972
rect 9088 2932 9094 2944
rect 9217 2941 9229 2944
rect 9263 2941 9275 2975
rect 9217 2935 9275 2941
rect 10505 2975 10563 2981
rect 10505 2941 10517 2975
rect 10551 2941 10563 2975
rect 10778 2972 10784 2984
rect 10739 2944 10784 2972
rect 10505 2935 10563 2941
rect 10778 2932 10784 2944
rect 10836 2932 10842 2984
rect 11330 2972 11336 2984
rect 11291 2944 11336 2972
rect 11330 2932 11336 2944
rect 11388 2932 11394 2984
rect 5445 2907 5503 2913
rect 5445 2873 5457 2907
rect 5491 2904 5503 2907
rect 5534 2904 5540 2916
rect 5491 2876 5540 2904
rect 5491 2873 5503 2876
rect 5445 2867 5503 2873
rect 5534 2864 5540 2876
rect 5592 2904 5598 2916
rect 9048 2904 9076 2932
rect 5592 2876 9076 2904
rect 10689 2907 10747 2913
rect 5592 2864 5598 2876
rect 10689 2873 10701 2907
rect 10735 2904 10747 2907
rect 12406 2904 12434 3080
rect 12802 3000 12808 3052
rect 12860 3040 12866 3052
rect 12989 3043 13047 3049
rect 12989 3040 13001 3043
rect 12860 3012 13001 3040
rect 12860 3000 12866 3012
rect 12989 3009 13001 3012
rect 13035 3040 13047 3043
rect 13170 3040 13176 3052
rect 13035 3012 13176 3040
rect 13035 3009 13047 3012
rect 12989 3003 13047 3009
rect 13170 3000 13176 3012
rect 13228 3040 13234 3052
rect 15381 3043 15439 3049
rect 15381 3040 15393 3043
rect 13228 3012 15393 3040
rect 13228 3000 13234 3012
rect 15381 3009 15393 3012
rect 15427 3040 15439 3043
rect 16482 3040 16488 3052
rect 15427 3012 16488 3040
rect 15427 3009 15439 3012
rect 15381 3003 15439 3009
rect 16482 3000 16488 3012
rect 16540 3040 16546 3052
rect 17681 3043 17739 3049
rect 17681 3040 17693 3043
rect 16540 3012 17693 3040
rect 16540 3000 16546 3012
rect 17681 3009 17693 3012
rect 17727 3009 17739 3043
rect 17681 3003 17739 3009
rect 15102 2932 15108 2984
rect 15160 2972 15166 2984
rect 15289 2975 15347 2981
rect 15289 2972 15301 2975
rect 15160 2944 15301 2972
rect 15160 2932 15166 2944
rect 15289 2941 15301 2944
rect 15335 2941 15347 2975
rect 15289 2935 15347 2941
rect 12805 2907 12863 2913
rect 12805 2904 12817 2907
rect 10735 2876 11560 2904
rect 12406 2876 12817 2904
rect 10735 2873 10747 2876
rect 10689 2867 10747 2873
rect 11532 2848 11560 2876
rect 12805 2873 12817 2876
rect 12851 2873 12863 2907
rect 12805 2867 12863 2873
rect 16853 2907 16911 2913
rect 16853 2873 16865 2907
rect 16899 2904 16911 2907
rect 17586 2904 17592 2916
rect 16899 2876 17592 2904
rect 16899 2873 16911 2876
rect 16853 2867 16911 2873
rect 17586 2864 17592 2876
rect 17644 2864 17650 2916
rect 5350 2836 5356 2848
rect 5311 2808 5356 2836
rect 5350 2796 5356 2808
rect 5408 2796 5414 2848
rect 9030 2796 9036 2848
rect 9088 2836 9094 2848
rect 9125 2839 9183 2845
rect 9125 2836 9137 2839
rect 9088 2808 9137 2836
rect 9088 2796 9094 2808
rect 9125 2805 9137 2808
rect 9171 2805 9183 2839
rect 9125 2799 9183 2805
rect 11514 2796 11520 2848
rect 11572 2796 11578 2848
rect 12897 2839 12955 2845
rect 12897 2805 12909 2839
rect 12943 2836 12955 2839
rect 13170 2836 13176 2848
rect 12943 2808 13176 2836
rect 12943 2805 12955 2808
rect 12897 2799 12955 2805
rect 13170 2796 13176 2808
rect 13228 2836 13234 2848
rect 13722 2836 13728 2848
rect 13228 2808 13728 2836
rect 13228 2796 13234 2808
rect 13722 2796 13728 2808
rect 13780 2796 13786 2848
rect 15194 2836 15200 2848
rect 15155 2808 15200 2836
rect 15194 2796 15200 2808
rect 15252 2796 15258 2848
rect 17494 2836 17500 2848
rect 17455 2808 17500 2836
rect 17494 2796 17500 2808
rect 17552 2796 17558 2848
rect 184 2746 18920 2768
rect 184 2694 3106 2746
rect 3158 2694 3170 2746
rect 3222 2694 3234 2746
rect 3286 2694 3298 2746
rect 3350 2694 3362 2746
rect 3414 2694 6206 2746
rect 6258 2694 6270 2746
rect 6322 2694 6334 2746
rect 6386 2694 6398 2746
rect 6450 2694 6462 2746
rect 6514 2694 9306 2746
rect 9358 2694 9370 2746
rect 9422 2694 9434 2746
rect 9486 2694 9498 2746
rect 9550 2694 9562 2746
rect 9614 2694 12406 2746
rect 12458 2694 12470 2746
rect 12522 2694 12534 2746
rect 12586 2694 12598 2746
rect 12650 2694 12662 2746
rect 12714 2694 15506 2746
rect 15558 2694 15570 2746
rect 15622 2694 15634 2746
rect 15686 2694 15698 2746
rect 15750 2694 15762 2746
rect 15814 2694 18606 2746
rect 18658 2694 18670 2746
rect 18722 2694 18734 2746
rect 18786 2694 18798 2746
rect 18850 2694 18862 2746
rect 18914 2694 18920 2746
rect 184 2672 18920 2694
rect 569 2635 627 2641
rect 569 2601 581 2635
rect 615 2632 627 2635
rect 750 2632 756 2644
rect 615 2604 756 2632
rect 615 2601 627 2604
rect 569 2595 627 2601
rect 750 2592 756 2604
rect 808 2592 814 2644
rect 1394 2592 1400 2644
rect 1452 2632 1458 2644
rect 1581 2635 1639 2641
rect 1581 2632 1593 2635
rect 1452 2604 1593 2632
rect 1452 2592 1458 2604
rect 1581 2601 1593 2604
rect 1627 2601 1639 2635
rect 1581 2595 1639 2601
rect 2041 2635 2099 2641
rect 2041 2601 2053 2635
rect 2087 2632 2099 2635
rect 2222 2632 2228 2644
rect 2087 2604 2228 2632
rect 2087 2601 2099 2604
rect 2041 2595 2099 2601
rect 2222 2592 2228 2604
rect 2280 2632 2286 2644
rect 2777 2635 2835 2641
rect 2777 2632 2789 2635
rect 2280 2604 2789 2632
rect 2280 2592 2286 2604
rect 2777 2601 2789 2604
rect 2823 2601 2835 2635
rect 5350 2632 5356 2644
rect 5311 2604 5356 2632
rect 2777 2595 2835 2601
rect 2792 2564 2820 2595
rect 5350 2592 5356 2604
rect 5408 2592 5414 2644
rect 5534 2592 5540 2644
rect 5592 2632 5598 2644
rect 5813 2635 5871 2641
rect 5813 2632 5825 2635
rect 5592 2604 5825 2632
rect 5592 2592 5598 2604
rect 5813 2601 5825 2604
rect 5859 2601 5871 2635
rect 8202 2632 8208 2644
rect 8163 2604 8208 2632
rect 5813 2595 5871 2601
rect 8202 2592 8208 2604
rect 8260 2592 8266 2644
rect 13173 2635 13231 2641
rect 13173 2601 13185 2635
rect 13219 2601 13231 2635
rect 13173 2595 13231 2601
rect 14277 2635 14335 2641
rect 14277 2601 14289 2635
rect 14323 2632 14335 2635
rect 14366 2632 14372 2644
rect 14323 2604 14372 2632
rect 14323 2601 14335 2604
rect 14277 2595 14335 2601
rect 4154 2564 4160 2576
rect 2792 2536 4160 2564
rect 4154 2524 4160 2536
rect 4212 2564 4218 2576
rect 7837 2567 7895 2573
rect 7837 2564 7849 2567
rect 4212 2536 7849 2564
rect 4212 2524 4218 2536
rect 7837 2533 7849 2536
rect 7883 2564 7895 2567
rect 8478 2564 8484 2576
rect 7883 2536 8484 2564
rect 7883 2533 7895 2536
rect 7837 2527 7895 2533
rect 8478 2524 8484 2536
rect 8536 2564 8542 2576
rect 8665 2567 8723 2573
rect 8665 2564 8677 2567
rect 8536 2536 8677 2564
rect 8536 2524 8542 2536
rect 8665 2533 8677 2536
rect 8711 2533 8723 2567
rect 13188 2564 13216 2595
rect 14366 2592 14372 2604
rect 14424 2592 14430 2644
rect 15194 2632 15200 2644
rect 15155 2604 15200 2632
rect 15194 2592 15200 2604
rect 15252 2592 15258 2644
rect 15378 2592 15384 2644
rect 15436 2632 15442 2644
rect 15565 2635 15623 2641
rect 15565 2632 15577 2635
rect 15436 2604 15577 2632
rect 15436 2592 15442 2604
rect 15565 2601 15577 2604
rect 15611 2601 15623 2635
rect 15565 2595 15623 2601
rect 17221 2635 17279 2641
rect 17221 2601 17233 2635
rect 17267 2632 17279 2635
rect 17494 2632 17500 2644
rect 17267 2604 17500 2632
rect 17267 2601 17279 2604
rect 17221 2595 17279 2601
rect 17494 2592 17500 2604
rect 17552 2592 17558 2644
rect 17586 2592 17592 2644
rect 17644 2632 17650 2644
rect 17681 2635 17739 2641
rect 17681 2632 17693 2635
rect 17644 2604 17693 2632
rect 17644 2592 17650 2604
rect 17681 2601 17693 2604
rect 17727 2601 17739 2635
rect 17681 2595 17739 2601
rect 13188 2536 13952 2564
rect 8665 2527 8723 2533
rect 934 2496 940 2508
rect 895 2468 940 2496
rect 934 2456 940 2468
rect 992 2456 998 2508
rect 1949 2499 2007 2505
rect 1949 2465 1961 2499
rect 1995 2496 2007 2499
rect 2866 2496 2872 2508
rect 1995 2468 2872 2496
rect 1995 2465 2007 2468
rect 1949 2459 2007 2465
rect 2866 2456 2872 2468
rect 2924 2456 2930 2508
rect 5626 2456 5632 2508
rect 5684 2496 5690 2508
rect 5721 2499 5779 2505
rect 5721 2496 5733 2499
rect 5684 2468 5733 2496
rect 5684 2456 5690 2468
rect 5721 2465 5733 2468
rect 5767 2465 5779 2499
rect 8570 2496 8576 2508
rect 8531 2468 8576 2496
rect 5721 2459 5779 2465
rect 8570 2456 8576 2468
rect 8628 2456 8634 2508
rect 13173 2499 13231 2505
rect 13173 2465 13185 2499
rect 13219 2496 13231 2499
rect 13722 2496 13728 2508
rect 13219 2468 13584 2496
rect 13683 2468 13728 2496
rect 13219 2465 13231 2468
rect 13173 2459 13231 2465
rect 1026 2428 1032 2440
rect 987 2400 1032 2428
rect 1026 2388 1032 2400
rect 1084 2388 1090 2440
rect 1213 2431 1271 2437
rect 1213 2397 1225 2431
rect 1259 2397 1271 2431
rect 1213 2391 1271 2397
rect 1228 2360 1256 2391
rect 2130 2388 2136 2440
rect 2188 2428 2194 2440
rect 2188 2400 2281 2428
rect 2188 2388 2194 2400
rect 4062 2388 4068 2440
rect 4120 2428 4126 2440
rect 5905 2431 5963 2437
rect 5905 2428 5917 2431
rect 4120 2400 5917 2428
rect 4120 2388 4126 2400
rect 5905 2397 5917 2400
rect 5951 2397 5963 2431
rect 5905 2391 5963 2397
rect 8757 2431 8815 2437
rect 8757 2397 8769 2431
rect 8803 2397 8815 2431
rect 8757 2391 8815 2397
rect 13449 2431 13507 2437
rect 13449 2397 13461 2431
rect 13495 2397 13507 2431
rect 13556 2428 13584 2468
rect 13722 2456 13728 2468
rect 13780 2456 13786 2508
rect 13924 2505 13952 2536
rect 15102 2524 15108 2576
rect 15160 2564 15166 2576
rect 15657 2567 15715 2573
rect 15657 2564 15669 2567
rect 15160 2536 15669 2564
rect 15160 2524 15166 2536
rect 15657 2533 15669 2536
rect 15703 2533 15715 2567
rect 15657 2527 15715 2533
rect 16761 2567 16819 2573
rect 16761 2533 16773 2567
rect 16807 2564 16819 2567
rect 17604 2564 17632 2592
rect 16807 2536 17632 2564
rect 16807 2533 16819 2536
rect 16761 2527 16819 2533
rect 13909 2499 13967 2505
rect 13909 2465 13921 2499
rect 13955 2465 13967 2499
rect 13909 2459 13967 2465
rect 14366 2456 14372 2508
rect 14424 2496 14430 2508
rect 16776 2496 16804 2527
rect 17586 2496 17592 2508
rect 14424 2468 16804 2496
rect 17547 2468 17592 2496
rect 14424 2456 14430 2468
rect 17586 2456 17592 2468
rect 17644 2456 17650 2508
rect 14458 2428 14464 2440
rect 13556 2400 14464 2428
rect 13449 2391 13507 2397
rect 2148 2360 2176 2388
rect 1228 2332 2176 2360
rect 7558 2320 7564 2372
rect 7616 2360 7622 2372
rect 8772 2360 8800 2391
rect 13262 2360 13268 2372
rect 7616 2332 8800 2360
rect 13223 2332 13268 2360
rect 7616 2320 7622 2332
rect 13262 2320 13268 2332
rect 13320 2320 13326 2372
rect 13464 2360 13492 2391
rect 14458 2388 14464 2400
rect 14516 2388 14522 2440
rect 15562 2388 15568 2440
rect 15620 2428 15626 2440
rect 15841 2431 15899 2437
rect 15841 2428 15853 2431
rect 15620 2400 15853 2428
rect 15620 2388 15626 2400
rect 15841 2397 15853 2400
rect 15887 2428 15899 2431
rect 16298 2428 16304 2440
rect 15887 2400 16304 2428
rect 15887 2397 15899 2400
rect 15841 2391 15899 2397
rect 16298 2388 16304 2400
rect 16356 2428 16362 2440
rect 17773 2431 17831 2437
rect 16356 2400 16574 2428
rect 16356 2388 16362 2400
rect 14366 2360 14372 2372
rect 13464 2332 14372 2360
rect 14366 2320 14372 2332
rect 14424 2320 14430 2372
rect 16546 2360 16574 2400
rect 17773 2397 17785 2431
rect 17819 2397 17831 2431
rect 17773 2391 17831 2397
rect 17788 2360 17816 2391
rect 16546 2332 17816 2360
rect 13722 2292 13728 2304
rect 13683 2264 13728 2292
rect 13722 2252 13728 2264
rect 13780 2252 13786 2304
rect 184 2202 18860 2224
rect 184 2150 1556 2202
rect 1608 2150 1620 2202
rect 1672 2150 1684 2202
rect 1736 2150 1748 2202
rect 1800 2150 1812 2202
rect 1864 2150 4656 2202
rect 4708 2150 4720 2202
rect 4772 2150 4784 2202
rect 4836 2150 4848 2202
rect 4900 2150 4912 2202
rect 4964 2150 7756 2202
rect 7808 2150 7820 2202
rect 7872 2150 7884 2202
rect 7936 2150 7948 2202
rect 8000 2150 8012 2202
rect 8064 2150 10856 2202
rect 10908 2150 10920 2202
rect 10972 2150 10984 2202
rect 11036 2150 11048 2202
rect 11100 2150 11112 2202
rect 11164 2150 13956 2202
rect 14008 2150 14020 2202
rect 14072 2150 14084 2202
rect 14136 2150 14148 2202
rect 14200 2150 14212 2202
rect 14264 2150 17056 2202
rect 17108 2150 17120 2202
rect 17172 2150 17184 2202
rect 17236 2150 17248 2202
rect 17300 2150 17312 2202
rect 17364 2150 18860 2202
rect 184 2128 18860 2150
rect 1026 2048 1032 2100
rect 1084 2088 1090 2100
rect 1581 2091 1639 2097
rect 1581 2088 1593 2091
rect 1084 2060 1593 2088
rect 1084 2048 1090 2060
rect 1581 2057 1593 2060
rect 1627 2057 1639 2091
rect 2866 2088 2872 2100
rect 2827 2060 2872 2088
rect 1581 2051 1639 2057
rect 1596 1952 1624 2051
rect 2866 2048 2872 2060
rect 2924 2048 2930 2100
rect 4065 2091 4123 2097
rect 4065 2057 4077 2091
rect 4111 2088 4123 2091
rect 4154 2088 4160 2100
rect 4111 2060 4160 2088
rect 4111 2057 4123 2060
rect 4065 2051 4123 2057
rect 4080 2020 4108 2051
rect 4154 2048 4160 2060
rect 4212 2048 4218 2100
rect 11606 2048 11612 2100
rect 11664 2088 11670 2100
rect 12161 2091 12219 2097
rect 12161 2088 12173 2091
rect 11664 2060 12173 2088
rect 11664 2048 11670 2060
rect 12161 2057 12173 2060
rect 12207 2057 12219 2091
rect 16206 2088 16212 2100
rect 12161 2051 12219 2057
rect 14844 2060 16212 2088
rect 7282 2020 7288 2032
rect 3344 1992 4108 2020
rect 7208 1992 7288 2020
rect 2866 1952 2872 1964
rect 1596 1924 2872 1952
rect 2866 1912 2872 1924
rect 2924 1912 2930 1964
rect 3344 1961 3372 1992
rect 3329 1955 3387 1961
rect 3329 1921 3341 1955
rect 3375 1921 3387 1955
rect 3329 1915 3387 1921
rect 3513 1955 3571 1961
rect 3513 1921 3525 1955
rect 3559 1952 3571 1955
rect 4062 1952 4068 1964
rect 3559 1924 4068 1952
rect 3559 1921 3571 1924
rect 3513 1915 3571 1921
rect 4062 1912 4068 1924
rect 4120 1912 4126 1964
rect 7208 1961 7236 1992
rect 7282 1980 7288 1992
rect 7340 1980 7346 2032
rect 11882 2020 11888 2032
rect 11843 1992 11888 2020
rect 11882 1980 11888 1992
rect 11940 1980 11946 2032
rect 13722 2020 13728 2032
rect 12636 1992 13728 2020
rect 7193 1955 7251 1961
rect 7193 1921 7205 1955
rect 7239 1921 7251 1955
rect 7193 1915 7251 1921
rect 8386 1912 8392 1964
rect 8444 1952 8450 1964
rect 9217 1955 9275 1961
rect 9217 1952 9229 1955
rect 8444 1924 9229 1952
rect 8444 1912 8450 1924
rect 9217 1921 9229 1924
rect 9263 1921 9275 1955
rect 9217 1915 9275 1921
rect 11333 1955 11391 1961
rect 11333 1921 11345 1955
rect 11379 1952 11391 1955
rect 12526 1952 12532 1964
rect 11379 1924 12532 1952
rect 11379 1921 11391 1924
rect 11333 1915 11391 1921
rect 12526 1912 12532 1924
rect 12584 1912 12590 1964
rect 12636 1961 12664 1992
rect 13722 1980 13728 1992
rect 13780 1980 13786 2032
rect 12621 1955 12679 1961
rect 12621 1921 12633 1955
rect 12667 1921 12679 1955
rect 12621 1915 12679 1921
rect 12710 1912 12716 1964
rect 12768 1952 12774 1964
rect 12768 1924 12813 1952
rect 12768 1912 12774 1924
rect 13262 1912 13268 1964
rect 13320 1952 13326 1964
rect 13998 1952 14004 1964
rect 13320 1924 13768 1952
rect 13911 1924 14004 1952
rect 13320 1912 13326 1924
rect 13740 1896 13768 1924
rect 13998 1912 14004 1924
rect 14056 1952 14062 1964
rect 14458 1952 14464 1964
rect 14056 1924 14464 1952
rect 14056 1912 14062 1924
rect 14458 1912 14464 1924
rect 14516 1912 14522 1964
rect 3970 1844 3976 1896
rect 4028 1884 4034 1896
rect 4341 1887 4399 1893
rect 4341 1884 4353 1887
rect 4028 1856 4353 1884
rect 4028 1844 4034 1856
rect 4341 1853 4353 1856
rect 4387 1853 4399 1887
rect 4341 1847 4399 1853
rect 4522 1844 4528 1896
rect 4580 1884 4586 1896
rect 4617 1887 4675 1893
rect 4617 1884 4629 1887
rect 4580 1856 4629 1884
rect 4580 1844 4586 1856
rect 4617 1853 4629 1856
rect 4663 1853 4675 1887
rect 5166 1884 5172 1896
rect 5127 1856 5172 1884
rect 4617 1847 4675 1853
rect 5166 1844 5172 1856
rect 5224 1844 5230 1896
rect 7377 1887 7435 1893
rect 7377 1853 7389 1887
rect 7423 1853 7435 1887
rect 7377 1847 7435 1853
rect 7653 1887 7711 1893
rect 7653 1853 7665 1887
rect 7699 1884 7711 1887
rect 8662 1884 8668 1896
rect 7699 1856 8668 1884
rect 7699 1853 7711 1856
rect 7653 1847 7711 1853
rect 7392 1816 7420 1847
rect 8662 1844 8668 1856
rect 8720 1844 8726 1896
rect 9585 1887 9643 1893
rect 9585 1853 9597 1887
rect 9631 1884 9643 1887
rect 9631 1856 13676 1884
rect 9631 1853 9643 1856
rect 9585 1847 9643 1853
rect 9122 1816 9128 1828
rect 7392 1788 9128 1816
rect 9122 1776 9128 1788
rect 9180 1776 9186 1828
rect 11425 1819 11483 1825
rect 11425 1785 11437 1819
rect 11471 1816 11483 1819
rect 13648 1816 13676 1856
rect 13722 1844 13728 1896
rect 13780 1884 13786 1896
rect 13909 1887 13967 1893
rect 13909 1884 13921 1887
rect 13780 1856 13921 1884
rect 13780 1844 13786 1856
rect 13909 1853 13921 1856
rect 13955 1884 13967 1887
rect 14844 1884 14872 2060
rect 16206 2048 16212 2060
rect 16264 2048 16270 2100
rect 16666 2088 16672 2100
rect 16627 2060 16672 2088
rect 16666 2048 16672 2060
rect 16724 2048 16730 2100
rect 17954 2020 17960 2032
rect 15028 1992 17960 2020
rect 15028 1893 15056 1992
rect 17954 1980 17960 1992
rect 18012 1980 18018 2032
rect 16117 1955 16175 1961
rect 15304 1924 15884 1952
rect 13955 1856 14872 1884
rect 15013 1887 15071 1893
rect 13955 1853 13967 1856
rect 13909 1847 13967 1853
rect 15013 1853 15025 1887
rect 15059 1884 15071 1887
rect 15102 1884 15108 1896
rect 15059 1856 15108 1884
rect 15059 1853 15071 1856
rect 15013 1847 15071 1853
rect 15102 1844 15108 1856
rect 15160 1844 15166 1896
rect 15304 1893 15332 1924
rect 15289 1887 15347 1893
rect 15289 1853 15301 1887
rect 15335 1853 15347 1887
rect 15289 1847 15347 1853
rect 15378 1844 15384 1896
rect 15436 1884 15442 1896
rect 15436 1856 15481 1884
rect 15436 1844 15442 1856
rect 15562 1844 15568 1896
rect 15620 1884 15626 1896
rect 15856 1884 15884 1924
rect 16117 1921 16129 1955
rect 16163 1952 16175 1955
rect 16298 1952 16304 1964
rect 16163 1924 16304 1952
rect 16163 1921 16175 1924
rect 16117 1915 16175 1921
rect 16298 1912 16304 1924
rect 16356 1912 16362 1964
rect 16850 1884 16856 1896
rect 15620 1856 15665 1884
rect 15856 1856 16856 1884
rect 15620 1844 15626 1856
rect 16850 1844 16856 1856
rect 16908 1844 16914 1896
rect 17681 1887 17739 1893
rect 17681 1853 17693 1887
rect 17727 1853 17739 1887
rect 17681 1847 17739 1853
rect 17957 1887 18015 1893
rect 17957 1853 17969 1887
rect 18003 1884 18015 1887
rect 18003 1856 18460 1884
rect 18003 1853 18015 1856
rect 17957 1847 18015 1853
rect 17696 1816 17724 1847
rect 11471 1788 13584 1816
rect 13648 1788 17724 1816
rect 11471 1785 11483 1788
rect 11425 1779 11483 1785
rect 2958 1708 2964 1760
rect 3016 1748 3022 1760
rect 3237 1751 3295 1757
rect 3237 1748 3249 1751
rect 3016 1720 3249 1748
rect 3016 1708 3022 1720
rect 3237 1717 3249 1720
rect 3283 1717 3295 1751
rect 3237 1711 3295 1717
rect 4062 1708 4068 1760
rect 4120 1748 4126 1760
rect 4433 1751 4491 1757
rect 4433 1748 4445 1751
rect 4120 1720 4445 1748
rect 4120 1708 4126 1720
rect 4433 1717 4445 1720
rect 4479 1717 4491 1751
rect 7558 1748 7564 1760
rect 7519 1720 7564 1748
rect 4433 1711 4491 1717
rect 7558 1708 7564 1720
rect 7616 1708 7622 1760
rect 11514 1748 11520 1760
rect 11475 1720 11520 1748
rect 11514 1708 11520 1720
rect 11572 1708 11578 1760
rect 12529 1751 12587 1757
rect 12529 1717 12541 1751
rect 12575 1748 12587 1751
rect 12802 1748 12808 1760
rect 12575 1720 12808 1748
rect 12575 1717 12587 1720
rect 12529 1711 12587 1717
rect 12802 1708 12808 1720
rect 12860 1708 12866 1760
rect 13556 1757 13584 1788
rect 18432 1760 18460 1856
rect 13541 1751 13599 1757
rect 13541 1717 13553 1751
rect 13587 1717 13599 1751
rect 16206 1748 16212 1760
rect 16167 1720 16212 1748
rect 13541 1711 13599 1717
rect 16206 1708 16212 1720
rect 16264 1708 16270 1760
rect 16298 1708 16304 1760
rect 16356 1748 16362 1760
rect 18414 1748 18420 1760
rect 16356 1720 16401 1748
rect 18375 1720 18420 1748
rect 16356 1708 16362 1720
rect 18414 1708 18420 1720
rect 18472 1708 18478 1760
rect 184 1658 18920 1680
rect 184 1606 3106 1658
rect 3158 1606 3170 1658
rect 3222 1606 3234 1658
rect 3286 1606 3298 1658
rect 3350 1606 3362 1658
rect 3414 1606 6206 1658
rect 6258 1606 6270 1658
rect 6322 1606 6334 1658
rect 6386 1606 6398 1658
rect 6450 1606 6462 1658
rect 6514 1606 9306 1658
rect 9358 1606 9370 1658
rect 9422 1606 9434 1658
rect 9486 1606 9498 1658
rect 9550 1606 9562 1658
rect 9614 1606 12406 1658
rect 12458 1606 12470 1658
rect 12522 1606 12534 1658
rect 12586 1606 12598 1658
rect 12650 1606 12662 1658
rect 12714 1606 15506 1658
rect 15558 1606 15570 1658
rect 15622 1606 15634 1658
rect 15686 1606 15698 1658
rect 15750 1606 15762 1658
rect 15814 1606 18606 1658
rect 18658 1606 18670 1658
rect 18722 1606 18734 1658
rect 18786 1606 18798 1658
rect 18850 1606 18862 1658
rect 18914 1606 18920 1658
rect 184 1584 18920 1606
rect 2225 1547 2283 1553
rect 2225 1513 2237 1547
rect 2271 1544 2283 1547
rect 3145 1547 3203 1553
rect 3145 1544 3157 1547
rect 2271 1516 3157 1544
rect 2271 1513 2283 1516
rect 2225 1507 2283 1513
rect 3145 1513 3157 1516
rect 3191 1513 3203 1547
rect 5626 1544 5632 1556
rect 3145 1507 3203 1513
rect 3804 1516 5488 1544
rect 5587 1516 5632 1544
rect 934 1436 940 1488
rect 992 1476 998 1488
rect 992 1448 2820 1476
rect 992 1436 998 1448
rect 2409 1411 2467 1417
rect 2409 1377 2421 1411
rect 2455 1408 2467 1411
rect 2682 1408 2688 1420
rect 2455 1380 2688 1408
rect 2455 1377 2467 1380
rect 2409 1371 2467 1377
rect 2682 1368 2688 1380
rect 2740 1368 2746 1420
rect 2792 1281 2820 1448
rect 2866 1436 2872 1488
rect 2924 1476 2930 1488
rect 3804 1485 3832 1516
rect 3237 1479 3295 1485
rect 3237 1476 3249 1479
rect 2924 1448 3249 1476
rect 2924 1436 2930 1448
rect 3237 1445 3249 1448
rect 3283 1476 3295 1479
rect 3789 1479 3847 1485
rect 3789 1476 3801 1479
rect 3283 1448 3801 1476
rect 3283 1445 3295 1448
rect 3237 1439 3295 1445
rect 3789 1445 3801 1448
rect 3835 1445 3847 1479
rect 3789 1439 3847 1445
rect 4801 1479 4859 1485
rect 4801 1445 4813 1479
rect 4847 1476 4859 1479
rect 5460 1476 5488 1516
rect 5626 1504 5632 1516
rect 5684 1504 5690 1556
rect 9122 1504 9128 1556
rect 9180 1504 9186 1556
rect 9582 1504 9588 1556
rect 9640 1544 9646 1556
rect 9640 1516 10272 1544
rect 9640 1504 9646 1516
rect 6546 1476 6552 1488
rect 4847 1448 5396 1476
rect 5460 1448 6552 1476
rect 4847 1445 4859 1448
rect 4801 1439 4859 1445
rect 3970 1368 3976 1420
rect 4028 1408 4034 1420
rect 4525 1411 4583 1417
rect 4525 1408 4537 1411
rect 4028 1380 4537 1408
rect 4028 1368 4034 1380
rect 4525 1377 4537 1380
rect 4571 1377 4583 1411
rect 5258 1408 5264 1420
rect 5219 1380 5264 1408
rect 4525 1371 4583 1377
rect 5258 1368 5264 1380
rect 5316 1368 5322 1420
rect 5368 1417 5396 1448
rect 6546 1436 6552 1448
rect 6604 1436 6610 1488
rect 7282 1436 7288 1488
rect 7340 1476 7346 1488
rect 7561 1479 7619 1485
rect 7561 1476 7573 1479
rect 7340 1448 7573 1476
rect 7340 1436 7346 1448
rect 7561 1445 7573 1448
rect 7607 1445 7619 1479
rect 9140 1476 9168 1504
rect 10244 1485 10272 1516
rect 11514 1504 11520 1556
rect 11572 1544 11578 1556
rect 11701 1547 11759 1553
rect 11701 1544 11713 1547
rect 11572 1516 11713 1544
rect 11572 1504 11578 1516
rect 11701 1513 11713 1516
rect 11747 1513 11759 1547
rect 13170 1544 13176 1556
rect 13131 1516 13176 1544
rect 11701 1507 11759 1513
rect 13170 1504 13176 1516
rect 13228 1504 13234 1556
rect 14001 1547 14059 1553
rect 14001 1544 14013 1547
rect 13372 1516 14013 1544
rect 10229 1479 10287 1485
rect 9140 1448 9996 1476
rect 7561 1439 7619 1445
rect 5354 1411 5412 1417
rect 5354 1377 5366 1411
rect 5400 1377 5412 1411
rect 5354 1371 5412 1377
rect 6825 1411 6883 1417
rect 6825 1377 6837 1411
rect 6871 1408 6883 1411
rect 8021 1411 8079 1417
rect 8021 1408 8033 1411
rect 6871 1380 8033 1408
rect 6871 1377 6883 1380
rect 6825 1371 6883 1377
rect 8021 1377 8033 1380
rect 8067 1408 8079 1411
rect 8110 1408 8116 1420
rect 8067 1380 8116 1408
rect 8067 1377 8079 1380
rect 8021 1371 8079 1377
rect 8110 1368 8116 1380
rect 8168 1408 8174 1420
rect 8754 1408 8760 1420
rect 8168 1380 8760 1408
rect 8168 1368 8174 1380
rect 8754 1368 8760 1380
rect 8812 1368 8818 1420
rect 8938 1368 8944 1420
rect 8996 1408 9002 1420
rect 9968 1417 9996 1448
rect 10229 1445 10241 1479
rect 10275 1445 10287 1479
rect 10229 1439 10287 1445
rect 9063 1411 9121 1417
rect 9063 1408 9075 1411
rect 8996 1380 9075 1408
rect 8996 1368 9002 1380
rect 9063 1377 9075 1380
rect 9109 1377 9121 1411
rect 9063 1371 9121 1377
rect 9217 1411 9275 1417
rect 9217 1377 9229 1411
rect 9263 1377 9275 1411
rect 9217 1371 9275 1377
rect 9953 1411 10011 1417
rect 9953 1377 9965 1411
rect 9999 1377 10011 1411
rect 9953 1371 10011 1377
rect 10965 1411 11023 1417
rect 10965 1377 10977 1411
rect 11011 1408 11023 1411
rect 11422 1408 11428 1420
rect 11011 1380 11428 1408
rect 11011 1377 11023 1380
rect 10965 1371 11023 1377
rect 3421 1343 3479 1349
rect 3421 1309 3433 1343
rect 3467 1340 3479 1343
rect 4062 1340 4068 1352
rect 3467 1312 4068 1340
rect 3467 1309 3479 1312
rect 3421 1303 3479 1309
rect 4062 1300 4068 1312
rect 4120 1300 4126 1352
rect 4614 1300 4620 1352
rect 4672 1340 4678 1352
rect 4801 1343 4859 1349
rect 4801 1340 4813 1343
rect 4672 1312 4813 1340
rect 4672 1300 4678 1312
rect 4801 1309 4813 1312
rect 4847 1340 4859 1343
rect 5442 1340 5448 1352
rect 4847 1312 5448 1340
rect 4847 1309 4859 1312
rect 4801 1303 4859 1309
rect 5442 1300 5448 1312
rect 5500 1300 5506 1352
rect 6733 1343 6791 1349
rect 6733 1309 6745 1343
rect 6779 1340 6791 1343
rect 9232 1340 9260 1371
rect 11422 1368 11428 1380
rect 11480 1368 11486 1420
rect 11790 1408 11796 1420
rect 11751 1380 11796 1408
rect 11790 1368 11796 1380
rect 11848 1368 11854 1420
rect 13372 1417 13400 1516
rect 14001 1513 14013 1516
rect 14047 1544 14059 1547
rect 14366 1544 14372 1556
rect 14047 1516 14372 1544
rect 14047 1513 14059 1516
rect 14001 1507 14059 1513
rect 14366 1504 14372 1516
rect 14424 1504 14430 1556
rect 15473 1547 15531 1553
rect 15473 1513 15485 1547
rect 15519 1544 15531 1547
rect 16298 1544 16304 1556
rect 15519 1516 16304 1544
rect 15519 1513 15531 1516
rect 15473 1507 15531 1513
rect 16298 1504 16304 1516
rect 16356 1504 16362 1556
rect 17405 1547 17463 1553
rect 17405 1513 17417 1547
rect 17451 1544 17463 1547
rect 17586 1544 17592 1556
rect 17451 1516 17592 1544
rect 17451 1513 17463 1516
rect 17405 1507 17463 1513
rect 17586 1504 17592 1516
rect 17644 1504 17650 1556
rect 18049 1547 18107 1553
rect 18049 1513 18061 1547
rect 18095 1513 18107 1547
rect 18049 1507 18107 1513
rect 15378 1436 15384 1488
rect 15436 1476 15442 1488
rect 15749 1479 15807 1485
rect 15749 1476 15761 1479
rect 15436 1448 15761 1476
rect 15436 1436 15442 1448
rect 15749 1445 15761 1448
rect 15795 1445 15807 1479
rect 18064 1476 18092 1507
rect 15749 1439 15807 1445
rect 17788 1448 18092 1476
rect 13357 1411 13415 1417
rect 13357 1377 13369 1411
rect 13403 1377 13415 1411
rect 13357 1371 13415 1377
rect 13541 1411 13599 1417
rect 13541 1377 13553 1411
rect 13587 1408 13599 1411
rect 13998 1408 14004 1420
rect 13587 1380 14004 1408
rect 13587 1377 13599 1380
rect 13541 1371 13599 1377
rect 13998 1368 14004 1380
rect 14056 1368 14062 1420
rect 15102 1408 15108 1420
rect 15063 1380 15108 1408
rect 15102 1368 15108 1380
rect 15160 1368 15166 1420
rect 15838 1408 15844 1420
rect 15799 1380 15844 1408
rect 15838 1368 15844 1380
rect 15896 1368 15902 1420
rect 17494 1368 17500 1420
rect 17552 1408 17558 1420
rect 17788 1417 17816 1448
rect 17619 1411 17677 1417
rect 17619 1408 17631 1411
rect 17552 1380 17631 1408
rect 17552 1368 17558 1380
rect 17619 1377 17631 1380
rect 17665 1377 17677 1411
rect 17619 1371 17677 1377
rect 17773 1411 17831 1417
rect 17773 1377 17785 1411
rect 17819 1377 17831 1411
rect 18049 1411 18107 1417
rect 18049 1408 18061 1411
rect 17773 1371 17831 1377
rect 17880 1380 18061 1408
rect 10873 1343 10931 1349
rect 6779 1312 8708 1340
rect 9232 1312 9996 1340
rect 6779 1309 6791 1312
rect 6733 1303 6791 1309
rect 8680 1284 8708 1312
rect 2777 1275 2835 1281
rect 2777 1241 2789 1275
rect 2823 1241 2835 1275
rect 2777 1235 2835 1241
rect 2866 1232 2872 1284
rect 2924 1272 2930 1284
rect 5166 1272 5172 1284
rect 2924 1244 5172 1272
rect 2924 1232 2930 1244
rect 4632 1213 4660 1244
rect 5166 1232 5172 1244
rect 5224 1232 5230 1284
rect 7193 1275 7251 1281
rect 7193 1241 7205 1275
rect 7239 1272 7251 1275
rect 8570 1272 8576 1284
rect 7239 1244 8576 1272
rect 7239 1241 7251 1244
rect 7193 1235 7251 1241
rect 8570 1232 8576 1244
rect 8628 1232 8634 1284
rect 8662 1232 8668 1284
rect 8720 1272 8726 1284
rect 9968 1281 9996 1312
rect 10873 1309 10885 1343
rect 10919 1340 10931 1343
rect 11808 1340 11836 1368
rect 10919 1312 11836 1340
rect 13633 1343 13691 1349
rect 10919 1309 10931 1312
rect 10873 1303 10931 1309
rect 13633 1309 13645 1343
rect 13679 1340 13691 1343
rect 13722 1340 13728 1352
rect 13679 1312 13728 1340
rect 13679 1309 13691 1312
rect 13633 1303 13691 1309
rect 13722 1300 13728 1312
rect 13780 1300 13786 1352
rect 15013 1343 15071 1349
rect 15013 1309 15025 1343
rect 15059 1340 15071 1343
rect 15856 1340 15884 1368
rect 15059 1312 15884 1340
rect 15059 1309 15071 1312
rect 15013 1303 15071 1309
rect 16850 1300 16856 1352
rect 16908 1340 16914 1352
rect 17402 1340 17408 1352
rect 16908 1312 17408 1340
rect 16908 1300 16914 1312
rect 17402 1300 17408 1312
rect 17460 1340 17466 1352
rect 17880 1340 17908 1380
rect 18049 1377 18061 1380
rect 18095 1377 18107 1411
rect 18049 1371 18107 1377
rect 18325 1411 18383 1417
rect 18325 1377 18337 1411
rect 18371 1377 18383 1411
rect 18325 1371 18383 1377
rect 17460 1312 17908 1340
rect 17460 1300 17466 1312
rect 17954 1300 17960 1352
rect 18012 1340 18018 1352
rect 18340 1340 18368 1371
rect 18012 1312 18368 1340
rect 18012 1300 18018 1312
rect 9953 1275 10011 1281
rect 8720 1244 9904 1272
rect 8720 1232 8726 1244
rect 4617 1207 4675 1213
rect 4617 1173 4629 1207
rect 4663 1173 4675 1207
rect 9030 1204 9036 1216
rect 8991 1176 9036 1204
rect 4617 1167 4675 1173
rect 9030 1164 9036 1176
rect 9088 1164 9094 1216
rect 9876 1204 9904 1244
rect 9953 1241 9965 1275
rect 9999 1241 10011 1275
rect 9953 1235 10011 1241
rect 10045 1275 10103 1281
rect 10045 1241 10057 1275
rect 10091 1241 10103 1275
rect 10045 1235 10103 1241
rect 11333 1275 11391 1281
rect 11333 1241 11345 1275
rect 11379 1272 11391 1275
rect 12802 1272 12808 1284
rect 11379 1244 12808 1272
rect 11379 1241 11391 1244
rect 11333 1235 11391 1241
rect 10060 1204 10088 1235
rect 12802 1232 12808 1244
rect 12860 1232 12866 1284
rect 17586 1232 17592 1284
rect 17644 1272 17650 1284
rect 18141 1275 18199 1281
rect 18141 1272 18153 1275
rect 17644 1244 18153 1272
rect 17644 1232 17650 1244
rect 18141 1241 18153 1244
rect 18187 1241 18199 1275
rect 18141 1235 18199 1241
rect 9876 1176 10088 1204
rect 184 1114 18860 1136
rect 184 1062 1556 1114
rect 1608 1062 1620 1114
rect 1672 1062 1684 1114
rect 1736 1062 1748 1114
rect 1800 1062 1812 1114
rect 1864 1062 4656 1114
rect 4708 1062 4720 1114
rect 4772 1062 4784 1114
rect 4836 1062 4848 1114
rect 4900 1062 4912 1114
rect 4964 1062 7756 1114
rect 7808 1062 7820 1114
rect 7872 1062 7884 1114
rect 7936 1062 7948 1114
rect 8000 1062 8012 1114
rect 8064 1062 10856 1114
rect 10908 1062 10920 1114
rect 10972 1062 10984 1114
rect 11036 1062 11048 1114
rect 11100 1062 11112 1114
rect 11164 1062 13956 1114
rect 14008 1062 14020 1114
rect 14072 1062 14084 1114
rect 14136 1062 14148 1114
rect 14200 1062 14212 1114
rect 14264 1062 17056 1114
rect 17108 1062 17120 1114
rect 17172 1062 17184 1114
rect 17236 1062 17248 1114
rect 17300 1062 17312 1114
rect 17364 1062 18860 1114
rect 184 1040 18860 1062
rect 2958 960 2964 1012
rect 3016 1000 3022 1012
rect 3237 1003 3295 1009
rect 3237 1000 3249 1003
rect 3016 972 3249 1000
rect 3016 960 3022 972
rect 3237 969 3249 972
rect 3283 969 3295 1003
rect 5258 1000 5264 1012
rect 5219 972 5264 1000
rect 3237 963 3295 969
rect 5258 960 5264 972
rect 5316 960 5322 1012
rect 8938 1000 8944 1012
rect 8899 972 8944 1000
rect 8938 960 8944 972
rect 8996 960 9002 1012
rect 17494 1000 17500 1012
rect 17455 972 17500 1000
rect 17494 960 17500 972
rect 17552 960 17558 1012
rect 17586 960 17592 1012
rect 17644 1000 17650 1012
rect 17644 972 17689 1000
rect 17644 960 17650 972
rect 5166 892 5172 944
rect 5224 932 5230 944
rect 5353 935 5411 941
rect 5353 932 5365 935
rect 5224 904 5365 932
rect 5224 892 5230 904
rect 5353 901 5365 904
rect 5399 901 5411 935
rect 5353 895 5411 901
rect 8662 892 8668 944
rect 8720 932 8726 944
rect 9033 935 9091 941
rect 9033 932 9045 935
rect 8720 904 9045 932
rect 8720 892 8726 904
rect 9033 901 9045 904
rect 9079 901 9091 935
rect 9033 895 9091 901
rect 9122 892 9128 944
rect 9180 892 9186 944
rect 15838 892 15844 944
rect 15896 932 15902 944
rect 17604 932 17632 960
rect 15896 904 17632 932
rect 15896 892 15902 904
rect 2774 824 2780 876
rect 2832 864 2838 876
rect 2869 867 2927 873
rect 2869 864 2881 867
rect 2832 836 2881 864
rect 2832 824 2838 836
rect 2869 833 2881 836
rect 2915 833 2927 867
rect 2869 827 2927 833
rect 8849 867 8907 873
rect 8849 833 8861 867
rect 8895 864 8907 867
rect 9140 864 9168 892
rect 17402 864 17408 876
rect 8895 836 9168 864
rect 17363 836 17408 864
rect 8895 833 8907 836
rect 8849 827 8907 833
rect 17402 824 17408 836
rect 17460 824 17466 876
rect 2961 799 3019 805
rect 2961 765 2973 799
rect 3007 796 3019 799
rect 3970 796 3976 808
rect 3007 768 3976 796
rect 3007 765 3019 768
rect 2961 759 3019 765
rect 3970 756 3976 768
rect 4028 796 4034 808
rect 5169 799 5227 805
rect 5169 796 5181 799
rect 4028 768 5181 796
rect 4028 756 4034 768
rect 5169 765 5181 768
rect 5215 765 5227 799
rect 5442 796 5448 808
rect 5403 768 5448 796
rect 5169 759 5227 765
rect 5442 756 5448 768
rect 5500 756 5506 808
rect 8754 756 8760 808
rect 8812 796 8818 808
rect 9125 799 9183 805
rect 9125 796 9137 799
rect 8812 768 9137 796
rect 8812 756 8818 768
rect 9125 765 9137 768
rect 9171 796 9183 799
rect 9582 796 9588 808
rect 9171 768 9588 796
rect 9171 765 9183 768
rect 9125 759 9183 765
rect 9582 756 9588 768
rect 9640 756 9646 808
rect 17681 799 17739 805
rect 17681 765 17693 799
rect 17727 796 17739 799
rect 17954 796 17960 808
rect 17727 768 17960 796
rect 17727 765 17739 768
rect 17681 759 17739 765
rect 17954 756 17960 768
rect 18012 756 18018 808
rect 184 570 18920 592
rect 184 518 3106 570
rect 3158 518 3170 570
rect 3222 518 3234 570
rect 3286 518 3298 570
rect 3350 518 3362 570
rect 3414 518 6206 570
rect 6258 518 6270 570
rect 6322 518 6334 570
rect 6386 518 6398 570
rect 6450 518 6462 570
rect 6514 518 9306 570
rect 9358 518 9370 570
rect 9422 518 9434 570
rect 9486 518 9498 570
rect 9550 518 9562 570
rect 9614 518 12406 570
rect 12458 518 12470 570
rect 12522 518 12534 570
rect 12586 518 12598 570
rect 12650 518 12662 570
rect 12714 518 15506 570
rect 15558 518 15570 570
rect 15622 518 15634 570
rect 15686 518 15698 570
rect 15750 518 15762 570
rect 15814 518 18606 570
rect 18658 518 18670 570
rect 18722 518 18734 570
rect 18786 518 18798 570
rect 18850 518 18862 570
rect 18914 518 18920 570
rect 184 496 18920 518
<< via1 >>
rect 1556 18470 1608 18522
rect 1620 18470 1672 18522
rect 1684 18470 1736 18522
rect 1748 18470 1800 18522
rect 1812 18470 1864 18522
rect 4656 18470 4708 18522
rect 4720 18470 4772 18522
rect 4784 18470 4836 18522
rect 4848 18470 4900 18522
rect 4912 18470 4964 18522
rect 7756 18470 7808 18522
rect 7820 18470 7872 18522
rect 7884 18470 7936 18522
rect 7948 18470 8000 18522
rect 8012 18470 8064 18522
rect 10856 18470 10908 18522
rect 10920 18470 10972 18522
rect 10984 18470 11036 18522
rect 11048 18470 11100 18522
rect 11112 18470 11164 18522
rect 13956 18470 14008 18522
rect 14020 18470 14072 18522
rect 14084 18470 14136 18522
rect 14148 18470 14200 18522
rect 14212 18470 14264 18522
rect 17056 18470 17108 18522
rect 17120 18470 17172 18522
rect 17184 18470 17236 18522
rect 17248 18470 17300 18522
rect 17312 18470 17364 18522
rect 1400 18368 1452 18420
rect 18420 18411 18472 18420
rect 18420 18377 18429 18411
rect 18429 18377 18463 18411
rect 18463 18377 18472 18411
rect 18420 18368 18472 18377
rect 1400 18164 1452 18216
rect 1952 18164 2004 18216
rect 4436 18232 4488 18284
rect 5724 18232 5776 18284
rect 1216 18028 1268 18080
rect 5448 18096 5500 18148
rect 6552 18096 6604 18148
rect 7104 18164 7156 18216
rect 7288 18164 7340 18216
rect 11152 18300 11204 18352
rect 9680 18232 9732 18284
rect 16028 18232 16080 18284
rect 8392 18139 8444 18148
rect 2964 18071 3016 18080
rect 2964 18037 2973 18071
rect 2973 18037 3007 18071
rect 3007 18037 3016 18071
rect 2964 18028 3016 18037
rect 4068 18071 4120 18080
rect 4068 18037 4077 18071
rect 4077 18037 4111 18071
rect 4111 18037 4120 18071
rect 4068 18028 4120 18037
rect 4344 18028 4396 18080
rect 4528 18071 4580 18080
rect 4528 18037 4537 18071
rect 4537 18037 4571 18071
rect 4571 18037 4580 18071
rect 5540 18071 5592 18080
rect 4528 18028 4580 18037
rect 5540 18037 5549 18071
rect 5549 18037 5583 18071
rect 5583 18037 5592 18071
rect 5540 18028 5592 18037
rect 7840 18028 7892 18080
rect 8392 18105 8401 18139
rect 8401 18105 8435 18139
rect 8435 18105 8444 18139
rect 8392 18096 8444 18105
rect 9956 18096 10008 18148
rect 11152 18207 11204 18216
rect 11152 18173 11161 18207
rect 11161 18173 11195 18207
rect 11195 18173 11204 18207
rect 11152 18164 11204 18173
rect 12440 18207 12492 18216
rect 12440 18173 12449 18207
rect 12449 18173 12483 18207
rect 12483 18173 12492 18207
rect 12440 18164 12492 18173
rect 11336 18096 11388 18148
rect 11428 18139 11480 18148
rect 11428 18105 11437 18139
rect 11437 18105 11471 18139
rect 11471 18105 11480 18139
rect 11428 18096 11480 18105
rect 8484 18028 8536 18080
rect 10140 18028 10192 18080
rect 11244 18028 11296 18080
rect 13452 18028 13504 18080
rect 18420 18164 18472 18216
rect 3106 17926 3158 17978
rect 3170 17926 3222 17978
rect 3234 17926 3286 17978
rect 3298 17926 3350 17978
rect 3362 17926 3414 17978
rect 6206 17926 6258 17978
rect 6270 17926 6322 17978
rect 6334 17926 6386 17978
rect 6398 17926 6450 17978
rect 6462 17926 6514 17978
rect 9306 17926 9358 17978
rect 9370 17926 9422 17978
rect 9434 17926 9486 17978
rect 9498 17926 9550 17978
rect 9562 17926 9614 17978
rect 12406 17926 12458 17978
rect 12470 17926 12522 17978
rect 12534 17926 12586 17978
rect 12598 17926 12650 17978
rect 12662 17926 12714 17978
rect 15506 17926 15558 17978
rect 15570 17926 15622 17978
rect 15634 17926 15686 17978
rect 15698 17926 15750 17978
rect 15762 17926 15814 17978
rect 18606 17926 18658 17978
rect 18670 17926 18722 17978
rect 18734 17926 18786 17978
rect 18798 17926 18850 17978
rect 18862 17926 18914 17978
rect 4528 17824 4580 17876
rect 12256 17824 12308 17876
rect 1216 17756 1268 17808
rect 2504 17756 2556 17808
rect 4252 17756 4304 17808
rect 7840 17799 7892 17808
rect 7840 17765 7849 17799
rect 7849 17765 7883 17799
rect 7883 17765 7892 17799
rect 7840 17756 7892 17765
rect 13084 17756 13136 17808
rect 9956 17731 10008 17740
rect 572 17620 624 17672
rect 4252 17620 4304 17672
rect 9956 17697 9965 17731
rect 9965 17697 9999 17731
rect 9999 17697 10008 17731
rect 9956 17688 10008 17697
rect 12256 17688 12308 17740
rect 17500 17731 17552 17740
rect 17500 17697 17509 17731
rect 17509 17697 17543 17731
rect 17543 17697 17552 17731
rect 17500 17688 17552 17697
rect 10324 17663 10376 17672
rect 10324 17629 10333 17663
rect 10333 17629 10367 17663
rect 10367 17629 10376 17663
rect 10324 17620 10376 17629
rect 13820 17620 13872 17672
rect 14740 17663 14792 17672
rect 14740 17629 14749 17663
rect 14749 17629 14783 17663
rect 14783 17629 14792 17663
rect 14740 17620 14792 17629
rect 15108 17663 15160 17672
rect 15108 17629 15117 17663
rect 15117 17629 15151 17663
rect 15151 17629 15160 17663
rect 15108 17620 15160 17629
rect 16948 17620 17000 17672
rect 17684 17620 17736 17672
rect 17868 17620 17920 17672
rect 2412 17527 2464 17536
rect 2412 17493 2421 17527
rect 2421 17493 2455 17527
rect 2455 17493 2464 17527
rect 2412 17484 2464 17493
rect 7012 17484 7064 17536
rect 14280 17552 14332 17604
rect 11980 17484 12032 17536
rect 16856 17484 16908 17536
rect 1556 17382 1608 17434
rect 1620 17382 1672 17434
rect 1684 17382 1736 17434
rect 1748 17382 1800 17434
rect 1812 17382 1864 17434
rect 4656 17382 4708 17434
rect 4720 17382 4772 17434
rect 4784 17382 4836 17434
rect 4848 17382 4900 17434
rect 4912 17382 4964 17434
rect 7756 17382 7808 17434
rect 7820 17382 7872 17434
rect 7884 17382 7936 17434
rect 7948 17382 8000 17434
rect 8012 17382 8064 17434
rect 10856 17382 10908 17434
rect 10920 17382 10972 17434
rect 10984 17382 11036 17434
rect 11048 17382 11100 17434
rect 11112 17382 11164 17434
rect 13956 17382 14008 17434
rect 14020 17382 14072 17434
rect 14084 17382 14136 17434
rect 14148 17382 14200 17434
rect 14212 17382 14264 17434
rect 17056 17382 17108 17434
rect 17120 17382 17172 17434
rect 17184 17382 17236 17434
rect 17248 17382 17300 17434
rect 17312 17382 17364 17434
rect 1952 17280 2004 17332
rect 4160 17280 4212 17332
rect 5540 17280 5592 17332
rect 10048 17280 10100 17332
rect 10324 17212 10376 17264
rect 2504 17187 2556 17196
rect 2504 17153 2513 17187
rect 2513 17153 2547 17187
rect 2547 17153 2556 17187
rect 2504 17144 2556 17153
rect 4344 17187 4396 17196
rect 4344 17153 4353 17187
rect 4353 17153 4387 17187
rect 4387 17153 4396 17187
rect 4344 17144 4396 17153
rect 6552 17187 6604 17196
rect 6552 17153 6561 17187
rect 6561 17153 6595 17187
rect 6595 17153 6604 17187
rect 6552 17144 6604 17153
rect 7288 17144 7340 17196
rect 8392 17144 8444 17196
rect 1584 17119 1636 17128
rect 1584 17085 1593 17119
rect 1593 17085 1627 17119
rect 1627 17085 1636 17119
rect 1584 17076 1636 17085
rect 1768 17119 1820 17128
rect 1768 17085 1777 17119
rect 1777 17085 1811 17119
rect 1811 17085 1820 17119
rect 1768 17076 1820 17085
rect 1860 17076 1912 17128
rect 2228 17076 2280 17128
rect 2320 17119 2372 17128
rect 2320 17085 2329 17119
rect 2329 17085 2363 17119
rect 2363 17085 2372 17119
rect 2320 17076 2372 17085
rect 2964 17076 3016 17128
rect 3516 17076 3568 17128
rect 2504 17008 2556 17060
rect 4436 17008 4488 17060
rect 6828 16940 6880 16992
rect 11244 17076 11296 17128
rect 13084 17008 13136 17060
rect 14740 17144 14792 17196
rect 16856 17144 16908 17196
rect 17684 17280 17736 17332
rect 16580 17008 16632 17060
rect 15936 16940 15988 16992
rect 3106 16838 3158 16890
rect 3170 16838 3222 16890
rect 3234 16838 3286 16890
rect 3298 16838 3350 16890
rect 3362 16838 3414 16890
rect 6206 16838 6258 16890
rect 6270 16838 6322 16890
rect 6334 16838 6386 16890
rect 6398 16838 6450 16890
rect 6462 16838 6514 16890
rect 9306 16838 9358 16890
rect 9370 16838 9422 16890
rect 9434 16838 9486 16890
rect 9498 16838 9550 16890
rect 9562 16838 9614 16890
rect 12406 16838 12458 16890
rect 12470 16838 12522 16890
rect 12534 16838 12586 16890
rect 12598 16838 12650 16890
rect 12662 16838 12714 16890
rect 15506 16838 15558 16890
rect 15570 16838 15622 16890
rect 15634 16838 15686 16890
rect 15698 16838 15750 16890
rect 15762 16838 15814 16890
rect 18606 16838 18658 16890
rect 18670 16838 18722 16890
rect 18734 16838 18786 16890
rect 18798 16838 18850 16890
rect 18862 16838 18914 16890
rect 1676 16779 1728 16788
rect 1676 16745 1685 16779
rect 1685 16745 1719 16779
rect 1719 16745 1728 16779
rect 1676 16736 1728 16745
rect 1584 16711 1636 16720
rect 1584 16677 1593 16711
rect 1593 16677 1627 16711
rect 1627 16677 1636 16711
rect 2412 16736 2464 16788
rect 1584 16668 1636 16677
rect 1860 16643 1912 16652
rect 1860 16609 1869 16643
rect 1869 16609 1903 16643
rect 1903 16609 1912 16643
rect 4344 16736 4396 16788
rect 12164 16736 12216 16788
rect 16028 16779 16080 16788
rect 4068 16668 4120 16720
rect 7012 16711 7064 16720
rect 7012 16677 7021 16711
rect 7021 16677 7055 16711
rect 7055 16677 7064 16711
rect 7012 16668 7064 16677
rect 10232 16668 10284 16720
rect 12532 16668 12584 16720
rect 13084 16668 13136 16720
rect 1860 16600 1912 16609
rect 1768 16575 1820 16584
rect 1768 16541 1777 16575
rect 1777 16541 1811 16575
rect 1811 16541 1820 16575
rect 1768 16532 1820 16541
rect 2228 16532 2280 16584
rect 572 16464 624 16516
rect 3516 16600 3568 16652
rect 16028 16745 16037 16779
rect 16037 16745 16071 16779
rect 16071 16745 16080 16779
rect 16028 16736 16080 16745
rect 17500 16736 17552 16788
rect 14280 16668 14332 16720
rect 17500 16600 17552 16652
rect 18420 16643 18472 16652
rect 18420 16609 18429 16643
rect 18429 16609 18463 16643
rect 18463 16609 18472 16643
rect 18420 16600 18472 16609
rect 7656 16532 7708 16584
rect 10140 16532 10192 16584
rect 1768 16396 1820 16448
rect 2044 16396 2096 16448
rect 2780 16396 2832 16448
rect 3424 16396 3476 16448
rect 7472 16396 7524 16448
rect 12072 16396 12124 16448
rect 12716 16396 12768 16448
rect 17684 16575 17736 16584
rect 17684 16541 17693 16575
rect 17693 16541 17727 16575
rect 17727 16541 17736 16575
rect 17684 16532 17736 16541
rect 17776 16575 17828 16584
rect 17776 16541 17785 16575
rect 17785 16541 17819 16575
rect 17819 16541 17828 16575
rect 17776 16532 17828 16541
rect 18052 16464 18104 16516
rect 1556 16294 1608 16346
rect 1620 16294 1672 16346
rect 1684 16294 1736 16346
rect 1748 16294 1800 16346
rect 1812 16294 1864 16346
rect 4656 16294 4708 16346
rect 4720 16294 4772 16346
rect 4784 16294 4836 16346
rect 4848 16294 4900 16346
rect 4912 16294 4964 16346
rect 7756 16294 7808 16346
rect 7820 16294 7872 16346
rect 7884 16294 7936 16346
rect 7948 16294 8000 16346
rect 8012 16294 8064 16346
rect 10856 16294 10908 16346
rect 10920 16294 10972 16346
rect 10984 16294 11036 16346
rect 11048 16294 11100 16346
rect 11112 16294 11164 16346
rect 13956 16294 14008 16346
rect 14020 16294 14072 16346
rect 14084 16294 14136 16346
rect 14148 16294 14200 16346
rect 14212 16294 14264 16346
rect 17056 16294 17108 16346
rect 17120 16294 17172 16346
rect 17184 16294 17236 16346
rect 17248 16294 17300 16346
rect 17312 16294 17364 16346
rect 5448 16192 5500 16244
rect 7104 16192 7156 16244
rect 11336 16192 11388 16244
rect 16120 16192 16172 16244
rect 17776 16192 17828 16244
rect 18420 16235 18472 16244
rect 18420 16201 18429 16235
rect 18429 16201 18463 16235
rect 18463 16201 18472 16235
rect 18420 16192 18472 16201
rect 17684 16167 17736 16176
rect 17684 16133 17693 16167
rect 17693 16133 17727 16167
rect 17727 16133 17736 16167
rect 17684 16124 17736 16133
rect 1952 16056 2004 16108
rect 2228 16099 2280 16108
rect 2228 16065 2237 16099
rect 2237 16065 2271 16099
rect 2271 16065 2280 16099
rect 2228 16056 2280 16065
rect 2780 16099 2832 16108
rect 2780 16065 2789 16099
rect 2789 16065 2823 16099
rect 2823 16065 2832 16099
rect 2780 16056 2832 16065
rect 12072 16056 12124 16108
rect 16028 16056 16080 16108
rect 16948 16056 17000 16108
rect 4252 16031 4304 16040
rect 4252 15997 4261 16031
rect 4261 15997 4295 16031
rect 4295 15997 4304 16031
rect 4252 15988 4304 15997
rect 10140 15988 10192 16040
rect 16120 16031 16172 16040
rect 16120 15997 16129 16031
rect 16129 15997 16163 16031
rect 16163 15997 16172 16031
rect 16120 15988 16172 15997
rect 2964 15920 3016 15972
rect 8760 15963 8812 15972
rect 848 15852 900 15904
rect 3700 15852 3752 15904
rect 8760 15929 8769 15963
rect 8769 15929 8803 15963
rect 8803 15929 8812 15963
rect 8760 15920 8812 15929
rect 12532 15920 12584 15972
rect 13084 15920 13136 15972
rect 15200 15920 15252 15972
rect 16304 15920 16356 15972
rect 17592 15988 17644 16040
rect 17868 15920 17920 15972
rect 15292 15895 15344 15904
rect 15292 15861 15301 15895
rect 15301 15861 15335 15895
rect 15335 15861 15344 15895
rect 15292 15852 15344 15861
rect 15936 15895 15988 15904
rect 15936 15861 15945 15895
rect 15945 15861 15979 15895
rect 15979 15861 15988 15895
rect 15936 15852 15988 15861
rect 3106 15750 3158 15802
rect 3170 15750 3222 15802
rect 3234 15750 3286 15802
rect 3298 15750 3350 15802
rect 3362 15750 3414 15802
rect 6206 15750 6258 15802
rect 6270 15750 6322 15802
rect 6334 15750 6386 15802
rect 6398 15750 6450 15802
rect 6462 15750 6514 15802
rect 9306 15750 9358 15802
rect 9370 15750 9422 15802
rect 9434 15750 9486 15802
rect 9498 15750 9550 15802
rect 9562 15750 9614 15802
rect 12406 15750 12458 15802
rect 12470 15750 12522 15802
rect 12534 15750 12586 15802
rect 12598 15750 12650 15802
rect 12662 15750 12714 15802
rect 15506 15750 15558 15802
rect 15570 15750 15622 15802
rect 15634 15750 15686 15802
rect 15698 15750 15750 15802
rect 15762 15750 15814 15802
rect 18606 15750 18658 15802
rect 18670 15750 18722 15802
rect 18734 15750 18786 15802
rect 18798 15750 18850 15802
rect 18862 15750 18914 15802
rect 848 15623 900 15632
rect 848 15589 857 15623
rect 857 15589 891 15623
rect 891 15589 900 15623
rect 848 15580 900 15589
rect 2136 15580 2188 15632
rect 2504 15580 2556 15632
rect 4160 15580 4212 15632
rect 5816 15580 5868 15632
rect 7564 15648 7616 15700
rect 9680 15648 9732 15700
rect 12808 15648 12860 15700
rect 12900 15648 12952 15700
rect 14280 15648 14332 15700
rect 15108 15648 15160 15700
rect 10140 15580 10192 15632
rect 11980 15623 12032 15632
rect 11980 15589 11989 15623
rect 11989 15589 12023 15623
rect 12023 15589 12032 15623
rect 11980 15580 12032 15589
rect 13084 15580 13136 15632
rect 16304 15648 16356 15700
rect 16580 15691 16632 15700
rect 16580 15657 16589 15691
rect 16589 15657 16623 15691
rect 16623 15657 16632 15691
rect 16580 15648 16632 15657
rect 17776 15648 17828 15700
rect 572 15555 624 15564
rect 572 15521 581 15555
rect 581 15521 615 15555
rect 615 15521 624 15555
rect 572 15512 624 15521
rect 1952 15376 2004 15428
rect 6828 15512 6880 15564
rect 5448 15487 5500 15496
rect 5448 15453 5457 15487
rect 5457 15453 5491 15487
rect 5491 15453 5500 15487
rect 5448 15444 5500 15453
rect 5724 15487 5776 15496
rect 5724 15453 5733 15487
rect 5733 15453 5767 15487
rect 5767 15453 5776 15487
rect 5724 15444 5776 15453
rect 7288 15444 7340 15496
rect 7656 15444 7708 15496
rect 11336 15444 11388 15496
rect 12164 15444 12216 15496
rect 15936 15580 15988 15632
rect 15844 15512 15896 15564
rect 16212 15555 16264 15564
rect 16212 15521 16221 15555
rect 16221 15521 16255 15555
rect 16255 15521 16264 15555
rect 16212 15512 16264 15521
rect 16488 15555 16540 15564
rect 16488 15521 16497 15555
rect 16497 15521 16531 15555
rect 16531 15521 16540 15555
rect 16488 15512 16540 15521
rect 16948 15512 17000 15564
rect 17408 15512 17460 15564
rect 15016 15444 15068 15496
rect 15936 15487 15988 15496
rect 8668 15308 8720 15360
rect 10140 15308 10192 15360
rect 15108 15308 15160 15360
rect 15936 15453 15945 15487
rect 15945 15453 15979 15487
rect 15979 15453 15988 15487
rect 15936 15444 15988 15453
rect 16948 15308 17000 15360
rect 17500 15308 17552 15360
rect 1556 15206 1608 15258
rect 1620 15206 1672 15258
rect 1684 15206 1736 15258
rect 1748 15206 1800 15258
rect 1812 15206 1864 15258
rect 4656 15206 4708 15258
rect 4720 15206 4772 15258
rect 4784 15206 4836 15258
rect 4848 15206 4900 15258
rect 4912 15206 4964 15258
rect 7756 15206 7808 15258
rect 7820 15206 7872 15258
rect 7884 15206 7936 15258
rect 7948 15206 8000 15258
rect 8012 15206 8064 15258
rect 10856 15206 10908 15258
rect 10920 15206 10972 15258
rect 10984 15206 11036 15258
rect 11048 15206 11100 15258
rect 11112 15206 11164 15258
rect 13956 15206 14008 15258
rect 14020 15206 14072 15258
rect 14084 15206 14136 15258
rect 14148 15206 14200 15258
rect 14212 15206 14264 15258
rect 17056 15206 17108 15258
rect 17120 15206 17172 15258
rect 17184 15206 17236 15258
rect 17248 15206 17300 15258
rect 17312 15206 17364 15258
rect 2228 15011 2280 15020
rect 2228 14977 2237 15011
rect 2237 14977 2271 15011
rect 2271 14977 2280 15011
rect 5080 15104 5132 15156
rect 8760 15104 8812 15156
rect 15844 15104 15896 15156
rect 3792 15036 3844 15088
rect 2228 14968 2280 14977
rect 2044 14943 2096 14952
rect 2044 14909 2053 14943
rect 2053 14909 2087 14943
rect 2087 14909 2096 14943
rect 2044 14900 2096 14909
rect 2412 14900 2464 14952
rect 3516 14900 3568 14952
rect 4436 14900 4488 14952
rect 7012 14968 7064 15020
rect 7564 14968 7616 15020
rect 14280 15011 14332 15020
rect 14280 14977 14289 15011
rect 14289 14977 14323 15011
rect 14323 14977 14332 15011
rect 14280 14968 14332 14977
rect 16120 14968 16172 15020
rect 4620 14943 4672 14952
rect 4620 14909 4629 14943
rect 4629 14909 4663 14943
rect 4663 14909 4672 14943
rect 5080 14943 5132 14952
rect 4620 14900 4672 14909
rect 5080 14909 5089 14943
rect 5089 14909 5123 14943
rect 5123 14909 5132 14943
rect 5080 14900 5132 14909
rect 4160 14875 4212 14884
rect 4160 14841 4169 14875
rect 4169 14841 4203 14875
rect 4203 14841 4212 14875
rect 4160 14832 4212 14841
rect 7472 14900 7524 14952
rect 11244 14900 11296 14952
rect 11520 14943 11572 14952
rect 11520 14909 11529 14943
rect 11529 14909 11563 14943
rect 11563 14909 11572 14943
rect 11520 14900 11572 14909
rect 13452 14900 13504 14952
rect 17592 14943 17644 14952
rect 9036 14875 9088 14884
rect 9036 14841 9045 14875
rect 9045 14841 9079 14875
rect 9079 14841 9088 14875
rect 9036 14832 9088 14841
rect 940 14764 992 14816
rect 1952 14807 2004 14816
rect 1952 14773 1961 14807
rect 1961 14773 1995 14807
rect 1995 14773 2004 14807
rect 1952 14764 2004 14773
rect 2504 14764 2556 14816
rect 5724 14807 5776 14816
rect 5724 14773 5733 14807
rect 5733 14773 5767 14807
rect 5767 14773 5776 14807
rect 5724 14764 5776 14773
rect 5816 14764 5868 14816
rect 7840 14807 7892 14816
rect 7840 14773 7849 14807
rect 7849 14773 7883 14807
rect 7883 14773 7892 14807
rect 7840 14764 7892 14773
rect 10324 14807 10376 14816
rect 10324 14773 10333 14807
rect 10333 14773 10367 14807
rect 10367 14773 10376 14807
rect 10324 14764 10376 14773
rect 11152 14764 11204 14816
rect 11888 14832 11940 14884
rect 17592 14909 17601 14943
rect 17601 14909 17635 14943
rect 17635 14909 17644 14943
rect 17592 14900 17644 14909
rect 17960 14832 18012 14884
rect 12808 14764 12860 14816
rect 15936 14764 15988 14816
rect 16120 14764 16172 14816
rect 16396 14807 16448 14816
rect 16396 14773 16405 14807
rect 16405 14773 16439 14807
rect 16439 14773 16448 14807
rect 16396 14764 16448 14773
rect 17132 14764 17184 14816
rect 17408 14764 17460 14816
rect 3106 14662 3158 14714
rect 3170 14662 3222 14714
rect 3234 14662 3286 14714
rect 3298 14662 3350 14714
rect 3362 14662 3414 14714
rect 6206 14662 6258 14714
rect 6270 14662 6322 14714
rect 6334 14662 6386 14714
rect 6398 14662 6450 14714
rect 6462 14662 6514 14714
rect 9306 14662 9358 14714
rect 9370 14662 9422 14714
rect 9434 14662 9486 14714
rect 9498 14662 9550 14714
rect 9562 14662 9614 14714
rect 12406 14662 12458 14714
rect 12470 14662 12522 14714
rect 12534 14662 12586 14714
rect 12598 14662 12650 14714
rect 12662 14662 12714 14714
rect 15506 14662 15558 14714
rect 15570 14662 15622 14714
rect 15634 14662 15686 14714
rect 15698 14662 15750 14714
rect 15762 14662 15814 14714
rect 18606 14662 18658 14714
rect 18670 14662 18722 14714
rect 18734 14662 18786 14714
rect 18798 14662 18850 14714
rect 18862 14662 18914 14714
rect 2964 14560 3016 14612
rect 3700 14603 3752 14612
rect 3700 14569 3709 14603
rect 3709 14569 3743 14603
rect 3743 14569 3752 14603
rect 3700 14560 3752 14569
rect 2136 14492 2188 14544
rect 2412 14535 2464 14544
rect 2412 14501 2421 14535
rect 2421 14501 2455 14535
rect 2455 14501 2464 14535
rect 2412 14492 2464 14501
rect 6736 14492 6788 14544
rect 8484 14492 8536 14544
rect 572 14467 624 14476
rect 572 14433 581 14467
rect 581 14433 615 14467
rect 615 14433 624 14467
rect 572 14424 624 14433
rect 940 14467 992 14476
rect 940 14433 949 14467
rect 949 14433 983 14467
rect 983 14433 992 14467
rect 940 14424 992 14433
rect 3700 14424 3752 14476
rect 4528 14424 4580 14476
rect 5448 14424 5500 14476
rect 5724 14467 5776 14476
rect 5724 14433 5733 14467
rect 5733 14433 5767 14467
rect 5767 14433 5776 14467
rect 5724 14424 5776 14433
rect 7840 14424 7892 14476
rect 8208 14424 8260 14476
rect 11428 14560 11480 14612
rect 11888 14560 11940 14612
rect 11336 14535 11388 14544
rect 11336 14501 11345 14535
rect 11345 14501 11379 14535
rect 11379 14501 11388 14535
rect 11336 14492 11388 14501
rect 16396 14560 16448 14612
rect 13084 14492 13136 14544
rect 16488 14492 16540 14544
rect 11244 14424 11296 14476
rect 12164 14424 12216 14476
rect 12808 14424 12860 14476
rect 15016 14467 15068 14476
rect 15016 14433 15025 14467
rect 15025 14433 15059 14467
rect 15059 14433 15068 14467
rect 15016 14424 15068 14433
rect 15752 14424 15804 14476
rect 3792 14399 3844 14408
rect 3792 14365 3801 14399
rect 3801 14365 3835 14399
rect 3835 14365 3844 14399
rect 3792 14356 3844 14365
rect 8116 14399 8168 14408
rect 8116 14365 8125 14399
rect 8125 14365 8159 14399
rect 8159 14365 8168 14399
rect 8116 14356 8168 14365
rect 11152 14356 11204 14408
rect 11336 14356 11388 14408
rect 15200 14356 15252 14408
rect 15568 14288 15620 14340
rect 15936 14467 15988 14476
rect 15936 14433 15945 14467
rect 15945 14433 15979 14467
rect 15979 14433 15988 14467
rect 15936 14424 15988 14433
rect 16028 14399 16080 14408
rect 16028 14365 16037 14399
rect 16037 14365 16071 14399
rect 16071 14365 16080 14399
rect 16028 14356 16080 14365
rect 17868 14467 17920 14476
rect 17868 14433 17877 14467
rect 17877 14433 17911 14467
rect 17911 14433 17920 14467
rect 17868 14424 17920 14433
rect 17960 14424 18012 14476
rect 16856 14356 16908 14408
rect 17408 14356 17460 14408
rect 17132 14288 17184 14340
rect 7012 14220 7064 14272
rect 7380 14220 7432 14272
rect 7472 14220 7524 14272
rect 11796 14220 11848 14272
rect 12900 14220 12952 14272
rect 15016 14220 15068 14272
rect 16212 14220 16264 14272
rect 16856 14220 16908 14272
rect 17592 14220 17644 14272
rect 18236 14263 18288 14272
rect 18236 14229 18245 14263
rect 18245 14229 18279 14263
rect 18279 14229 18288 14263
rect 18236 14220 18288 14229
rect 1556 14118 1608 14170
rect 1620 14118 1672 14170
rect 1684 14118 1736 14170
rect 1748 14118 1800 14170
rect 1812 14118 1864 14170
rect 4656 14118 4708 14170
rect 4720 14118 4772 14170
rect 4784 14118 4836 14170
rect 4848 14118 4900 14170
rect 4912 14118 4964 14170
rect 7756 14118 7808 14170
rect 7820 14118 7872 14170
rect 7884 14118 7936 14170
rect 7948 14118 8000 14170
rect 8012 14118 8064 14170
rect 10856 14118 10908 14170
rect 10920 14118 10972 14170
rect 10984 14118 11036 14170
rect 11048 14118 11100 14170
rect 11112 14118 11164 14170
rect 13956 14118 14008 14170
rect 14020 14118 14072 14170
rect 14084 14118 14136 14170
rect 14148 14118 14200 14170
rect 14212 14118 14264 14170
rect 17056 14118 17108 14170
rect 17120 14118 17172 14170
rect 17184 14118 17236 14170
rect 17248 14118 17300 14170
rect 17312 14118 17364 14170
rect 1952 14016 2004 14068
rect 5816 14016 5868 14068
rect 6644 14016 6696 14068
rect 8668 14016 8720 14068
rect 10140 14016 10192 14068
rect 11520 14016 11572 14068
rect 12256 13948 12308 14000
rect 2504 13923 2556 13932
rect 2504 13889 2513 13923
rect 2513 13889 2547 13923
rect 2547 13889 2556 13923
rect 2504 13880 2556 13889
rect 3792 13880 3844 13932
rect 2596 13812 2648 13864
rect 5080 13744 5132 13796
rect 6828 13812 6880 13864
rect 7104 13855 7156 13864
rect 7104 13821 7113 13855
rect 7113 13821 7147 13855
rect 7147 13821 7156 13855
rect 7104 13812 7156 13821
rect 8208 13880 8260 13932
rect 14280 13948 14332 14000
rect 15292 13948 15344 14000
rect 15568 13948 15620 14000
rect 18144 13948 18196 14000
rect 7472 13855 7524 13864
rect 7472 13821 7481 13855
rect 7481 13821 7515 13855
rect 7515 13821 7524 13855
rect 7472 13812 7524 13821
rect 11796 13855 11848 13864
rect 11796 13821 11805 13855
rect 11805 13821 11839 13855
rect 11839 13821 11848 13855
rect 11796 13812 11848 13821
rect 15200 13880 15252 13932
rect 12808 13855 12860 13864
rect 7196 13744 7248 13796
rect 6828 13676 6880 13728
rect 8484 13744 8536 13796
rect 8944 13744 8996 13796
rect 12808 13821 12817 13855
rect 12817 13821 12851 13855
rect 12851 13821 12860 13855
rect 12808 13812 12860 13821
rect 14832 13812 14884 13864
rect 14924 13812 14976 13864
rect 13728 13744 13780 13796
rect 13820 13744 13872 13796
rect 16304 13812 16356 13864
rect 16212 13787 16264 13796
rect 14740 13676 14792 13728
rect 16212 13753 16221 13787
rect 16221 13753 16255 13787
rect 16255 13753 16264 13787
rect 16948 13880 17000 13932
rect 17408 13855 17460 13864
rect 17408 13821 17416 13855
rect 17416 13821 17450 13855
rect 17450 13821 17460 13855
rect 17408 13812 17460 13821
rect 18236 13880 18288 13932
rect 19064 13812 19116 13864
rect 16212 13744 16264 13753
rect 16028 13676 16080 13728
rect 16856 13676 16908 13728
rect 3106 13574 3158 13626
rect 3170 13574 3222 13626
rect 3234 13574 3286 13626
rect 3298 13574 3350 13626
rect 3362 13574 3414 13626
rect 6206 13574 6258 13626
rect 6270 13574 6322 13626
rect 6334 13574 6386 13626
rect 6398 13574 6450 13626
rect 6462 13574 6514 13626
rect 9306 13574 9358 13626
rect 9370 13574 9422 13626
rect 9434 13574 9486 13626
rect 9498 13574 9550 13626
rect 9562 13574 9614 13626
rect 12406 13574 12458 13626
rect 12470 13574 12522 13626
rect 12534 13574 12586 13626
rect 12598 13574 12650 13626
rect 12662 13574 12714 13626
rect 15506 13574 15558 13626
rect 15570 13574 15622 13626
rect 15634 13574 15686 13626
rect 15698 13574 15750 13626
rect 15762 13574 15814 13626
rect 18606 13574 18658 13626
rect 18670 13574 18722 13626
rect 18734 13574 18786 13626
rect 18798 13574 18850 13626
rect 18862 13574 18914 13626
rect 8024 13472 8076 13524
rect 11244 13472 11296 13524
rect 13820 13472 13872 13524
rect 15200 13472 15252 13524
rect 4528 13404 4580 13456
rect 572 13268 624 13320
rect 3700 13379 3752 13388
rect 3700 13345 3734 13379
rect 3734 13345 3752 13379
rect 6092 13404 6144 13456
rect 5448 13379 5500 13388
rect 3700 13336 3752 13345
rect 5448 13345 5457 13379
rect 5457 13345 5491 13379
rect 5491 13345 5500 13379
rect 5448 13336 5500 13345
rect 6552 13404 6604 13456
rect 6828 13404 6880 13456
rect 11980 13447 12032 13456
rect 6644 13379 6696 13388
rect 6644 13345 6653 13379
rect 6653 13345 6687 13379
rect 6687 13345 6696 13379
rect 6644 13336 6696 13345
rect 6736 13336 6788 13388
rect 5724 13311 5776 13320
rect 5724 13277 5733 13311
rect 5733 13277 5767 13311
rect 5767 13277 5776 13311
rect 5724 13268 5776 13277
rect 6000 13268 6052 13320
rect 11980 13413 11989 13447
rect 11989 13413 12023 13447
rect 12023 13413 12032 13447
rect 11980 13404 12032 13413
rect 14648 13404 14700 13456
rect 14372 13379 14424 13388
rect 14372 13345 14381 13379
rect 14381 13345 14415 13379
rect 14415 13345 14424 13379
rect 14372 13336 14424 13345
rect 14740 13379 14792 13388
rect 14740 13345 14749 13379
rect 14749 13345 14783 13379
rect 14783 13345 14792 13379
rect 14740 13336 14792 13345
rect 14924 13336 14976 13388
rect 8852 13268 8904 13320
rect 9312 13268 9364 13320
rect 14832 13311 14884 13320
rect 14832 13277 14841 13311
rect 14841 13277 14875 13311
rect 14875 13277 14884 13311
rect 14832 13268 14884 13277
rect 15016 13268 15068 13320
rect 16212 13336 16264 13388
rect 16304 13268 16356 13320
rect 5080 13200 5132 13252
rect 6920 13243 6972 13252
rect 6920 13209 6929 13243
rect 6929 13209 6963 13243
rect 6963 13209 6972 13243
rect 6920 13200 6972 13209
rect 4988 13132 5040 13184
rect 5632 13175 5684 13184
rect 5632 13141 5641 13175
rect 5641 13141 5675 13175
rect 5675 13141 5684 13175
rect 5632 13132 5684 13141
rect 7656 13132 7708 13184
rect 16212 13132 16264 13184
rect 1556 13030 1608 13082
rect 1620 13030 1672 13082
rect 1684 13030 1736 13082
rect 1748 13030 1800 13082
rect 1812 13030 1864 13082
rect 4656 13030 4708 13082
rect 4720 13030 4772 13082
rect 4784 13030 4836 13082
rect 4848 13030 4900 13082
rect 4912 13030 4964 13082
rect 7756 13030 7808 13082
rect 7820 13030 7872 13082
rect 7884 13030 7936 13082
rect 7948 13030 8000 13082
rect 8012 13030 8064 13082
rect 10856 13030 10908 13082
rect 10920 13030 10972 13082
rect 10984 13030 11036 13082
rect 11048 13030 11100 13082
rect 11112 13030 11164 13082
rect 13956 13030 14008 13082
rect 14020 13030 14072 13082
rect 14084 13030 14136 13082
rect 14148 13030 14200 13082
rect 14212 13030 14264 13082
rect 17056 13030 17108 13082
rect 17120 13030 17172 13082
rect 17184 13030 17236 13082
rect 17248 13030 17300 13082
rect 17312 13030 17364 13082
rect 4988 12971 5040 12980
rect 4988 12937 4997 12971
rect 4997 12937 5031 12971
rect 5031 12937 5040 12971
rect 4988 12928 5040 12937
rect 7012 12928 7064 12980
rect 5448 12860 5500 12912
rect 7288 12792 7340 12844
rect 9036 12928 9088 12980
rect 12808 12928 12860 12980
rect 17960 12971 18012 12980
rect 17960 12937 17969 12971
rect 17969 12937 18003 12971
rect 18003 12937 18012 12971
rect 17960 12928 18012 12937
rect 9220 12792 9272 12844
rect 13820 12792 13872 12844
rect 5080 12724 5132 12776
rect 6000 12724 6052 12776
rect 6644 12767 6696 12776
rect 6644 12733 6653 12767
rect 6653 12733 6687 12767
rect 6687 12733 6696 12767
rect 6644 12724 6696 12733
rect 6920 12767 6972 12776
rect 6920 12733 6929 12767
rect 6929 12733 6963 12767
rect 6963 12733 6972 12767
rect 6920 12724 6972 12733
rect 7012 12724 7064 12776
rect 7196 12724 7248 12776
rect 8668 12724 8720 12776
rect 11152 12767 11204 12776
rect 11152 12733 11161 12767
rect 11161 12733 11195 12767
rect 11195 12733 11204 12767
rect 11152 12724 11204 12733
rect 11520 12767 11572 12776
rect 11520 12733 11529 12767
rect 11529 12733 11563 12767
rect 11563 12733 11572 12767
rect 11520 12724 11572 12733
rect 13728 12767 13780 12776
rect 13728 12733 13737 12767
rect 13737 12733 13771 12767
rect 13771 12733 13780 12767
rect 13728 12724 13780 12733
rect 16856 12792 16908 12844
rect 8944 12656 8996 12708
rect 9956 12656 10008 12708
rect 4344 12588 4396 12640
rect 6920 12588 6972 12640
rect 8668 12588 8720 12640
rect 11888 12656 11940 12708
rect 12900 12656 12952 12708
rect 16120 12724 16172 12776
rect 15200 12656 15252 12708
rect 12256 12588 12308 12640
rect 15292 12588 15344 12640
rect 16212 12588 16264 12640
rect 3106 12486 3158 12538
rect 3170 12486 3222 12538
rect 3234 12486 3286 12538
rect 3298 12486 3350 12538
rect 3362 12486 3414 12538
rect 6206 12486 6258 12538
rect 6270 12486 6322 12538
rect 6334 12486 6386 12538
rect 6398 12486 6450 12538
rect 6462 12486 6514 12538
rect 9306 12486 9358 12538
rect 9370 12486 9422 12538
rect 9434 12486 9486 12538
rect 9498 12486 9550 12538
rect 9562 12486 9614 12538
rect 12406 12486 12458 12538
rect 12470 12486 12522 12538
rect 12534 12486 12586 12538
rect 12598 12486 12650 12538
rect 12662 12486 12714 12538
rect 15506 12486 15558 12538
rect 15570 12486 15622 12538
rect 15634 12486 15686 12538
rect 15698 12486 15750 12538
rect 15762 12486 15814 12538
rect 18606 12486 18658 12538
rect 18670 12486 18722 12538
rect 18734 12486 18786 12538
rect 18798 12486 18850 12538
rect 18862 12486 18914 12538
rect 7564 12384 7616 12436
rect 11520 12384 11572 12436
rect 12256 12384 12308 12436
rect 16856 12384 16908 12436
rect 17960 12384 18012 12436
rect 18512 12384 18564 12436
rect 572 12248 624 12300
rect 1124 12248 1176 12300
rect 2228 12248 2280 12300
rect 2596 12248 2648 12300
rect 8576 12316 8628 12368
rect 11152 12316 11204 12368
rect 2412 12155 2464 12164
rect 2412 12121 2421 12155
rect 2421 12121 2455 12155
rect 2455 12121 2464 12155
rect 2964 12248 3016 12300
rect 3516 12248 3568 12300
rect 7196 12248 7248 12300
rect 10600 12291 10652 12300
rect 10600 12257 10609 12291
rect 10609 12257 10643 12291
rect 10643 12257 10652 12291
rect 10600 12248 10652 12257
rect 10784 12291 10836 12300
rect 10784 12257 10793 12291
rect 10793 12257 10827 12291
rect 10827 12257 10836 12291
rect 10784 12248 10836 12257
rect 13820 12316 13872 12368
rect 15108 12316 15160 12368
rect 12900 12248 12952 12300
rect 15016 12248 15068 12300
rect 15200 12291 15252 12300
rect 15200 12257 15209 12291
rect 15209 12257 15243 12291
rect 15243 12257 15252 12291
rect 15200 12248 15252 12257
rect 15292 12248 15344 12300
rect 5172 12223 5224 12232
rect 5172 12189 5181 12223
rect 5181 12189 5215 12223
rect 5215 12189 5224 12223
rect 5172 12180 5224 12189
rect 8576 12180 8628 12232
rect 2412 12112 2464 12121
rect 3700 12087 3752 12096
rect 3700 12053 3709 12087
rect 3709 12053 3743 12087
rect 3743 12053 3752 12087
rect 3700 12044 3752 12053
rect 7564 12044 7616 12096
rect 14648 12180 14700 12232
rect 13820 12155 13872 12164
rect 13820 12121 13829 12155
rect 13829 12121 13863 12155
rect 13863 12121 13872 12155
rect 13820 12112 13872 12121
rect 14280 12112 14332 12164
rect 16580 12223 16632 12232
rect 16580 12189 16589 12223
rect 16589 12189 16623 12223
rect 16623 12189 16632 12223
rect 16580 12180 16632 12189
rect 11612 12044 11664 12096
rect 16948 12044 17000 12096
rect 1556 11942 1608 11994
rect 1620 11942 1672 11994
rect 1684 11942 1736 11994
rect 1748 11942 1800 11994
rect 1812 11942 1864 11994
rect 4656 11942 4708 11994
rect 4720 11942 4772 11994
rect 4784 11942 4836 11994
rect 4848 11942 4900 11994
rect 4912 11942 4964 11994
rect 7756 11942 7808 11994
rect 7820 11942 7872 11994
rect 7884 11942 7936 11994
rect 7948 11942 8000 11994
rect 8012 11942 8064 11994
rect 10856 11942 10908 11994
rect 10920 11942 10972 11994
rect 10984 11942 11036 11994
rect 11048 11942 11100 11994
rect 11112 11942 11164 11994
rect 13956 11942 14008 11994
rect 14020 11942 14072 11994
rect 14084 11942 14136 11994
rect 14148 11942 14200 11994
rect 14212 11942 14264 11994
rect 17056 11942 17108 11994
rect 17120 11942 17172 11994
rect 17184 11942 17236 11994
rect 17248 11942 17300 11994
rect 17312 11942 17364 11994
rect 4160 11840 4212 11892
rect 5540 11883 5592 11892
rect 3516 11772 3568 11824
rect 5540 11849 5549 11883
rect 5549 11849 5583 11883
rect 5583 11849 5592 11883
rect 5540 11840 5592 11849
rect 5724 11840 5776 11892
rect 7104 11883 7156 11892
rect 7104 11849 7113 11883
rect 7113 11849 7147 11883
rect 7147 11849 7156 11883
rect 7104 11840 7156 11849
rect 7196 11840 7248 11892
rect 15384 11840 15436 11892
rect 4528 11772 4580 11824
rect 5264 11704 5316 11756
rect 2228 11679 2280 11688
rect 2228 11645 2237 11679
rect 2237 11645 2271 11679
rect 2271 11645 2280 11679
rect 2228 11636 2280 11645
rect 2412 11679 2464 11688
rect 2412 11645 2425 11679
rect 2425 11645 2464 11679
rect 2412 11636 2464 11645
rect 4344 11636 4396 11688
rect 3700 11568 3752 11620
rect 5632 11636 5684 11688
rect 6552 11704 6604 11756
rect 10784 11772 10836 11824
rect 7656 11747 7708 11756
rect 7656 11713 7665 11747
rect 7665 11713 7699 11747
rect 7699 11713 7708 11747
rect 7656 11704 7708 11713
rect 8300 11704 8352 11756
rect 9220 11704 9272 11756
rect 6000 11679 6052 11688
rect 6000 11645 6009 11679
rect 6009 11645 6043 11679
rect 6043 11645 6052 11679
rect 6000 11636 6052 11645
rect 6552 11611 6604 11620
rect 6552 11577 6561 11611
rect 6561 11577 6595 11611
rect 6595 11577 6604 11611
rect 6552 11568 6604 11577
rect 7380 11636 7432 11688
rect 11336 11679 11388 11688
rect 11336 11645 11345 11679
rect 11345 11645 11379 11679
rect 11379 11645 11388 11679
rect 11336 11636 11388 11645
rect 11704 11772 11756 11824
rect 11796 11704 11848 11756
rect 11612 11679 11664 11688
rect 11612 11645 11621 11679
rect 11621 11645 11655 11679
rect 11655 11645 11664 11679
rect 11612 11636 11664 11645
rect 15108 11636 15160 11688
rect 4988 11500 5040 11552
rect 5448 11500 5500 11552
rect 6092 11500 6144 11552
rect 8668 11568 8720 11620
rect 8944 11568 8996 11620
rect 18236 11840 18288 11892
rect 16120 11747 16172 11756
rect 16120 11713 16129 11747
rect 16129 11713 16163 11747
rect 16163 11713 16172 11747
rect 16120 11704 16172 11713
rect 17960 11704 18012 11756
rect 16488 11679 16540 11688
rect 16488 11645 16497 11679
rect 16497 11645 16531 11679
rect 16531 11645 16540 11679
rect 16488 11636 16540 11645
rect 16856 11568 16908 11620
rect 9956 11500 10008 11552
rect 14372 11500 14424 11552
rect 17316 11500 17368 11552
rect 3106 11398 3158 11450
rect 3170 11398 3222 11450
rect 3234 11398 3286 11450
rect 3298 11398 3350 11450
rect 3362 11398 3414 11450
rect 6206 11398 6258 11450
rect 6270 11398 6322 11450
rect 6334 11398 6386 11450
rect 6398 11398 6450 11450
rect 6462 11398 6514 11450
rect 9306 11398 9358 11450
rect 9370 11398 9422 11450
rect 9434 11398 9486 11450
rect 9498 11398 9550 11450
rect 9562 11398 9614 11450
rect 12406 11398 12458 11450
rect 12470 11398 12522 11450
rect 12534 11398 12586 11450
rect 12598 11398 12650 11450
rect 12662 11398 12714 11450
rect 15506 11398 15558 11450
rect 15570 11398 15622 11450
rect 15634 11398 15686 11450
rect 15698 11398 15750 11450
rect 15762 11398 15814 11450
rect 18606 11398 18658 11450
rect 18670 11398 18722 11450
rect 18734 11398 18786 11450
rect 18798 11398 18850 11450
rect 18862 11398 18914 11450
rect 2964 11296 3016 11348
rect 6920 11339 6972 11348
rect 6920 11305 6929 11339
rect 6929 11305 6963 11339
rect 6963 11305 6972 11339
rect 6920 11296 6972 11305
rect 8300 11339 8352 11348
rect 8300 11305 8309 11339
rect 8309 11305 8343 11339
rect 8343 11305 8352 11339
rect 8300 11296 8352 11305
rect 10600 11296 10652 11348
rect 15200 11339 15252 11348
rect 15200 11305 15209 11339
rect 15209 11305 15243 11339
rect 15243 11305 15252 11339
rect 15200 11296 15252 11305
rect 16028 11296 16080 11348
rect 16488 11296 16540 11348
rect 16672 11296 16724 11348
rect 18052 11296 18104 11348
rect 1124 11228 1176 11280
rect 5448 11271 5500 11280
rect 5448 11237 5457 11271
rect 5457 11237 5491 11271
rect 5491 11237 5500 11271
rect 5448 11228 5500 11237
rect 6736 11228 6788 11280
rect 10324 11228 10376 11280
rect 2136 11160 2188 11212
rect 2780 11160 2832 11212
rect 4528 11160 4580 11212
rect 11612 11228 11664 11280
rect 11336 11160 11388 11212
rect 11796 11160 11848 11212
rect 13728 11160 13780 11212
rect 2964 11024 3016 11076
rect 3516 11024 3568 11076
rect 11704 11092 11756 11144
rect 14832 11160 14884 11212
rect 16764 11228 16816 11280
rect 17316 11160 17368 11212
rect 17500 11203 17552 11212
rect 17500 11169 17509 11203
rect 17509 11169 17543 11203
rect 17543 11169 17552 11203
rect 17500 11160 17552 11169
rect 18420 11203 18472 11212
rect 18420 11169 18429 11203
rect 18429 11169 18463 11203
rect 18463 11169 18472 11203
rect 18420 11160 18472 11169
rect 2228 10956 2280 11008
rect 4988 10956 5040 11008
rect 12808 11024 12860 11076
rect 5632 10956 5684 11008
rect 12440 10956 12492 11008
rect 13452 10956 13504 11008
rect 15200 11092 15252 11144
rect 15108 11024 15160 11076
rect 15936 11067 15988 11076
rect 15936 11033 15945 11067
rect 15945 11033 15979 11067
rect 15979 11033 15988 11067
rect 15936 11024 15988 11033
rect 16764 10956 16816 11008
rect 1556 10854 1608 10906
rect 1620 10854 1672 10906
rect 1684 10854 1736 10906
rect 1748 10854 1800 10906
rect 1812 10854 1864 10906
rect 4656 10854 4708 10906
rect 4720 10854 4772 10906
rect 4784 10854 4836 10906
rect 4848 10854 4900 10906
rect 4912 10854 4964 10906
rect 7756 10854 7808 10906
rect 7820 10854 7872 10906
rect 7884 10854 7936 10906
rect 7948 10854 8000 10906
rect 8012 10854 8064 10906
rect 10856 10854 10908 10906
rect 10920 10854 10972 10906
rect 10984 10854 11036 10906
rect 11048 10854 11100 10906
rect 11112 10854 11164 10906
rect 13956 10854 14008 10906
rect 14020 10854 14072 10906
rect 14084 10854 14136 10906
rect 14148 10854 14200 10906
rect 14212 10854 14264 10906
rect 17056 10854 17108 10906
rect 17120 10854 17172 10906
rect 17184 10854 17236 10906
rect 17248 10854 17300 10906
rect 17312 10854 17364 10906
rect 4344 10752 4396 10804
rect 6552 10752 6604 10804
rect 12808 10752 12860 10804
rect 13452 10752 13504 10804
rect 15936 10752 15988 10804
rect 16672 10752 16724 10804
rect 17500 10752 17552 10804
rect 17684 10752 17736 10804
rect 4160 10684 4212 10736
rect 5264 10727 5316 10736
rect 5264 10693 5273 10727
rect 5273 10693 5307 10727
rect 5307 10693 5316 10727
rect 5264 10684 5316 10693
rect 14832 10727 14884 10736
rect 14832 10693 14841 10727
rect 14841 10693 14875 10727
rect 14875 10693 14884 10727
rect 14832 10684 14884 10693
rect 1124 10591 1176 10600
rect 1124 10557 1133 10591
rect 1133 10557 1167 10591
rect 1167 10557 1176 10591
rect 1124 10548 1176 10557
rect 1952 10591 2004 10600
rect 1952 10557 1961 10591
rect 1961 10557 1995 10591
rect 1995 10557 2004 10591
rect 1952 10548 2004 10557
rect 4068 10548 4120 10600
rect 4620 10548 4672 10600
rect 2320 10480 2372 10532
rect 4344 10480 4396 10532
rect 14280 10616 14332 10668
rect 16120 10616 16172 10668
rect 10048 10548 10100 10600
rect 12440 10591 12492 10600
rect 12440 10557 12449 10591
rect 12449 10557 12483 10591
rect 12483 10557 12492 10591
rect 12440 10548 12492 10557
rect 13084 10548 13136 10600
rect 14464 10591 14516 10600
rect 14464 10557 14473 10591
rect 14473 10557 14507 10591
rect 14507 10557 14516 10591
rect 14464 10548 14516 10557
rect 2780 10412 2832 10464
rect 4988 10480 5040 10532
rect 10508 10480 10560 10532
rect 16488 10523 16540 10532
rect 10140 10412 10192 10464
rect 12256 10412 12308 10464
rect 16488 10489 16497 10523
rect 16497 10489 16531 10523
rect 16531 10489 16540 10523
rect 16488 10480 16540 10489
rect 16028 10412 16080 10464
rect 16212 10412 16264 10464
rect 3106 10310 3158 10362
rect 3170 10310 3222 10362
rect 3234 10310 3286 10362
rect 3298 10310 3350 10362
rect 3362 10310 3414 10362
rect 6206 10310 6258 10362
rect 6270 10310 6322 10362
rect 6334 10310 6386 10362
rect 6398 10310 6450 10362
rect 6462 10310 6514 10362
rect 9306 10310 9358 10362
rect 9370 10310 9422 10362
rect 9434 10310 9486 10362
rect 9498 10310 9550 10362
rect 9562 10310 9614 10362
rect 12406 10310 12458 10362
rect 12470 10310 12522 10362
rect 12534 10310 12586 10362
rect 12598 10310 12650 10362
rect 12662 10310 12714 10362
rect 15506 10310 15558 10362
rect 15570 10310 15622 10362
rect 15634 10310 15686 10362
rect 15698 10310 15750 10362
rect 15762 10310 15814 10362
rect 18606 10310 18658 10362
rect 18670 10310 18722 10362
rect 18734 10310 18786 10362
rect 18798 10310 18850 10362
rect 18862 10310 18914 10362
rect 1952 10208 2004 10260
rect 6644 10208 6696 10260
rect 7012 10208 7064 10260
rect 12256 10208 12308 10260
rect 13084 10251 13136 10260
rect 13084 10217 13093 10251
rect 13093 10217 13127 10251
rect 13127 10217 13136 10251
rect 13084 10208 13136 10217
rect 16488 10208 16540 10260
rect 1124 10140 1176 10192
rect 4528 10183 4580 10192
rect 4528 10149 4537 10183
rect 4537 10149 4571 10183
rect 4571 10149 4580 10183
rect 4528 10140 4580 10149
rect 5172 10140 5224 10192
rect 8484 10140 8536 10192
rect 11428 10140 11480 10192
rect 2872 10072 2924 10124
rect 7012 10115 7064 10124
rect 2228 10047 2280 10056
rect 2228 10013 2237 10047
rect 2237 10013 2271 10047
rect 2271 10013 2280 10047
rect 2228 10004 2280 10013
rect 7012 10081 7021 10115
rect 7021 10081 7055 10115
rect 7055 10081 7064 10115
rect 7012 10072 7064 10081
rect 7564 10115 7616 10124
rect 7564 10081 7573 10115
rect 7573 10081 7607 10115
rect 7607 10081 7616 10115
rect 7564 10072 7616 10081
rect 10140 10115 10192 10124
rect 10140 10081 10149 10115
rect 10149 10081 10183 10115
rect 10183 10081 10192 10115
rect 10140 10072 10192 10081
rect 10508 10115 10560 10124
rect 10508 10081 10517 10115
rect 10517 10081 10551 10115
rect 10551 10081 10560 10115
rect 10508 10072 10560 10081
rect 12900 10140 12952 10192
rect 12808 10115 12860 10124
rect 12808 10081 12817 10115
rect 12817 10081 12851 10115
rect 12851 10081 12860 10115
rect 16948 10140 17000 10192
rect 12808 10072 12860 10081
rect 6828 10047 6880 10056
rect 6828 10013 6837 10047
rect 6837 10013 6871 10047
rect 6871 10013 6880 10047
rect 6828 10004 6880 10013
rect 8300 10004 8352 10056
rect 14464 10072 14516 10124
rect 17316 10115 17368 10124
rect 17316 10081 17345 10115
rect 17345 10081 17368 10115
rect 17316 10072 17368 10081
rect 17684 10115 17736 10124
rect 17684 10081 17693 10115
rect 17693 10081 17727 10115
rect 17727 10081 17736 10115
rect 17684 10072 17736 10081
rect 2780 9936 2832 9988
rect 11336 9936 11388 9988
rect 16580 9936 16632 9988
rect 17592 9979 17644 9988
rect 17592 9945 17601 9979
rect 17601 9945 17635 9979
rect 17635 9945 17644 9979
rect 17592 9936 17644 9945
rect 9036 9868 9088 9920
rect 12348 9868 12400 9920
rect 16028 9911 16080 9920
rect 16028 9877 16037 9911
rect 16037 9877 16071 9911
rect 16071 9877 16080 9911
rect 16028 9868 16080 9877
rect 1556 9766 1608 9818
rect 1620 9766 1672 9818
rect 1684 9766 1736 9818
rect 1748 9766 1800 9818
rect 1812 9766 1864 9818
rect 4656 9766 4708 9818
rect 4720 9766 4772 9818
rect 4784 9766 4836 9818
rect 4848 9766 4900 9818
rect 4912 9766 4964 9818
rect 7756 9766 7808 9818
rect 7820 9766 7872 9818
rect 7884 9766 7936 9818
rect 7948 9766 8000 9818
rect 8012 9766 8064 9818
rect 10856 9766 10908 9818
rect 10920 9766 10972 9818
rect 10984 9766 11036 9818
rect 11048 9766 11100 9818
rect 11112 9766 11164 9818
rect 13956 9766 14008 9818
rect 14020 9766 14072 9818
rect 14084 9766 14136 9818
rect 14148 9766 14200 9818
rect 14212 9766 14264 9818
rect 17056 9766 17108 9818
rect 17120 9766 17172 9818
rect 17184 9766 17236 9818
rect 17248 9766 17300 9818
rect 17312 9766 17364 9818
rect 2872 9639 2924 9648
rect 2872 9605 2881 9639
rect 2881 9605 2915 9639
rect 2915 9605 2924 9639
rect 2872 9596 2924 9605
rect 8300 9639 8352 9648
rect 8300 9605 8309 9639
rect 8309 9605 8343 9639
rect 8343 9605 8352 9639
rect 8300 9596 8352 9605
rect 4252 9528 4304 9580
rect 7012 9528 7064 9580
rect 2412 9460 2464 9512
rect 3516 9460 3568 9512
rect 7564 9460 7616 9512
rect 9036 9503 9088 9512
rect 2136 9324 2188 9376
rect 4160 9392 4212 9444
rect 2320 9324 2372 9376
rect 4988 9324 5040 9376
rect 5264 9324 5316 9376
rect 9036 9469 9045 9503
rect 9045 9469 9079 9503
rect 9079 9469 9088 9503
rect 9036 9460 9088 9469
rect 14280 9503 14332 9512
rect 14280 9469 14289 9503
rect 14289 9469 14323 9503
rect 14323 9469 14332 9503
rect 14280 9460 14332 9469
rect 14648 9503 14700 9512
rect 14648 9469 14657 9503
rect 14657 9469 14691 9503
rect 14691 9469 14700 9503
rect 14648 9460 14700 9469
rect 8300 9392 8352 9444
rect 14464 9392 14516 9444
rect 9036 9324 9088 9376
rect 11428 9324 11480 9376
rect 11796 9324 11848 9376
rect 12348 9324 12400 9376
rect 15108 9324 15160 9376
rect 3106 9222 3158 9274
rect 3170 9222 3222 9274
rect 3234 9222 3286 9274
rect 3298 9222 3350 9274
rect 3362 9222 3414 9274
rect 6206 9222 6258 9274
rect 6270 9222 6322 9274
rect 6334 9222 6386 9274
rect 6398 9222 6450 9274
rect 6462 9222 6514 9274
rect 9306 9222 9358 9274
rect 9370 9222 9422 9274
rect 9434 9222 9486 9274
rect 9498 9222 9550 9274
rect 9562 9222 9614 9274
rect 12406 9222 12458 9274
rect 12470 9222 12522 9274
rect 12534 9222 12586 9274
rect 12598 9222 12650 9274
rect 12662 9222 12714 9274
rect 15506 9222 15558 9274
rect 15570 9222 15622 9274
rect 15634 9222 15686 9274
rect 15698 9222 15750 9274
rect 15762 9222 15814 9274
rect 18606 9222 18658 9274
rect 18670 9222 18722 9274
rect 18734 9222 18786 9274
rect 18798 9222 18850 9274
rect 18862 9222 18914 9274
rect 4436 9120 4488 9172
rect 5632 9120 5684 9172
rect 14648 9120 14700 9172
rect 8484 9052 8536 9104
rect 11796 9052 11848 9104
rect 2320 8984 2372 9036
rect 3976 8984 4028 9036
rect 4344 9027 4396 9036
rect 4344 8993 4353 9027
rect 4353 8993 4387 9027
rect 4387 8993 4396 9027
rect 4344 8984 4396 8993
rect 5080 8984 5132 9036
rect 5264 9027 5316 9036
rect 5264 8993 5273 9027
rect 5273 8993 5307 9027
rect 5307 8993 5316 9027
rect 5264 8984 5316 8993
rect 12900 9052 12952 9104
rect 14464 9052 14516 9104
rect 2228 8916 2280 8968
rect 2412 8916 2464 8968
rect 4252 8916 4304 8968
rect 4988 8916 5040 8968
rect 5632 8959 5684 8968
rect 5632 8925 5641 8959
rect 5641 8925 5675 8959
rect 5675 8925 5684 8959
rect 5632 8916 5684 8925
rect 848 8780 900 8832
rect 5172 8780 5224 8832
rect 5908 8780 5960 8832
rect 6828 8780 6880 8832
rect 10048 8780 10100 8832
rect 11244 8916 11296 8968
rect 12808 8984 12860 9036
rect 13728 8984 13780 9036
rect 14648 8984 14700 9036
rect 12808 8848 12860 8900
rect 14280 8891 14332 8900
rect 14280 8857 14289 8891
rect 14289 8857 14323 8891
rect 14323 8857 14332 8891
rect 14280 8848 14332 8857
rect 17408 9120 17460 9172
rect 18236 9163 18288 9172
rect 18236 9129 18245 9163
rect 18245 9129 18279 9163
rect 18279 9129 18288 9163
rect 18236 9120 18288 9129
rect 17500 9052 17552 9104
rect 15108 8891 15160 8900
rect 15108 8857 15117 8891
rect 15117 8857 15151 8891
rect 15151 8857 15160 8891
rect 15108 8848 15160 8857
rect 16304 8984 16356 9036
rect 17960 8984 18012 9036
rect 18420 9027 18472 9036
rect 18420 8993 18429 9027
rect 18429 8993 18463 9027
rect 18463 8993 18472 9027
rect 18420 8984 18472 8993
rect 12072 8780 12124 8832
rect 14464 8780 14516 8832
rect 18420 8848 18472 8900
rect 15568 8823 15620 8832
rect 15568 8789 15577 8823
rect 15577 8789 15611 8823
rect 15611 8789 15620 8823
rect 15568 8780 15620 8789
rect 1556 8678 1608 8730
rect 1620 8678 1672 8730
rect 1684 8678 1736 8730
rect 1748 8678 1800 8730
rect 1812 8678 1864 8730
rect 4656 8678 4708 8730
rect 4720 8678 4772 8730
rect 4784 8678 4836 8730
rect 4848 8678 4900 8730
rect 4912 8678 4964 8730
rect 7756 8678 7808 8730
rect 7820 8678 7872 8730
rect 7884 8678 7936 8730
rect 7948 8678 8000 8730
rect 8012 8678 8064 8730
rect 10856 8678 10908 8730
rect 10920 8678 10972 8730
rect 10984 8678 11036 8730
rect 11048 8678 11100 8730
rect 11112 8678 11164 8730
rect 13956 8678 14008 8730
rect 14020 8678 14072 8730
rect 14084 8678 14136 8730
rect 14148 8678 14200 8730
rect 14212 8678 14264 8730
rect 17056 8678 17108 8730
rect 17120 8678 17172 8730
rect 17184 8678 17236 8730
rect 17248 8678 17300 8730
rect 17312 8678 17364 8730
rect 2964 8576 3016 8628
rect 3976 8619 4028 8628
rect 3976 8585 3985 8619
rect 3985 8585 4019 8619
rect 4019 8585 4028 8619
rect 3976 8576 4028 8585
rect 5172 8576 5224 8628
rect 5632 8576 5684 8628
rect 11244 8619 11296 8628
rect 11244 8585 11253 8619
rect 11253 8585 11287 8619
rect 11287 8585 11296 8619
rect 11244 8576 11296 8585
rect 14280 8576 14332 8628
rect 15568 8576 15620 8628
rect 17960 8619 18012 8628
rect 17960 8585 17969 8619
rect 17969 8585 18003 8619
rect 18003 8585 18012 8619
rect 17960 8576 18012 8585
rect 14556 8551 14608 8560
rect 2780 8440 2832 8492
rect 3976 8440 4028 8492
rect 12072 8440 12124 8492
rect 4436 8415 4488 8424
rect 2320 8304 2372 8356
rect 4436 8381 4445 8415
rect 4445 8381 4479 8415
rect 4479 8381 4488 8415
rect 4436 8372 4488 8381
rect 5264 8415 5316 8424
rect 5264 8381 5273 8415
rect 5273 8381 5307 8415
rect 5307 8381 5316 8415
rect 5264 8372 5316 8381
rect 5632 8372 5684 8424
rect 6828 8415 6880 8424
rect 6828 8381 6837 8415
rect 6837 8381 6871 8415
rect 6871 8381 6880 8415
rect 6828 8372 6880 8381
rect 11336 8415 11388 8424
rect 11336 8381 11345 8415
rect 11345 8381 11379 8415
rect 11379 8381 11388 8415
rect 11336 8372 11388 8381
rect 14556 8517 14565 8551
rect 14565 8517 14599 8551
rect 14599 8517 14608 8551
rect 14556 8508 14608 8517
rect 16304 8551 16356 8560
rect 16304 8517 16313 8551
rect 16313 8517 16347 8551
rect 16347 8517 16356 8551
rect 16304 8508 16356 8517
rect 13728 8440 13780 8492
rect 16212 8440 16264 8492
rect 5816 8304 5868 8356
rect 15292 8304 15344 8356
rect 16396 8372 16448 8424
rect 17224 8372 17276 8424
rect 4344 8279 4396 8288
rect 4344 8245 4353 8279
rect 4353 8245 4387 8279
rect 4387 8245 4396 8279
rect 4344 8236 4396 8245
rect 13912 8279 13964 8288
rect 13912 8245 13921 8279
rect 13921 8245 13955 8279
rect 13955 8245 13964 8279
rect 13912 8236 13964 8245
rect 16672 8304 16724 8356
rect 3106 8134 3158 8186
rect 3170 8134 3222 8186
rect 3234 8134 3286 8186
rect 3298 8134 3350 8186
rect 3362 8134 3414 8186
rect 6206 8134 6258 8186
rect 6270 8134 6322 8186
rect 6334 8134 6386 8186
rect 6398 8134 6450 8186
rect 6462 8134 6514 8186
rect 9306 8134 9358 8186
rect 9370 8134 9422 8186
rect 9434 8134 9486 8186
rect 9498 8134 9550 8186
rect 9562 8134 9614 8186
rect 12406 8134 12458 8186
rect 12470 8134 12522 8186
rect 12534 8134 12586 8186
rect 12598 8134 12650 8186
rect 12662 8134 12714 8186
rect 15506 8134 15558 8186
rect 15570 8134 15622 8186
rect 15634 8134 15686 8186
rect 15698 8134 15750 8186
rect 15762 8134 15814 8186
rect 18606 8134 18658 8186
rect 18670 8134 18722 8186
rect 18734 8134 18786 8186
rect 18798 8134 18850 8186
rect 18862 8134 18914 8186
rect 848 8007 900 8016
rect 848 7973 857 8007
rect 857 7973 891 8007
rect 891 7973 900 8007
rect 848 7964 900 7973
rect 2136 7964 2188 8016
rect 572 7939 624 7948
rect 572 7905 581 7939
rect 581 7905 615 7939
rect 615 7905 624 7939
rect 572 7896 624 7905
rect 5264 8032 5316 8084
rect 13912 8032 13964 8084
rect 15108 8075 15160 8084
rect 15108 8041 15117 8075
rect 15117 8041 15151 8075
rect 15151 8041 15160 8075
rect 15108 8032 15160 8041
rect 17500 8075 17552 8084
rect 17500 8041 17509 8075
rect 17509 8041 17543 8075
rect 17543 8041 17552 8075
rect 17500 8032 17552 8041
rect 4528 8007 4580 8016
rect 4528 7973 4537 8007
rect 4537 7973 4571 8007
rect 4571 7973 4580 8007
rect 4528 7964 4580 7973
rect 8484 7964 8536 8016
rect 7564 7939 7616 7948
rect 7564 7905 7573 7939
rect 7573 7905 7607 7939
rect 7607 7905 7616 7939
rect 7564 7896 7616 7905
rect 11244 7964 11296 8016
rect 12808 8007 12860 8016
rect 12808 7973 12817 8007
rect 12817 7973 12851 8007
rect 12851 7973 12860 8007
rect 12808 7964 12860 7973
rect 14372 8007 14424 8016
rect 14372 7973 14381 8007
rect 14381 7973 14415 8007
rect 14415 7973 14424 8007
rect 14372 7964 14424 7973
rect 14556 7964 14608 8016
rect 10784 7939 10836 7948
rect 10784 7905 10793 7939
rect 10793 7905 10827 7939
rect 10827 7905 10836 7939
rect 10784 7896 10836 7905
rect 12440 7896 12492 7948
rect 13728 7896 13780 7948
rect 16672 7896 16724 7948
rect 17224 7939 17276 7948
rect 17224 7905 17234 7939
rect 17234 7905 17268 7939
rect 17268 7905 17276 7939
rect 17224 7896 17276 7905
rect 2320 7871 2372 7880
rect 2320 7837 2329 7871
rect 2329 7837 2363 7871
rect 2363 7837 2372 7871
rect 2320 7828 2372 7837
rect 5540 7871 5592 7880
rect 5540 7837 5549 7871
rect 5549 7837 5583 7871
rect 5583 7837 5592 7871
rect 5540 7828 5592 7837
rect 5264 7760 5316 7812
rect 4068 7692 4120 7744
rect 5816 7871 5868 7880
rect 5816 7837 5825 7871
rect 5825 7837 5859 7871
rect 5859 7837 5868 7871
rect 5816 7828 5868 7837
rect 8208 7828 8260 7880
rect 15016 7828 15068 7880
rect 11336 7760 11388 7812
rect 8668 7692 8720 7744
rect 9312 7735 9364 7744
rect 9312 7701 9321 7735
rect 9321 7701 9355 7735
rect 9355 7701 9364 7735
rect 9312 7692 9364 7701
rect 1556 7590 1608 7642
rect 1620 7590 1672 7642
rect 1684 7590 1736 7642
rect 1748 7590 1800 7642
rect 1812 7590 1864 7642
rect 4656 7590 4708 7642
rect 4720 7590 4772 7642
rect 4784 7590 4836 7642
rect 4848 7590 4900 7642
rect 4912 7590 4964 7642
rect 7756 7590 7808 7642
rect 7820 7590 7872 7642
rect 7884 7590 7936 7642
rect 7948 7590 8000 7642
rect 8012 7590 8064 7642
rect 10856 7590 10908 7642
rect 10920 7590 10972 7642
rect 10984 7590 11036 7642
rect 11048 7590 11100 7642
rect 11112 7590 11164 7642
rect 13956 7590 14008 7642
rect 14020 7590 14072 7642
rect 14084 7590 14136 7642
rect 14148 7590 14200 7642
rect 14212 7590 14264 7642
rect 17056 7590 17108 7642
rect 17120 7590 17172 7642
rect 17184 7590 17236 7642
rect 17248 7590 17300 7642
rect 17312 7590 17364 7642
rect 4344 7488 4396 7540
rect 5632 7531 5684 7540
rect 5632 7497 5641 7531
rect 5641 7497 5675 7531
rect 5675 7497 5684 7531
rect 5632 7488 5684 7497
rect 11336 7531 11388 7540
rect 11336 7497 11345 7531
rect 11345 7497 11379 7531
rect 11379 7497 11388 7531
rect 11336 7488 11388 7497
rect 13728 7488 13780 7540
rect 9036 7463 9088 7472
rect 9036 7429 9045 7463
rect 9045 7429 9079 7463
rect 9079 7429 9088 7463
rect 9036 7420 9088 7429
rect 2412 7352 2464 7404
rect 4068 7352 4120 7404
rect 5816 7352 5868 7404
rect 2964 7284 3016 7336
rect 3976 7327 4028 7336
rect 3976 7293 3985 7327
rect 3985 7293 4019 7327
rect 4019 7293 4028 7327
rect 3976 7284 4028 7293
rect 2320 7216 2372 7268
rect 5908 7284 5960 7336
rect 6828 7284 6880 7336
rect 8668 7352 8720 7404
rect 9312 7352 9364 7404
rect 7288 7284 7340 7336
rect 4436 7216 4488 7268
rect 5264 7259 5316 7268
rect 5264 7225 5273 7259
rect 5273 7225 5307 7259
rect 5307 7225 5316 7259
rect 5264 7216 5316 7225
rect 5448 7216 5500 7268
rect 8116 7284 8168 7336
rect 8300 7284 8352 7336
rect 8944 7284 8996 7336
rect 12900 7352 12952 7404
rect 12164 7327 12216 7336
rect 12164 7293 12173 7327
rect 12173 7293 12207 7327
rect 12207 7293 12216 7327
rect 12164 7284 12216 7293
rect 12440 7284 12492 7336
rect 16672 7488 16724 7540
rect 14372 7352 14424 7404
rect 15384 7352 15436 7404
rect 16396 7395 16448 7404
rect 16396 7361 16405 7395
rect 16405 7361 16439 7395
rect 16439 7361 16448 7395
rect 16396 7352 16448 7361
rect 15292 7284 15344 7336
rect 9220 7216 9272 7268
rect 15200 7216 15252 7268
rect 16304 7216 16356 7268
rect 848 7148 900 7200
rect 2780 7148 2832 7200
rect 7104 7191 7156 7200
rect 7104 7157 7113 7191
rect 7113 7157 7147 7191
rect 7147 7157 7156 7191
rect 7104 7148 7156 7157
rect 7656 7191 7708 7200
rect 7656 7157 7665 7191
rect 7665 7157 7699 7191
rect 7699 7157 7708 7191
rect 7656 7148 7708 7157
rect 8300 7191 8352 7200
rect 8300 7157 8309 7191
rect 8309 7157 8343 7191
rect 8343 7157 8352 7191
rect 8300 7148 8352 7157
rect 8944 7148 8996 7200
rect 9128 7191 9180 7200
rect 9128 7157 9137 7191
rect 9137 7157 9171 7191
rect 9171 7157 9180 7191
rect 9128 7148 9180 7157
rect 11152 7191 11204 7200
rect 11152 7157 11161 7191
rect 11161 7157 11195 7191
rect 11195 7157 11204 7191
rect 11152 7148 11204 7157
rect 14464 7191 14516 7200
rect 14464 7157 14473 7191
rect 14473 7157 14507 7191
rect 14507 7157 14516 7191
rect 14464 7148 14516 7157
rect 3106 7046 3158 7098
rect 3170 7046 3222 7098
rect 3234 7046 3286 7098
rect 3298 7046 3350 7098
rect 3362 7046 3414 7098
rect 6206 7046 6258 7098
rect 6270 7046 6322 7098
rect 6334 7046 6386 7098
rect 6398 7046 6450 7098
rect 6462 7046 6514 7098
rect 9306 7046 9358 7098
rect 9370 7046 9422 7098
rect 9434 7046 9486 7098
rect 9498 7046 9550 7098
rect 9562 7046 9614 7098
rect 12406 7046 12458 7098
rect 12470 7046 12522 7098
rect 12534 7046 12586 7098
rect 12598 7046 12650 7098
rect 12662 7046 12714 7098
rect 15506 7046 15558 7098
rect 15570 7046 15622 7098
rect 15634 7046 15686 7098
rect 15698 7046 15750 7098
rect 15762 7046 15814 7098
rect 18606 7046 18658 7098
rect 18670 7046 18722 7098
rect 18734 7046 18786 7098
rect 18798 7046 18850 7098
rect 18862 7046 18914 7098
rect 2136 6876 2188 6928
rect 2780 6987 2832 6996
rect 2780 6953 2789 6987
rect 2789 6953 2823 6987
rect 2823 6953 2832 6987
rect 2780 6944 2832 6953
rect 4344 6944 4396 6996
rect 8208 6987 8260 6996
rect 8208 6953 8217 6987
rect 8217 6953 8251 6987
rect 8251 6953 8260 6987
rect 8208 6944 8260 6953
rect 10784 6944 10836 6996
rect 11704 6944 11756 6996
rect 2964 6876 3016 6928
rect 572 6851 624 6860
rect 572 6817 581 6851
rect 581 6817 615 6851
rect 615 6817 624 6851
rect 572 6808 624 6817
rect 6644 6876 6696 6928
rect 848 6783 900 6792
rect 848 6749 857 6783
rect 857 6749 891 6783
rect 891 6749 900 6783
rect 848 6740 900 6749
rect 2228 6740 2280 6792
rect 3516 6740 3568 6792
rect 4344 6783 4396 6792
rect 4344 6749 4353 6783
rect 4353 6749 4387 6783
rect 4387 6749 4396 6783
rect 6828 6851 6880 6860
rect 6828 6817 6837 6851
rect 6837 6817 6871 6851
rect 6871 6817 6880 6851
rect 7104 6876 7156 6928
rect 6828 6808 6880 6817
rect 4344 6740 4396 6749
rect 7288 6740 7340 6792
rect 7472 6808 7524 6860
rect 11796 6876 11848 6928
rect 12072 6876 12124 6928
rect 7748 6740 7800 6792
rect 2412 6672 2464 6724
rect 9220 6808 9272 6860
rect 14464 6944 14516 6996
rect 10048 6740 10100 6792
rect 11152 6740 11204 6792
rect 12164 6740 12216 6792
rect 13452 6783 13504 6792
rect 8852 6672 8904 6724
rect 8576 6647 8628 6656
rect 8576 6613 8585 6647
rect 8585 6613 8619 6647
rect 8619 6613 8628 6647
rect 8576 6604 8628 6613
rect 8944 6647 8996 6656
rect 8944 6613 8953 6647
rect 8953 6613 8987 6647
rect 8987 6613 8996 6647
rect 8944 6604 8996 6613
rect 12900 6672 12952 6724
rect 13452 6749 13461 6783
rect 13461 6749 13495 6783
rect 13495 6749 13504 6783
rect 13452 6740 13504 6749
rect 15200 6944 15252 6996
rect 15016 6876 15068 6928
rect 15108 6851 15160 6860
rect 15108 6817 15117 6851
rect 15117 6817 15151 6851
rect 15151 6817 15160 6851
rect 15108 6808 15160 6817
rect 15200 6783 15252 6792
rect 15200 6749 15209 6783
rect 15209 6749 15243 6783
rect 15243 6749 15252 6783
rect 15200 6740 15252 6749
rect 15384 6808 15436 6860
rect 18420 6851 18472 6860
rect 18420 6817 18429 6851
rect 18429 6817 18463 6851
rect 18463 6817 18472 6851
rect 18420 6808 18472 6817
rect 16764 6604 16816 6656
rect 1556 6502 1608 6554
rect 1620 6502 1672 6554
rect 1684 6502 1736 6554
rect 1748 6502 1800 6554
rect 1812 6502 1864 6554
rect 4656 6502 4708 6554
rect 4720 6502 4772 6554
rect 4784 6502 4836 6554
rect 4848 6502 4900 6554
rect 4912 6502 4964 6554
rect 7756 6502 7808 6554
rect 7820 6502 7872 6554
rect 7884 6502 7936 6554
rect 7948 6502 8000 6554
rect 8012 6502 8064 6554
rect 10856 6502 10908 6554
rect 10920 6502 10972 6554
rect 10984 6502 11036 6554
rect 11048 6502 11100 6554
rect 11112 6502 11164 6554
rect 13956 6502 14008 6554
rect 14020 6502 14072 6554
rect 14084 6502 14136 6554
rect 14148 6502 14200 6554
rect 14212 6502 14264 6554
rect 17056 6502 17108 6554
rect 17120 6502 17172 6554
rect 17184 6502 17236 6554
rect 17248 6502 17300 6554
rect 17312 6502 17364 6554
rect 2228 6443 2280 6452
rect 2228 6409 2237 6443
rect 2237 6409 2271 6443
rect 2271 6409 2280 6443
rect 2228 6400 2280 6409
rect 4252 6264 4304 6316
rect 5172 6400 5224 6452
rect 6092 6400 6144 6452
rect 8944 6400 8996 6452
rect 13452 6400 13504 6452
rect 14556 6400 14608 6452
rect 15108 6400 15160 6452
rect 2228 6196 2280 6248
rect 4436 6239 4488 6248
rect 4436 6205 4445 6239
rect 4445 6205 4479 6239
rect 4479 6205 4488 6239
rect 4436 6196 4488 6205
rect 4988 6239 5040 6248
rect 4988 6205 4997 6239
rect 4997 6205 5031 6239
rect 5031 6205 5040 6239
rect 4988 6196 5040 6205
rect 5080 6196 5132 6248
rect 5448 6239 5500 6248
rect 5448 6205 5457 6239
rect 5457 6205 5491 6239
rect 5491 6205 5500 6239
rect 5448 6196 5500 6205
rect 8300 6332 8352 6384
rect 8760 6264 8812 6316
rect 12164 6264 12216 6316
rect 14280 6264 14332 6316
rect 7656 6196 7708 6248
rect 8576 6196 8628 6248
rect 12900 6196 12952 6248
rect 16396 6264 16448 6316
rect 16488 6239 16540 6248
rect 16488 6205 16497 6239
rect 16497 6205 16531 6239
rect 16531 6205 16540 6239
rect 16488 6196 16540 6205
rect 6644 6128 6696 6180
rect 6828 6128 6880 6180
rect 16028 6128 16080 6180
rect 17500 6128 17552 6180
rect 17960 6171 18012 6180
rect 17960 6137 17969 6171
rect 17969 6137 18003 6171
rect 18003 6137 18012 6171
rect 17960 6128 18012 6137
rect 8024 6060 8076 6112
rect 12072 6103 12124 6112
rect 12072 6069 12081 6103
rect 12081 6069 12115 6103
rect 12115 6069 12124 6103
rect 12072 6060 12124 6069
rect 13268 6060 13320 6112
rect 14556 6060 14608 6112
rect 16948 6060 17000 6112
rect 3106 5958 3158 6010
rect 3170 5958 3222 6010
rect 3234 5958 3286 6010
rect 3298 5958 3350 6010
rect 3362 5958 3414 6010
rect 6206 5958 6258 6010
rect 6270 5958 6322 6010
rect 6334 5958 6386 6010
rect 6398 5958 6450 6010
rect 6462 5958 6514 6010
rect 9306 5958 9358 6010
rect 9370 5958 9422 6010
rect 9434 5958 9486 6010
rect 9498 5958 9550 6010
rect 9562 5958 9614 6010
rect 12406 5958 12458 6010
rect 12470 5958 12522 6010
rect 12534 5958 12586 6010
rect 12598 5958 12650 6010
rect 12662 5958 12714 6010
rect 15506 5958 15558 6010
rect 15570 5958 15622 6010
rect 15634 5958 15686 6010
rect 15698 5958 15750 6010
rect 15762 5958 15814 6010
rect 18606 5958 18658 6010
rect 18670 5958 18722 6010
rect 18734 5958 18786 6010
rect 18798 5958 18850 6010
rect 18862 5958 18914 6010
rect 4344 5856 4396 5908
rect 4436 5856 4488 5908
rect 5264 5856 5316 5908
rect 16488 5856 16540 5908
rect 3516 5788 3568 5840
rect 7656 5788 7708 5840
rect 8024 5831 8076 5840
rect 8024 5797 8033 5831
rect 8033 5797 8067 5831
rect 8067 5797 8076 5831
rect 8024 5788 8076 5797
rect 8484 5788 8536 5840
rect 12072 5788 12124 5840
rect 15200 5788 15252 5840
rect 572 5720 624 5772
rect 4252 5763 4304 5772
rect 4252 5729 4261 5763
rect 4261 5729 4295 5763
rect 4295 5729 4304 5763
rect 4252 5720 4304 5729
rect 5540 5720 5592 5772
rect 5908 5720 5960 5772
rect 7564 5720 7616 5772
rect 6552 5652 6604 5704
rect 10048 5695 10100 5704
rect 10048 5661 10057 5695
rect 10057 5661 10091 5695
rect 10091 5661 10100 5695
rect 10048 5652 10100 5661
rect 11336 5652 11388 5704
rect 13820 5763 13872 5772
rect 13820 5729 13830 5763
rect 13830 5729 13864 5763
rect 13864 5729 13872 5763
rect 13820 5720 13872 5729
rect 13176 5695 13228 5704
rect 13176 5661 13185 5695
rect 13185 5661 13219 5695
rect 13219 5661 13228 5695
rect 13176 5652 13228 5661
rect 13268 5695 13320 5704
rect 13268 5661 13277 5695
rect 13277 5661 13311 5695
rect 13311 5661 13320 5695
rect 13268 5652 13320 5661
rect 14924 5584 14976 5636
rect 1952 5516 2004 5568
rect 5080 5516 5132 5568
rect 6736 5516 6788 5568
rect 9220 5516 9272 5568
rect 11520 5516 11572 5568
rect 12072 5516 12124 5568
rect 12440 5559 12492 5568
rect 12440 5525 12449 5559
rect 12449 5525 12483 5559
rect 12483 5525 12492 5559
rect 12440 5516 12492 5525
rect 12716 5559 12768 5568
rect 12716 5525 12725 5559
rect 12725 5525 12759 5559
rect 12759 5525 12768 5559
rect 12716 5516 12768 5525
rect 15660 5720 15712 5772
rect 15844 5720 15896 5772
rect 16304 5720 16356 5772
rect 16948 5788 17000 5840
rect 16764 5720 16816 5772
rect 17408 5720 17460 5772
rect 15936 5584 15988 5636
rect 16304 5584 16356 5636
rect 17960 5652 18012 5704
rect 1556 5414 1608 5466
rect 1620 5414 1672 5466
rect 1684 5414 1736 5466
rect 1748 5414 1800 5466
rect 1812 5414 1864 5466
rect 4656 5414 4708 5466
rect 4720 5414 4772 5466
rect 4784 5414 4836 5466
rect 4848 5414 4900 5466
rect 4912 5414 4964 5466
rect 7756 5414 7808 5466
rect 7820 5414 7872 5466
rect 7884 5414 7936 5466
rect 7948 5414 8000 5466
rect 8012 5414 8064 5466
rect 10856 5414 10908 5466
rect 10920 5414 10972 5466
rect 10984 5414 11036 5466
rect 11048 5414 11100 5466
rect 11112 5414 11164 5466
rect 13956 5414 14008 5466
rect 14020 5414 14072 5466
rect 14084 5414 14136 5466
rect 14148 5414 14200 5466
rect 14212 5414 14264 5466
rect 17056 5414 17108 5466
rect 17120 5414 17172 5466
rect 17184 5414 17236 5466
rect 17248 5414 17300 5466
rect 17312 5414 17364 5466
rect 1952 5176 2004 5228
rect 2044 5151 2096 5160
rect 2044 5117 2053 5151
rect 2053 5117 2087 5151
rect 2087 5117 2096 5151
rect 2044 5108 2096 5117
rect 3056 5040 3108 5092
rect 5816 5312 5868 5364
rect 11336 5312 11388 5364
rect 15660 5312 15712 5364
rect 17592 5312 17644 5364
rect 12440 5244 12492 5296
rect 7656 5176 7708 5228
rect 8116 5176 8168 5228
rect 9128 5176 9180 5228
rect 12716 5176 12768 5228
rect 13268 5176 13320 5228
rect 10048 5108 10100 5160
rect 13544 5151 13596 5160
rect 13544 5117 13553 5151
rect 13553 5117 13587 5151
rect 13587 5117 13596 5151
rect 13544 5108 13596 5117
rect 16396 5176 16448 5228
rect 16028 5108 16080 5160
rect 17500 5108 17552 5160
rect 4528 5083 4580 5092
rect 4528 5049 4537 5083
rect 4537 5049 4571 5083
rect 4571 5049 4580 5083
rect 4528 5040 4580 5049
rect 5816 5040 5868 5092
rect 6644 5083 6696 5092
rect 3976 4972 4028 5024
rect 5172 4972 5224 5024
rect 6644 5049 6653 5083
rect 6653 5049 6687 5083
rect 6687 5049 6696 5083
rect 6644 5040 6696 5049
rect 8484 5040 8536 5092
rect 11520 5083 11572 5092
rect 11520 5049 11529 5083
rect 11529 5049 11563 5083
rect 11563 5049 11572 5083
rect 11520 5040 11572 5049
rect 13820 5083 13872 5092
rect 13820 5049 13829 5083
rect 13829 5049 13863 5083
rect 13863 5049 13872 5083
rect 13820 5040 13872 5049
rect 15844 5040 15896 5092
rect 16672 5040 16724 5092
rect 9956 4972 10008 5024
rect 11888 4972 11940 5024
rect 3106 4870 3158 4922
rect 3170 4870 3222 4922
rect 3234 4870 3286 4922
rect 3298 4870 3350 4922
rect 3362 4870 3414 4922
rect 6206 4870 6258 4922
rect 6270 4870 6322 4922
rect 6334 4870 6386 4922
rect 6398 4870 6450 4922
rect 6462 4870 6514 4922
rect 9306 4870 9358 4922
rect 9370 4870 9422 4922
rect 9434 4870 9486 4922
rect 9498 4870 9550 4922
rect 9562 4870 9614 4922
rect 12406 4870 12458 4922
rect 12470 4870 12522 4922
rect 12534 4870 12586 4922
rect 12598 4870 12650 4922
rect 12662 4870 12714 4922
rect 15506 4870 15558 4922
rect 15570 4870 15622 4922
rect 15634 4870 15686 4922
rect 15698 4870 15750 4922
rect 15762 4870 15814 4922
rect 18606 4870 18658 4922
rect 18670 4870 18722 4922
rect 18734 4870 18786 4922
rect 18798 4870 18850 4922
rect 18862 4870 18914 4922
rect 4528 4811 4580 4820
rect 4528 4777 4537 4811
rect 4537 4777 4571 4811
rect 4571 4777 4580 4811
rect 4528 4768 4580 4777
rect 6644 4768 6696 4820
rect 13820 4768 13872 4820
rect 16028 4811 16080 4820
rect 16028 4777 16037 4811
rect 16037 4777 16071 4811
rect 16071 4777 16080 4811
rect 16028 4768 16080 4777
rect 17500 4768 17552 4820
rect 2136 4700 2188 4752
rect 2964 4700 3016 4752
rect 572 4675 624 4684
rect 572 4641 581 4675
rect 581 4641 615 4675
rect 615 4641 624 4675
rect 572 4632 624 4641
rect 4252 4700 4304 4752
rect 12072 4700 12124 4752
rect 13268 4700 13320 4752
rect 13544 4700 13596 4752
rect 848 4607 900 4616
rect 848 4573 857 4607
rect 857 4573 891 4607
rect 891 4573 900 4607
rect 848 4564 900 4573
rect 2780 4564 2832 4616
rect 3516 4675 3568 4684
rect 3516 4641 3525 4675
rect 3525 4641 3559 4675
rect 3559 4641 3568 4675
rect 3516 4632 3568 4641
rect 5264 4632 5316 4684
rect 7288 4632 7340 4684
rect 9956 4675 10008 4684
rect 9956 4641 9965 4675
rect 9965 4641 9999 4675
rect 9999 4641 10008 4675
rect 9956 4632 10008 4641
rect 16396 4700 16448 4752
rect 14924 4675 14976 4684
rect 14924 4641 14933 4675
rect 14933 4641 14967 4675
rect 14967 4641 14976 4675
rect 14924 4632 14976 4641
rect 15384 4632 15436 4684
rect 4528 4607 4580 4616
rect 4528 4573 4537 4607
rect 4537 4573 4571 4607
rect 4571 4573 4580 4607
rect 4528 4564 4580 4573
rect 5080 4564 5132 4616
rect 6736 4564 6788 4616
rect 11244 4564 11296 4616
rect 13820 4607 13872 4616
rect 13820 4573 13829 4607
rect 13829 4573 13863 4607
rect 13863 4573 13872 4607
rect 13820 4564 13872 4573
rect 14740 4607 14792 4616
rect 14740 4573 14749 4607
rect 14749 4573 14783 4607
rect 14783 4573 14792 4607
rect 14740 4564 14792 4573
rect 3148 4471 3200 4480
rect 3148 4437 3157 4471
rect 3157 4437 3191 4471
rect 3191 4437 3200 4471
rect 3148 4428 3200 4437
rect 6828 4428 6880 4480
rect 11612 4428 11664 4480
rect 12256 4428 12308 4480
rect 1556 4326 1608 4378
rect 1620 4326 1672 4378
rect 1684 4326 1736 4378
rect 1748 4326 1800 4378
rect 1812 4326 1864 4378
rect 4656 4326 4708 4378
rect 4720 4326 4772 4378
rect 4784 4326 4836 4378
rect 4848 4326 4900 4378
rect 4912 4326 4964 4378
rect 7756 4326 7808 4378
rect 7820 4326 7872 4378
rect 7884 4326 7936 4378
rect 7948 4326 8000 4378
rect 8012 4326 8064 4378
rect 10856 4326 10908 4378
rect 10920 4326 10972 4378
rect 10984 4326 11036 4378
rect 11048 4326 11100 4378
rect 11112 4326 11164 4378
rect 13956 4326 14008 4378
rect 14020 4326 14072 4378
rect 14084 4326 14136 4378
rect 14148 4326 14200 4378
rect 14212 4326 14264 4378
rect 17056 4326 17108 4378
rect 17120 4326 17172 4378
rect 17184 4326 17236 4378
rect 17248 4326 17300 4378
rect 17312 4326 17364 4378
rect 848 4224 900 4276
rect 4528 4224 4580 4276
rect 11244 4224 11296 4276
rect 14740 4224 14792 4276
rect 5080 4156 5132 4208
rect 8208 4156 8260 4208
rect 3148 4088 3200 4140
rect 756 4063 808 4072
rect 756 4029 765 4063
rect 765 4029 799 4063
rect 799 4029 808 4063
rect 756 4020 808 4029
rect 3516 4020 3568 4072
rect 4712 4088 4764 4140
rect 5172 4088 5224 4140
rect 12808 4156 12860 4208
rect 16856 4156 16908 4208
rect 17592 4156 17644 4208
rect 14832 4088 14884 4140
rect 16488 4131 16540 4140
rect 16488 4097 16497 4131
rect 16497 4097 16531 4131
rect 16531 4097 16540 4131
rect 16488 4088 16540 4097
rect 16672 4088 16724 4140
rect 17408 4131 17460 4140
rect 17408 4097 17417 4131
rect 17417 4097 17451 4131
rect 17451 4097 17460 4131
rect 17408 4088 17460 4097
rect 4252 3952 4304 4004
rect 11244 4020 11296 4072
rect 11612 4020 11664 4072
rect 14372 4020 14424 4072
rect 8208 3952 8260 4004
rect 9036 3952 9088 4004
rect 12808 3952 12860 4004
rect 14188 3952 14240 4004
rect 16212 4020 16264 4072
rect 17500 4063 17552 4072
rect 17500 4029 17509 4063
rect 17509 4029 17543 4063
rect 17543 4029 17552 4063
rect 17500 4020 17552 4029
rect 7472 3884 7524 3936
rect 8484 3884 8536 3936
rect 8760 3927 8812 3936
rect 8760 3893 8769 3927
rect 8769 3893 8803 3927
rect 8803 3893 8812 3927
rect 8760 3884 8812 3893
rect 9128 3927 9180 3936
rect 9128 3893 9137 3927
rect 9137 3893 9171 3927
rect 9171 3893 9180 3927
rect 9128 3884 9180 3893
rect 11612 3927 11664 3936
rect 11612 3893 11621 3927
rect 11621 3893 11655 3927
rect 11655 3893 11664 3927
rect 11612 3884 11664 3893
rect 12256 3884 12308 3936
rect 13820 3884 13872 3936
rect 16120 3884 16172 3936
rect 16672 3952 16724 4004
rect 16580 3884 16632 3936
rect 17408 3884 17460 3936
rect 3106 3782 3158 3834
rect 3170 3782 3222 3834
rect 3234 3782 3286 3834
rect 3298 3782 3350 3834
rect 3362 3782 3414 3834
rect 6206 3782 6258 3834
rect 6270 3782 6322 3834
rect 6334 3782 6386 3834
rect 6398 3782 6450 3834
rect 6462 3782 6514 3834
rect 9306 3782 9358 3834
rect 9370 3782 9422 3834
rect 9434 3782 9486 3834
rect 9498 3782 9550 3834
rect 9562 3782 9614 3834
rect 12406 3782 12458 3834
rect 12470 3782 12522 3834
rect 12534 3782 12586 3834
rect 12598 3782 12650 3834
rect 12662 3782 12714 3834
rect 15506 3782 15558 3834
rect 15570 3782 15622 3834
rect 15634 3782 15686 3834
rect 15698 3782 15750 3834
rect 15762 3782 15814 3834
rect 18606 3782 18658 3834
rect 18670 3782 18722 3834
rect 18734 3782 18786 3834
rect 18798 3782 18850 3834
rect 18862 3782 18914 3834
rect 2044 3680 2096 3732
rect 5264 3723 5316 3732
rect 5264 3689 5273 3723
rect 5273 3689 5307 3723
rect 5307 3689 5316 3723
rect 5264 3680 5316 3689
rect 6092 3723 6144 3732
rect 6092 3689 6101 3723
rect 6101 3689 6135 3723
rect 6135 3689 6144 3723
rect 6092 3680 6144 3689
rect 6552 3680 6604 3732
rect 8484 3723 8536 3732
rect 8484 3689 8493 3723
rect 8493 3689 8527 3723
rect 8527 3689 8536 3723
rect 8484 3680 8536 3689
rect 14188 3723 14240 3732
rect 14188 3689 14197 3723
rect 14197 3689 14231 3723
rect 14231 3689 14240 3723
rect 14188 3680 14240 3689
rect 14556 3680 14608 3732
rect 16304 3723 16356 3732
rect 16304 3689 16313 3723
rect 16313 3689 16347 3723
rect 16347 3689 16356 3723
rect 16304 3680 16356 3689
rect 1400 3544 1452 3596
rect 3516 3587 3568 3596
rect 3516 3553 3525 3587
rect 3525 3553 3559 3587
rect 3559 3553 3568 3587
rect 4252 3612 4304 3664
rect 6644 3612 6696 3664
rect 3516 3544 3568 3553
rect 3976 3587 4028 3596
rect 3976 3553 3985 3587
rect 3985 3553 4019 3587
rect 4019 3553 4028 3587
rect 3976 3544 4028 3553
rect 4988 3544 5040 3596
rect 6828 3587 6880 3596
rect 6828 3553 6837 3587
rect 6837 3553 6871 3587
rect 6871 3553 6880 3587
rect 6828 3544 6880 3553
rect 11244 3587 11296 3596
rect 11244 3553 11253 3587
rect 11253 3553 11287 3587
rect 11287 3553 11296 3587
rect 11244 3544 11296 3553
rect 11336 3544 11388 3596
rect 12256 3544 12308 3596
rect 14372 3612 14424 3664
rect 14464 3544 14516 3596
rect 15108 3544 15160 3596
rect 16120 3587 16172 3596
rect 16120 3553 16129 3587
rect 16129 3553 16163 3587
rect 16163 3553 16172 3587
rect 16120 3544 16172 3553
rect 16580 3680 16632 3732
rect 17500 3680 17552 3732
rect 18144 3680 18196 3732
rect 16488 3544 16540 3596
rect 17408 3544 17460 3596
rect 18420 3587 18472 3596
rect 18420 3553 18429 3587
rect 18429 3553 18463 3587
rect 18463 3553 18472 3587
rect 18420 3544 18472 3553
rect 19064 3544 19116 3596
rect 10784 3408 10836 3460
rect 16212 3408 16264 3460
rect 2136 3340 2188 3392
rect 3516 3340 3568 3392
rect 16948 3340 17000 3392
rect 1556 3238 1608 3290
rect 1620 3238 1672 3290
rect 1684 3238 1736 3290
rect 1748 3238 1800 3290
rect 1812 3238 1864 3290
rect 4656 3238 4708 3290
rect 4720 3238 4772 3290
rect 4784 3238 4836 3290
rect 4848 3238 4900 3290
rect 4912 3238 4964 3290
rect 7756 3238 7808 3290
rect 7820 3238 7872 3290
rect 7884 3238 7936 3290
rect 7948 3238 8000 3290
rect 8012 3238 8064 3290
rect 10856 3238 10908 3290
rect 10920 3238 10972 3290
rect 10984 3238 11036 3290
rect 11048 3238 11100 3290
rect 11112 3238 11164 3290
rect 13956 3238 14008 3290
rect 14020 3238 14072 3290
rect 14084 3238 14136 3290
rect 14148 3238 14200 3290
rect 14212 3238 14264 3290
rect 17056 3238 17108 3290
rect 17120 3238 17172 3290
rect 17184 3238 17236 3290
rect 17248 3238 17300 3290
rect 17312 3238 17364 3290
rect 756 3136 808 3188
rect 4988 3179 5040 3188
rect 4988 3145 4997 3179
rect 4997 3145 5031 3179
rect 5031 3145 5040 3179
rect 4988 3136 5040 3145
rect 6644 3179 6696 3188
rect 6644 3145 6653 3179
rect 6653 3145 6687 3179
rect 6687 3145 6696 3179
rect 6644 3136 6696 3145
rect 6828 3136 6880 3188
rect 9128 3136 9180 3188
rect 11520 3179 11572 3188
rect 11520 3145 11529 3179
rect 11529 3145 11563 3179
rect 11563 3145 11572 3179
rect 11520 3136 11572 3145
rect 11796 3136 11848 3188
rect 12808 3136 12860 3188
rect 14832 3179 14884 3188
rect 14832 3145 14841 3179
rect 14841 3145 14875 3179
rect 14875 3145 14884 3179
rect 14832 3136 14884 3145
rect 16948 3136 17000 3188
rect 18420 3179 18472 3188
rect 18420 3145 18429 3179
rect 18429 3145 18463 3179
rect 18463 3145 18472 3179
rect 18420 3136 18472 3145
rect 5908 3000 5960 3052
rect 6644 3000 6696 3052
rect 7564 3043 7616 3052
rect 7564 3009 7573 3043
rect 7573 3009 7607 3043
rect 7607 3009 7616 3043
rect 7564 3000 7616 3009
rect 756 2975 808 2984
rect 756 2941 765 2975
rect 765 2941 799 2975
rect 799 2941 808 2975
rect 756 2932 808 2941
rect 7288 2975 7340 2984
rect 7288 2941 7297 2975
rect 7297 2941 7331 2975
rect 7331 2941 7340 2975
rect 7288 2932 7340 2941
rect 9036 2932 9088 2984
rect 11244 3000 11296 3052
rect 11428 3000 11480 3052
rect 10784 2975 10836 2984
rect 10784 2941 10793 2975
rect 10793 2941 10827 2975
rect 10827 2941 10836 2975
rect 10784 2932 10836 2941
rect 11336 2975 11388 2984
rect 11336 2941 11345 2975
rect 11345 2941 11379 2975
rect 11379 2941 11388 2975
rect 11336 2932 11388 2941
rect 5540 2864 5592 2916
rect 12808 3000 12860 3052
rect 13176 3000 13228 3052
rect 16488 3000 16540 3052
rect 15108 2932 15160 2984
rect 17592 2907 17644 2916
rect 17592 2873 17601 2907
rect 17601 2873 17635 2907
rect 17635 2873 17644 2907
rect 17592 2864 17644 2873
rect 5356 2839 5408 2848
rect 5356 2805 5365 2839
rect 5365 2805 5399 2839
rect 5399 2805 5408 2839
rect 5356 2796 5408 2805
rect 9036 2796 9088 2848
rect 11520 2796 11572 2848
rect 13176 2796 13228 2848
rect 13728 2796 13780 2848
rect 15200 2839 15252 2848
rect 15200 2805 15209 2839
rect 15209 2805 15243 2839
rect 15243 2805 15252 2839
rect 15200 2796 15252 2805
rect 17500 2839 17552 2848
rect 17500 2805 17509 2839
rect 17509 2805 17543 2839
rect 17543 2805 17552 2839
rect 17500 2796 17552 2805
rect 3106 2694 3158 2746
rect 3170 2694 3222 2746
rect 3234 2694 3286 2746
rect 3298 2694 3350 2746
rect 3362 2694 3414 2746
rect 6206 2694 6258 2746
rect 6270 2694 6322 2746
rect 6334 2694 6386 2746
rect 6398 2694 6450 2746
rect 6462 2694 6514 2746
rect 9306 2694 9358 2746
rect 9370 2694 9422 2746
rect 9434 2694 9486 2746
rect 9498 2694 9550 2746
rect 9562 2694 9614 2746
rect 12406 2694 12458 2746
rect 12470 2694 12522 2746
rect 12534 2694 12586 2746
rect 12598 2694 12650 2746
rect 12662 2694 12714 2746
rect 15506 2694 15558 2746
rect 15570 2694 15622 2746
rect 15634 2694 15686 2746
rect 15698 2694 15750 2746
rect 15762 2694 15814 2746
rect 18606 2694 18658 2746
rect 18670 2694 18722 2746
rect 18734 2694 18786 2746
rect 18798 2694 18850 2746
rect 18862 2694 18914 2746
rect 756 2592 808 2644
rect 1400 2592 1452 2644
rect 2228 2592 2280 2644
rect 5356 2635 5408 2644
rect 5356 2601 5365 2635
rect 5365 2601 5399 2635
rect 5399 2601 5408 2635
rect 5356 2592 5408 2601
rect 5540 2592 5592 2644
rect 8208 2635 8260 2644
rect 8208 2601 8217 2635
rect 8217 2601 8251 2635
rect 8251 2601 8260 2635
rect 8208 2592 8260 2601
rect 4160 2524 4212 2576
rect 8484 2524 8536 2576
rect 14372 2592 14424 2644
rect 15200 2635 15252 2644
rect 15200 2601 15209 2635
rect 15209 2601 15243 2635
rect 15243 2601 15252 2635
rect 15200 2592 15252 2601
rect 15384 2592 15436 2644
rect 17500 2592 17552 2644
rect 17592 2592 17644 2644
rect 940 2499 992 2508
rect 940 2465 949 2499
rect 949 2465 983 2499
rect 983 2465 992 2499
rect 940 2456 992 2465
rect 2872 2456 2924 2508
rect 5632 2456 5684 2508
rect 8576 2499 8628 2508
rect 8576 2465 8585 2499
rect 8585 2465 8619 2499
rect 8619 2465 8628 2499
rect 8576 2456 8628 2465
rect 13728 2499 13780 2508
rect 1032 2431 1084 2440
rect 1032 2397 1041 2431
rect 1041 2397 1075 2431
rect 1075 2397 1084 2431
rect 1032 2388 1084 2397
rect 2136 2431 2188 2440
rect 2136 2397 2145 2431
rect 2145 2397 2179 2431
rect 2179 2397 2188 2431
rect 2136 2388 2188 2397
rect 4068 2388 4120 2440
rect 13728 2465 13737 2499
rect 13737 2465 13771 2499
rect 13771 2465 13780 2499
rect 13728 2456 13780 2465
rect 15108 2524 15160 2576
rect 14372 2456 14424 2508
rect 17592 2499 17644 2508
rect 17592 2465 17601 2499
rect 17601 2465 17635 2499
rect 17635 2465 17644 2499
rect 17592 2456 17644 2465
rect 7564 2320 7616 2372
rect 13268 2363 13320 2372
rect 13268 2329 13277 2363
rect 13277 2329 13311 2363
rect 13311 2329 13320 2363
rect 13268 2320 13320 2329
rect 14464 2388 14516 2440
rect 15568 2388 15620 2440
rect 16304 2388 16356 2440
rect 14372 2320 14424 2372
rect 13728 2295 13780 2304
rect 13728 2261 13737 2295
rect 13737 2261 13771 2295
rect 13771 2261 13780 2295
rect 13728 2252 13780 2261
rect 1556 2150 1608 2202
rect 1620 2150 1672 2202
rect 1684 2150 1736 2202
rect 1748 2150 1800 2202
rect 1812 2150 1864 2202
rect 4656 2150 4708 2202
rect 4720 2150 4772 2202
rect 4784 2150 4836 2202
rect 4848 2150 4900 2202
rect 4912 2150 4964 2202
rect 7756 2150 7808 2202
rect 7820 2150 7872 2202
rect 7884 2150 7936 2202
rect 7948 2150 8000 2202
rect 8012 2150 8064 2202
rect 10856 2150 10908 2202
rect 10920 2150 10972 2202
rect 10984 2150 11036 2202
rect 11048 2150 11100 2202
rect 11112 2150 11164 2202
rect 13956 2150 14008 2202
rect 14020 2150 14072 2202
rect 14084 2150 14136 2202
rect 14148 2150 14200 2202
rect 14212 2150 14264 2202
rect 17056 2150 17108 2202
rect 17120 2150 17172 2202
rect 17184 2150 17236 2202
rect 17248 2150 17300 2202
rect 17312 2150 17364 2202
rect 1032 2048 1084 2100
rect 2872 2091 2924 2100
rect 2872 2057 2881 2091
rect 2881 2057 2915 2091
rect 2915 2057 2924 2091
rect 2872 2048 2924 2057
rect 4160 2048 4212 2100
rect 11612 2048 11664 2100
rect 2872 1912 2924 1964
rect 4068 1912 4120 1964
rect 7288 1980 7340 2032
rect 11888 2023 11940 2032
rect 11888 1989 11897 2023
rect 11897 1989 11931 2023
rect 11931 1989 11940 2023
rect 11888 1980 11940 1989
rect 8392 1912 8444 1964
rect 12532 1912 12584 1964
rect 13728 1980 13780 2032
rect 12716 1955 12768 1964
rect 12716 1921 12725 1955
rect 12725 1921 12759 1955
rect 12759 1921 12768 1955
rect 12716 1912 12768 1921
rect 13268 1912 13320 1964
rect 14004 1955 14056 1964
rect 14004 1921 14013 1955
rect 14013 1921 14047 1955
rect 14047 1921 14056 1955
rect 14004 1912 14056 1921
rect 14464 1912 14516 1964
rect 3976 1844 4028 1896
rect 4528 1844 4580 1896
rect 5172 1887 5224 1896
rect 5172 1853 5181 1887
rect 5181 1853 5215 1887
rect 5215 1853 5224 1887
rect 5172 1844 5224 1853
rect 8668 1844 8720 1896
rect 9128 1776 9180 1828
rect 13728 1844 13780 1896
rect 16212 2048 16264 2100
rect 16672 2091 16724 2100
rect 16672 2057 16681 2091
rect 16681 2057 16715 2091
rect 16715 2057 16724 2091
rect 16672 2048 16724 2057
rect 17960 1980 18012 2032
rect 15108 1844 15160 1896
rect 15384 1887 15436 1896
rect 15384 1853 15393 1887
rect 15393 1853 15427 1887
rect 15427 1853 15436 1887
rect 15384 1844 15436 1853
rect 15568 1887 15620 1896
rect 15568 1853 15577 1887
rect 15577 1853 15611 1887
rect 15611 1853 15620 1887
rect 16304 1912 16356 1964
rect 15568 1844 15620 1853
rect 16856 1844 16908 1896
rect 2964 1708 3016 1760
rect 4068 1708 4120 1760
rect 7564 1751 7616 1760
rect 7564 1717 7573 1751
rect 7573 1717 7607 1751
rect 7607 1717 7616 1751
rect 7564 1708 7616 1717
rect 11520 1751 11572 1760
rect 11520 1717 11529 1751
rect 11529 1717 11563 1751
rect 11563 1717 11572 1751
rect 11520 1708 11572 1717
rect 12808 1708 12860 1760
rect 16212 1751 16264 1760
rect 16212 1717 16221 1751
rect 16221 1717 16255 1751
rect 16255 1717 16264 1751
rect 16212 1708 16264 1717
rect 16304 1751 16356 1760
rect 16304 1717 16313 1751
rect 16313 1717 16347 1751
rect 16347 1717 16356 1751
rect 18420 1751 18472 1760
rect 16304 1708 16356 1717
rect 18420 1717 18429 1751
rect 18429 1717 18463 1751
rect 18463 1717 18472 1751
rect 18420 1708 18472 1717
rect 3106 1606 3158 1658
rect 3170 1606 3222 1658
rect 3234 1606 3286 1658
rect 3298 1606 3350 1658
rect 3362 1606 3414 1658
rect 6206 1606 6258 1658
rect 6270 1606 6322 1658
rect 6334 1606 6386 1658
rect 6398 1606 6450 1658
rect 6462 1606 6514 1658
rect 9306 1606 9358 1658
rect 9370 1606 9422 1658
rect 9434 1606 9486 1658
rect 9498 1606 9550 1658
rect 9562 1606 9614 1658
rect 12406 1606 12458 1658
rect 12470 1606 12522 1658
rect 12534 1606 12586 1658
rect 12598 1606 12650 1658
rect 12662 1606 12714 1658
rect 15506 1606 15558 1658
rect 15570 1606 15622 1658
rect 15634 1606 15686 1658
rect 15698 1606 15750 1658
rect 15762 1606 15814 1658
rect 18606 1606 18658 1658
rect 18670 1606 18722 1658
rect 18734 1606 18786 1658
rect 18798 1606 18850 1658
rect 18862 1606 18914 1658
rect 5632 1547 5684 1556
rect 940 1436 992 1488
rect 2688 1368 2740 1420
rect 2872 1436 2924 1488
rect 5632 1513 5641 1547
rect 5641 1513 5675 1547
rect 5675 1513 5684 1547
rect 5632 1504 5684 1513
rect 9128 1504 9180 1556
rect 9588 1504 9640 1556
rect 3976 1368 4028 1420
rect 5264 1411 5316 1420
rect 5264 1377 5273 1411
rect 5273 1377 5307 1411
rect 5307 1377 5316 1411
rect 5264 1368 5316 1377
rect 6552 1436 6604 1488
rect 7288 1436 7340 1488
rect 11520 1504 11572 1556
rect 13176 1547 13228 1556
rect 13176 1513 13185 1547
rect 13185 1513 13219 1547
rect 13219 1513 13228 1547
rect 13176 1504 13228 1513
rect 8116 1368 8168 1420
rect 8760 1368 8812 1420
rect 8944 1368 8996 1420
rect 4068 1300 4120 1352
rect 4620 1300 4672 1352
rect 5448 1300 5500 1352
rect 11428 1368 11480 1420
rect 11796 1411 11848 1420
rect 11796 1377 11805 1411
rect 11805 1377 11839 1411
rect 11839 1377 11848 1411
rect 11796 1368 11848 1377
rect 14372 1504 14424 1556
rect 16304 1504 16356 1556
rect 17592 1504 17644 1556
rect 15384 1436 15436 1488
rect 14004 1368 14056 1420
rect 15108 1411 15160 1420
rect 15108 1377 15117 1411
rect 15117 1377 15151 1411
rect 15151 1377 15160 1411
rect 15108 1368 15160 1377
rect 15844 1411 15896 1420
rect 15844 1377 15853 1411
rect 15853 1377 15887 1411
rect 15887 1377 15896 1411
rect 15844 1368 15896 1377
rect 17500 1368 17552 1420
rect 2872 1232 2924 1284
rect 5172 1232 5224 1284
rect 8576 1232 8628 1284
rect 8668 1232 8720 1284
rect 13728 1300 13780 1352
rect 16856 1300 16908 1352
rect 17408 1300 17460 1352
rect 17960 1300 18012 1352
rect 9036 1207 9088 1216
rect 9036 1173 9045 1207
rect 9045 1173 9079 1207
rect 9079 1173 9088 1207
rect 9036 1164 9088 1173
rect 12808 1232 12860 1284
rect 17592 1232 17644 1284
rect 1556 1062 1608 1114
rect 1620 1062 1672 1114
rect 1684 1062 1736 1114
rect 1748 1062 1800 1114
rect 1812 1062 1864 1114
rect 4656 1062 4708 1114
rect 4720 1062 4772 1114
rect 4784 1062 4836 1114
rect 4848 1062 4900 1114
rect 4912 1062 4964 1114
rect 7756 1062 7808 1114
rect 7820 1062 7872 1114
rect 7884 1062 7936 1114
rect 7948 1062 8000 1114
rect 8012 1062 8064 1114
rect 10856 1062 10908 1114
rect 10920 1062 10972 1114
rect 10984 1062 11036 1114
rect 11048 1062 11100 1114
rect 11112 1062 11164 1114
rect 13956 1062 14008 1114
rect 14020 1062 14072 1114
rect 14084 1062 14136 1114
rect 14148 1062 14200 1114
rect 14212 1062 14264 1114
rect 17056 1062 17108 1114
rect 17120 1062 17172 1114
rect 17184 1062 17236 1114
rect 17248 1062 17300 1114
rect 17312 1062 17364 1114
rect 2964 960 3016 1012
rect 5264 1003 5316 1012
rect 5264 969 5273 1003
rect 5273 969 5307 1003
rect 5307 969 5316 1003
rect 5264 960 5316 969
rect 8944 1003 8996 1012
rect 8944 969 8953 1003
rect 8953 969 8987 1003
rect 8987 969 8996 1003
rect 8944 960 8996 969
rect 17500 1003 17552 1012
rect 17500 969 17509 1003
rect 17509 969 17543 1003
rect 17543 969 17552 1003
rect 17500 960 17552 969
rect 17592 1003 17644 1012
rect 17592 969 17601 1003
rect 17601 969 17635 1003
rect 17635 969 17644 1003
rect 17592 960 17644 969
rect 5172 892 5224 944
rect 8668 892 8720 944
rect 9128 892 9180 944
rect 15844 892 15896 944
rect 2780 824 2832 876
rect 17408 867 17460 876
rect 17408 833 17417 867
rect 17417 833 17451 867
rect 17451 833 17460 867
rect 17408 824 17460 833
rect 3976 756 4028 808
rect 5448 799 5500 808
rect 5448 765 5457 799
rect 5457 765 5491 799
rect 5491 765 5500 799
rect 5448 756 5500 765
rect 8760 756 8812 808
rect 9588 756 9640 808
rect 17960 756 18012 808
rect 3106 518 3158 570
rect 3170 518 3222 570
rect 3234 518 3286 570
rect 3298 518 3350 570
rect 3362 518 3414 570
rect 6206 518 6258 570
rect 6270 518 6322 570
rect 6334 518 6386 570
rect 6398 518 6450 570
rect 6462 518 6514 570
rect 9306 518 9358 570
rect 9370 518 9422 570
rect 9434 518 9486 570
rect 9498 518 9550 570
rect 9562 518 9614 570
rect 12406 518 12458 570
rect 12470 518 12522 570
rect 12534 518 12586 570
rect 12598 518 12650 570
rect 12662 518 12714 570
rect 15506 518 15558 570
rect 15570 518 15622 570
rect 15634 518 15686 570
rect 15698 518 15750 570
rect 15762 518 15814 570
rect 18606 518 18658 570
rect 18670 518 18722 570
rect 18734 518 18786 570
rect 18798 518 18850 570
rect 18862 518 18914 570
<< metal2 >>
rect 1398 19200 1454 20000
rect 4250 19200 4306 20000
rect 7102 19200 7158 20000
rect 9954 19200 10010 20000
rect 12806 19200 12862 20000
rect 15396 19230 15608 19258
rect 1412 18426 1440 19200
rect 1556 18524 1864 18533
rect 1556 18522 1562 18524
rect 1618 18522 1642 18524
rect 1698 18522 1722 18524
rect 1778 18522 1802 18524
rect 1858 18522 1864 18524
rect 1618 18470 1620 18522
rect 1800 18470 1802 18522
rect 1556 18468 1562 18470
rect 1618 18468 1642 18470
rect 1698 18468 1722 18470
rect 1778 18468 1802 18470
rect 1858 18468 1864 18470
rect 1556 18459 1864 18468
rect 1400 18420 1452 18426
rect 1400 18362 1452 18368
rect 1400 18216 1452 18222
rect 1400 18158 1452 18164
rect 1952 18216 2004 18222
rect 1952 18158 2004 18164
rect 1216 18080 1268 18086
rect 1216 18022 1268 18028
rect 1228 17814 1256 18022
rect 1216 17808 1268 17814
rect 1216 17750 1268 17756
rect 572 17672 624 17678
rect 572 17614 624 17620
rect 584 16522 612 17614
rect 1412 17218 1440 18158
rect 1556 17436 1864 17445
rect 1556 17434 1562 17436
rect 1618 17434 1642 17436
rect 1698 17434 1722 17436
rect 1778 17434 1802 17436
rect 1858 17434 1864 17436
rect 1618 17382 1620 17434
rect 1800 17382 1802 17434
rect 1556 17380 1562 17382
rect 1618 17380 1642 17382
rect 1698 17380 1722 17382
rect 1778 17380 1802 17382
rect 1858 17380 1864 17382
rect 1556 17371 1864 17380
rect 1964 17338 1992 18158
rect 2964 18080 3016 18086
rect 2964 18022 3016 18028
rect 4068 18080 4120 18086
rect 4068 18022 4120 18028
rect 2504 17808 2556 17814
rect 2504 17750 2556 17756
rect 2412 17536 2464 17542
rect 2412 17478 2464 17484
rect 1952 17332 2004 17338
rect 1952 17274 2004 17280
rect 1412 17190 1716 17218
rect 1584 17128 1636 17134
rect 1584 17070 1636 17076
rect 1596 16726 1624 17070
rect 1688 16794 1716 17190
rect 1768 17128 1820 17134
rect 1768 17070 1820 17076
rect 1860 17128 1912 17134
rect 1860 17070 1912 17076
rect 2228 17128 2280 17134
rect 2228 17070 2280 17076
rect 2320 17128 2372 17134
rect 2320 17070 2372 17076
rect 1676 16788 1728 16794
rect 1676 16730 1728 16736
rect 1584 16720 1636 16726
rect 1584 16662 1636 16668
rect 1780 16590 1808 17070
rect 1872 16658 1900 17070
rect 1860 16652 1912 16658
rect 1860 16594 1912 16600
rect 1768 16584 1820 16590
rect 1768 16526 1820 16532
rect 1872 16538 1900 16594
rect 2240 16590 2268 17070
rect 2228 16584 2280 16590
rect 572 16516 624 16522
rect 572 16458 624 16464
rect 584 15570 612 16458
rect 1780 16454 1808 16526
rect 1872 16510 1992 16538
rect 2228 16526 2280 16532
rect 1768 16448 1820 16454
rect 1768 16390 1820 16396
rect 1556 16348 1864 16357
rect 1556 16346 1562 16348
rect 1618 16346 1642 16348
rect 1698 16346 1722 16348
rect 1778 16346 1802 16348
rect 1858 16346 1864 16348
rect 1618 16294 1620 16346
rect 1800 16294 1802 16346
rect 1556 16292 1562 16294
rect 1618 16292 1642 16294
rect 1698 16292 1722 16294
rect 1778 16292 1802 16294
rect 1858 16292 1864 16294
rect 1556 16283 1864 16292
rect 1964 16114 1992 16510
rect 2044 16448 2096 16454
rect 2044 16390 2096 16396
rect 1952 16108 2004 16114
rect 1952 16050 2004 16056
rect 848 15904 900 15910
rect 848 15846 900 15852
rect 860 15638 888 15846
rect 848 15632 900 15638
rect 848 15574 900 15580
rect 572 15564 624 15570
rect 572 15506 624 15512
rect 584 14482 612 15506
rect 1964 15434 1992 16050
rect 1952 15428 2004 15434
rect 1952 15370 2004 15376
rect 1556 15260 1864 15269
rect 1556 15258 1562 15260
rect 1618 15258 1642 15260
rect 1698 15258 1722 15260
rect 1778 15258 1802 15260
rect 1858 15258 1864 15260
rect 1618 15206 1620 15258
rect 1800 15206 1802 15258
rect 1556 15204 1562 15206
rect 1618 15204 1642 15206
rect 1698 15204 1722 15206
rect 1778 15204 1802 15206
rect 1858 15204 1864 15206
rect 1556 15195 1864 15204
rect 2056 14958 2084 16390
rect 2240 16114 2268 16526
rect 2228 16108 2280 16114
rect 2228 16050 2280 16056
rect 2136 15632 2188 15638
rect 2136 15574 2188 15580
rect 2044 14952 2096 14958
rect 2044 14894 2096 14900
rect 940 14816 992 14822
rect 940 14758 992 14764
rect 1952 14816 2004 14822
rect 1952 14758 2004 14764
rect 952 14482 980 14758
rect 572 14476 624 14482
rect 572 14418 624 14424
rect 940 14476 992 14482
rect 940 14418 992 14424
rect 584 13326 612 14418
rect 1556 14172 1864 14181
rect 1556 14170 1562 14172
rect 1618 14170 1642 14172
rect 1698 14170 1722 14172
rect 1778 14170 1802 14172
rect 1858 14170 1864 14172
rect 1618 14118 1620 14170
rect 1800 14118 1802 14170
rect 1556 14116 1562 14118
rect 1618 14116 1642 14118
rect 1698 14116 1722 14118
rect 1778 14116 1802 14118
rect 1858 14116 1864 14118
rect 1556 14107 1864 14116
rect 1964 14074 1992 14758
rect 2148 14550 2176 15574
rect 2240 15026 2268 16050
rect 2228 15020 2280 15026
rect 2228 14962 2280 14968
rect 2136 14544 2188 14550
rect 2136 14486 2188 14492
rect 1952 14068 2004 14074
rect 1952 14010 2004 14016
rect 572 13320 624 13326
rect 572 13262 624 13268
rect 584 12306 612 13262
rect 1556 13084 1864 13093
rect 1556 13082 1562 13084
rect 1618 13082 1642 13084
rect 1698 13082 1722 13084
rect 1778 13082 1802 13084
rect 1858 13082 1864 13084
rect 1618 13030 1620 13082
rect 1800 13030 1802 13082
rect 1556 13028 1562 13030
rect 1618 13028 1642 13030
rect 1698 13028 1722 13030
rect 1778 13028 1802 13030
rect 1858 13028 1864 13030
rect 1556 13019 1864 13028
rect 2240 12424 2268 14962
rect 2148 12396 2268 12424
rect 572 12300 624 12306
rect 572 12242 624 12248
rect 1124 12300 1176 12306
rect 1124 12242 1176 12248
rect 1136 11286 1164 12242
rect 1556 11996 1864 12005
rect 1556 11994 1562 11996
rect 1618 11994 1642 11996
rect 1698 11994 1722 11996
rect 1778 11994 1802 11996
rect 1858 11994 1864 11996
rect 1618 11942 1620 11994
rect 1800 11942 1802 11994
rect 1556 11940 1562 11942
rect 1618 11940 1642 11942
rect 1698 11940 1722 11942
rect 1778 11940 1802 11942
rect 1858 11940 1864 11942
rect 1556 11931 1864 11940
rect 1124 11280 1176 11286
rect 1124 11222 1176 11228
rect 1136 10606 1164 11222
rect 2148 11218 2176 12396
rect 2228 12300 2280 12306
rect 2228 12242 2280 12248
rect 2240 11694 2268 12242
rect 2228 11688 2280 11694
rect 2228 11630 2280 11636
rect 2136 11212 2188 11218
rect 2136 11154 2188 11160
rect 2228 11008 2280 11014
rect 2228 10950 2280 10956
rect 2332 10962 2360 17070
rect 2424 16794 2452 17478
rect 2516 17202 2544 17750
rect 2504 17196 2556 17202
rect 2504 17138 2556 17144
rect 2516 17066 2544 17138
rect 2976 17134 3004 18022
rect 3106 17980 3414 17989
rect 3106 17978 3112 17980
rect 3168 17978 3192 17980
rect 3248 17978 3272 17980
rect 3328 17978 3352 17980
rect 3408 17978 3414 17980
rect 3168 17926 3170 17978
rect 3350 17926 3352 17978
rect 3106 17924 3112 17926
rect 3168 17924 3192 17926
rect 3248 17924 3272 17926
rect 3328 17924 3352 17926
rect 3408 17924 3414 17926
rect 3106 17915 3414 17924
rect 2964 17128 3016 17134
rect 2964 17070 3016 17076
rect 3516 17128 3568 17134
rect 3516 17070 3568 17076
rect 2504 17060 2556 17066
rect 2504 17002 2556 17008
rect 2412 16788 2464 16794
rect 2412 16730 2464 16736
rect 2516 15638 2544 17002
rect 3106 16892 3414 16901
rect 3106 16890 3112 16892
rect 3168 16890 3192 16892
rect 3248 16890 3272 16892
rect 3328 16890 3352 16892
rect 3408 16890 3414 16892
rect 3168 16838 3170 16890
rect 3350 16838 3352 16890
rect 3106 16836 3112 16838
rect 3168 16836 3192 16838
rect 3248 16836 3272 16838
rect 3328 16836 3352 16838
rect 3408 16836 3414 16838
rect 3106 16827 3414 16836
rect 3528 16658 3556 17070
rect 4080 16726 4108 18022
rect 4264 17814 4292 19200
rect 4656 18524 4964 18533
rect 4656 18522 4662 18524
rect 4718 18522 4742 18524
rect 4798 18522 4822 18524
rect 4878 18522 4902 18524
rect 4958 18522 4964 18524
rect 4718 18470 4720 18522
rect 4900 18470 4902 18522
rect 4656 18468 4662 18470
rect 4718 18468 4742 18470
rect 4798 18468 4822 18470
rect 4878 18468 4902 18470
rect 4958 18468 4964 18470
rect 4656 18459 4964 18468
rect 4436 18284 4488 18290
rect 4436 18226 4488 18232
rect 5724 18284 5776 18290
rect 5724 18226 5776 18232
rect 4344 18080 4396 18086
rect 4344 18022 4396 18028
rect 4252 17808 4304 17814
rect 4172 17768 4252 17796
rect 4172 17338 4200 17768
rect 4252 17750 4304 17756
rect 4252 17672 4304 17678
rect 4252 17614 4304 17620
rect 4160 17332 4212 17338
rect 4160 17274 4212 17280
rect 4068 16720 4120 16726
rect 4068 16662 4120 16668
rect 3516 16652 3568 16658
rect 3516 16594 3568 16600
rect 2780 16448 2832 16454
rect 2780 16390 2832 16396
rect 3424 16448 3476 16454
rect 3476 16408 3556 16436
rect 3424 16390 3476 16396
rect 2792 16114 2820 16390
rect 2780 16108 2832 16114
rect 2780 16050 2832 16056
rect 2964 15972 3016 15978
rect 2964 15914 3016 15920
rect 2504 15632 2556 15638
rect 2504 15574 2556 15580
rect 2412 14952 2464 14958
rect 2412 14894 2464 14900
rect 2424 14550 2452 14894
rect 2504 14816 2556 14822
rect 2504 14758 2556 14764
rect 2412 14544 2464 14550
rect 2412 14486 2464 14492
rect 2516 13938 2544 14758
rect 2976 14618 3004 15914
rect 3106 15804 3414 15813
rect 3106 15802 3112 15804
rect 3168 15802 3192 15804
rect 3248 15802 3272 15804
rect 3328 15802 3352 15804
rect 3408 15802 3414 15804
rect 3168 15750 3170 15802
rect 3350 15750 3352 15802
rect 3106 15748 3112 15750
rect 3168 15748 3192 15750
rect 3248 15748 3272 15750
rect 3328 15748 3352 15750
rect 3408 15748 3414 15750
rect 3106 15739 3414 15748
rect 3528 14958 3556 16408
rect 4264 16046 4292 17614
rect 4356 17202 4384 18022
rect 4344 17196 4396 17202
rect 4344 17138 4396 17144
rect 4356 16794 4384 17138
rect 4448 17066 4476 18226
rect 5448 18148 5500 18154
rect 5448 18090 5500 18096
rect 4528 18080 4580 18086
rect 4528 18022 4580 18028
rect 4540 17882 4568 18022
rect 4528 17876 4580 17882
rect 4528 17818 4580 17824
rect 4656 17436 4964 17445
rect 4656 17434 4662 17436
rect 4718 17434 4742 17436
rect 4798 17434 4822 17436
rect 4878 17434 4902 17436
rect 4958 17434 4964 17436
rect 4718 17382 4720 17434
rect 4900 17382 4902 17434
rect 4656 17380 4662 17382
rect 4718 17380 4742 17382
rect 4798 17380 4822 17382
rect 4878 17380 4902 17382
rect 4958 17380 4964 17382
rect 4656 17371 4964 17380
rect 4436 17060 4488 17066
rect 4436 17002 4488 17008
rect 4344 16788 4396 16794
rect 4344 16730 4396 16736
rect 4656 16348 4964 16357
rect 4656 16346 4662 16348
rect 4718 16346 4742 16348
rect 4798 16346 4822 16348
rect 4878 16346 4902 16348
rect 4958 16346 4964 16348
rect 4718 16294 4720 16346
rect 4900 16294 4902 16346
rect 4656 16292 4662 16294
rect 4718 16292 4742 16294
rect 4798 16292 4822 16294
rect 4878 16292 4902 16294
rect 4958 16292 4964 16294
rect 4656 16283 4964 16292
rect 5460 16250 5488 18090
rect 5540 18080 5592 18086
rect 5540 18022 5592 18028
rect 5552 17338 5580 18022
rect 5540 17332 5592 17338
rect 5540 17274 5592 17280
rect 5448 16244 5500 16250
rect 5448 16186 5500 16192
rect 4252 16040 4304 16046
rect 4252 15982 4304 15988
rect 3700 15904 3752 15910
rect 3700 15846 3752 15852
rect 3516 14952 3568 14958
rect 3516 14894 3568 14900
rect 3106 14716 3414 14725
rect 3106 14714 3112 14716
rect 3168 14714 3192 14716
rect 3248 14714 3272 14716
rect 3328 14714 3352 14716
rect 3408 14714 3414 14716
rect 3168 14662 3170 14714
rect 3350 14662 3352 14714
rect 3106 14660 3112 14662
rect 3168 14660 3192 14662
rect 3248 14660 3272 14662
rect 3328 14660 3352 14662
rect 3408 14660 3414 14662
rect 3106 14651 3414 14660
rect 3712 14618 3740 15846
rect 4160 15632 4212 15638
rect 4160 15574 4212 15580
rect 3792 15088 3844 15094
rect 3792 15030 3844 15036
rect 2964 14612 3016 14618
rect 2964 14554 3016 14560
rect 3700 14612 3752 14618
rect 3700 14554 3752 14560
rect 3700 14476 3752 14482
rect 3700 14418 3752 14424
rect 2504 13932 2556 13938
rect 2504 13874 2556 13880
rect 2596 13864 2648 13870
rect 2596 13806 2648 13812
rect 2608 12306 2636 13806
rect 3106 13628 3414 13637
rect 3106 13626 3112 13628
rect 3168 13626 3192 13628
rect 3248 13626 3272 13628
rect 3328 13626 3352 13628
rect 3408 13626 3414 13628
rect 3168 13574 3170 13626
rect 3350 13574 3352 13626
rect 3106 13572 3112 13574
rect 3168 13572 3192 13574
rect 3248 13572 3272 13574
rect 3328 13572 3352 13574
rect 3408 13572 3414 13574
rect 3106 13563 3414 13572
rect 3712 13394 3740 14418
rect 3804 14414 3832 15030
rect 4172 14890 4200 15574
rect 5736 15502 5764 18226
rect 7116 18222 7144 19200
rect 7756 18524 8064 18533
rect 7756 18522 7762 18524
rect 7818 18522 7842 18524
rect 7898 18522 7922 18524
rect 7978 18522 8002 18524
rect 8058 18522 8064 18524
rect 7818 18470 7820 18522
rect 8000 18470 8002 18522
rect 7756 18468 7762 18470
rect 7818 18468 7842 18470
rect 7898 18468 7922 18470
rect 7978 18468 8002 18470
rect 8058 18468 8064 18470
rect 7756 18459 8064 18468
rect 9968 18306 9996 19200
rect 10856 18524 11164 18533
rect 10856 18522 10862 18524
rect 10918 18522 10942 18524
rect 10998 18522 11022 18524
rect 11078 18522 11102 18524
rect 11158 18522 11164 18524
rect 10918 18470 10920 18522
rect 11100 18470 11102 18522
rect 10856 18468 10862 18470
rect 10918 18468 10942 18470
rect 10998 18468 11022 18470
rect 11078 18468 11102 18470
rect 11158 18468 11164 18470
rect 10856 18459 11164 18468
rect 11152 18352 11204 18358
rect 9680 18284 9732 18290
rect 9968 18278 10088 18306
rect 11152 18294 11204 18300
rect 9680 18226 9732 18232
rect 7104 18216 7156 18222
rect 7104 18158 7156 18164
rect 7288 18216 7340 18222
rect 7288 18158 7340 18164
rect 6552 18148 6604 18154
rect 6552 18090 6604 18096
rect 6206 17980 6514 17989
rect 6206 17978 6212 17980
rect 6268 17978 6292 17980
rect 6348 17978 6372 17980
rect 6428 17978 6452 17980
rect 6508 17978 6514 17980
rect 6268 17926 6270 17978
rect 6450 17926 6452 17978
rect 6206 17924 6212 17926
rect 6268 17924 6292 17926
rect 6348 17924 6372 17926
rect 6428 17924 6452 17926
rect 6508 17924 6514 17926
rect 6206 17915 6514 17924
rect 6564 17202 6592 18090
rect 7012 17536 7064 17542
rect 7012 17478 7064 17484
rect 6552 17196 6604 17202
rect 6552 17138 6604 17144
rect 6828 16992 6880 16998
rect 6828 16934 6880 16940
rect 6206 16892 6514 16901
rect 6206 16890 6212 16892
rect 6268 16890 6292 16892
rect 6348 16890 6372 16892
rect 6428 16890 6452 16892
rect 6508 16890 6514 16892
rect 6268 16838 6270 16890
rect 6450 16838 6452 16890
rect 6206 16836 6212 16838
rect 6268 16836 6292 16838
rect 6348 16836 6372 16838
rect 6428 16836 6452 16838
rect 6508 16836 6514 16838
rect 6206 16827 6514 16836
rect 6206 15804 6514 15813
rect 6206 15802 6212 15804
rect 6268 15802 6292 15804
rect 6348 15802 6372 15804
rect 6428 15802 6452 15804
rect 6508 15802 6514 15804
rect 6268 15750 6270 15802
rect 6450 15750 6452 15802
rect 6206 15748 6212 15750
rect 6268 15748 6292 15750
rect 6348 15748 6372 15750
rect 6428 15748 6452 15750
rect 6508 15748 6514 15750
rect 6206 15739 6514 15748
rect 5816 15632 5868 15638
rect 5816 15574 5868 15580
rect 5448 15496 5500 15502
rect 5448 15438 5500 15444
rect 5724 15496 5776 15502
rect 5724 15438 5776 15444
rect 4656 15260 4964 15269
rect 4656 15258 4662 15260
rect 4718 15258 4742 15260
rect 4798 15258 4822 15260
rect 4878 15258 4902 15260
rect 4958 15258 4964 15260
rect 4718 15206 4720 15258
rect 4900 15206 4902 15258
rect 4656 15204 4662 15206
rect 4718 15204 4742 15206
rect 4798 15204 4822 15206
rect 4878 15204 4902 15206
rect 4958 15204 4964 15206
rect 4656 15195 4964 15204
rect 5080 15156 5132 15162
rect 5080 15098 5132 15104
rect 5092 14958 5120 15098
rect 4436 14952 4488 14958
rect 4620 14952 4672 14958
rect 4488 14912 4620 14940
rect 4436 14894 4488 14900
rect 4620 14894 4672 14900
rect 5080 14952 5132 14958
rect 5080 14894 5132 14900
rect 4160 14884 4212 14890
rect 4160 14826 4212 14832
rect 3792 14408 3844 14414
rect 3792 14350 3844 14356
rect 3804 13938 3832 14350
rect 3792 13932 3844 13938
rect 3792 13874 3844 13880
rect 3700 13388 3752 13394
rect 3700 13330 3752 13336
rect 3106 12540 3414 12549
rect 3106 12538 3112 12540
rect 3168 12538 3192 12540
rect 3248 12538 3272 12540
rect 3328 12538 3352 12540
rect 3408 12538 3414 12540
rect 3168 12486 3170 12538
rect 3350 12486 3352 12538
rect 3106 12484 3112 12486
rect 3168 12484 3192 12486
rect 3248 12484 3272 12486
rect 3328 12484 3352 12486
rect 3408 12484 3414 12486
rect 3106 12475 3414 12484
rect 2596 12300 2648 12306
rect 2596 12242 2648 12248
rect 2964 12300 3016 12306
rect 2964 12242 3016 12248
rect 3516 12300 3568 12306
rect 3516 12242 3568 12248
rect 2412 12164 2464 12170
rect 2412 12106 2464 12112
rect 2424 11694 2452 12106
rect 2412 11688 2464 11694
rect 2412 11630 2464 11636
rect 2976 11354 3004 12242
rect 3528 11830 3556 12242
rect 3700 12096 3752 12102
rect 3700 12038 3752 12044
rect 3516 11824 3568 11830
rect 3516 11766 3568 11772
rect 3712 11626 3740 12038
rect 4172 11898 4200 14826
rect 4528 14476 4580 14482
rect 4528 14418 4580 14424
rect 4540 13462 4568 14418
rect 4656 14172 4964 14181
rect 4656 14170 4662 14172
rect 4718 14170 4742 14172
rect 4798 14170 4822 14172
rect 4878 14170 4902 14172
rect 4958 14170 4964 14172
rect 4718 14118 4720 14170
rect 4900 14118 4902 14170
rect 4656 14116 4662 14118
rect 4718 14116 4742 14118
rect 4798 14116 4822 14118
rect 4878 14116 4902 14118
rect 4958 14116 4964 14118
rect 4656 14107 4964 14116
rect 5092 13802 5120 14894
rect 5460 14482 5488 15438
rect 5828 14822 5856 15574
rect 6840 15570 6868 16934
rect 7024 16726 7052 17478
rect 7012 16720 7064 16726
rect 7012 16662 7064 16668
rect 7116 16250 7144 18158
rect 7300 17202 7328 18158
rect 8392 18148 8444 18154
rect 8392 18090 8444 18096
rect 7840 18080 7892 18086
rect 7840 18022 7892 18028
rect 7852 17814 7880 18022
rect 7840 17808 7892 17814
rect 7840 17750 7892 17756
rect 7756 17436 8064 17445
rect 7756 17434 7762 17436
rect 7818 17434 7842 17436
rect 7898 17434 7922 17436
rect 7978 17434 8002 17436
rect 8058 17434 8064 17436
rect 7818 17382 7820 17434
rect 8000 17382 8002 17434
rect 7756 17380 7762 17382
rect 7818 17380 7842 17382
rect 7898 17380 7922 17382
rect 7978 17380 8002 17382
rect 8058 17380 8064 17382
rect 7756 17371 8064 17380
rect 8404 17202 8432 18090
rect 8484 18080 8536 18086
rect 8484 18022 8536 18028
rect 7288 17196 7340 17202
rect 7288 17138 7340 17144
rect 8392 17196 8444 17202
rect 8392 17138 8444 17144
rect 7656 16584 7708 16590
rect 7656 16526 7708 16532
rect 7472 16448 7524 16454
rect 7472 16390 7524 16396
rect 7104 16244 7156 16250
rect 7104 16186 7156 16192
rect 6828 15564 6880 15570
rect 6828 15506 6880 15512
rect 6840 15450 6868 15506
rect 6748 15422 6868 15450
rect 7288 15496 7340 15502
rect 7288 15438 7340 15444
rect 5724 14816 5776 14822
rect 5724 14758 5776 14764
rect 5816 14816 5868 14822
rect 5816 14758 5868 14764
rect 5736 14482 5764 14758
rect 5448 14476 5500 14482
rect 5448 14418 5500 14424
rect 5724 14476 5776 14482
rect 5724 14418 5776 14424
rect 5828 14074 5856 14758
rect 6206 14716 6514 14725
rect 6206 14714 6212 14716
rect 6268 14714 6292 14716
rect 6348 14714 6372 14716
rect 6428 14714 6452 14716
rect 6508 14714 6514 14716
rect 6268 14662 6270 14714
rect 6450 14662 6452 14714
rect 6206 14660 6212 14662
rect 6268 14660 6292 14662
rect 6348 14660 6372 14662
rect 6428 14660 6452 14662
rect 6508 14660 6514 14662
rect 6206 14651 6514 14660
rect 6748 14550 6776 15422
rect 7012 15020 7064 15026
rect 7012 14962 7064 14968
rect 6736 14544 6788 14550
rect 6736 14486 6788 14492
rect 5816 14068 5868 14074
rect 5816 14010 5868 14016
rect 6644 14068 6696 14074
rect 6644 14010 6696 14016
rect 5080 13796 5132 13802
rect 5080 13738 5132 13744
rect 6206 13628 6514 13637
rect 6206 13626 6212 13628
rect 6268 13626 6292 13628
rect 6348 13626 6372 13628
rect 6428 13626 6452 13628
rect 6508 13626 6514 13628
rect 6268 13574 6270 13626
rect 6450 13574 6452 13626
rect 6206 13572 6212 13574
rect 6268 13572 6292 13574
rect 6348 13572 6372 13574
rect 6428 13572 6452 13574
rect 6508 13572 6514 13574
rect 6206 13563 6514 13572
rect 4528 13456 4580 13462
rect 4528 13398 4580 13404
rect 6092 13456 6144 13462
rect 6092 13398 6144 13404
rect 6552 13456 6604 13462
rect 6552 13398 6604 13404
rect 4344 12640 4396 12646
rect 4344 12582 4396 12588
rect 4160 11892 4212 11898
rect 4080 11852 4160 11880
rect 3700 11620 3752 11626
rect 3700 11562 3752 11568
rect 3106 11452 3414 11461
rect 3106 11450 3112 11452
rect 3168 11450 3192 11452
rect 3248 11450 3272 11452
rect 3328 11450 3352 11452
rect 3408 11450 3414 11452
rect 3168 11398 3170 11450
rect 3350 11398 3352 11450
rect 3106 11396 3112 11398
rect 3168 11396 3192 11398
rect 3248 11396 3272 11398
rect 3328 11396 3352 11398
rect 3408 11396 3414 11398
rect 3106 11387 3414 11396
rect 2964 11348 3016 11354
rect 2964 11290 3016 11296
rect 2780 11212 2832 11218
rect 2780 11154 2832 11160
rect 1556 10908 1864 10917
rect 1556 10906 1562 10908
rect 1618 10906 1642 10908
rect 1698 10906 1722 10908
rect 1778 10906 1802 10908
rect 1858 10906 1864 10908
rect 1618 10854 1620 10906
rect 1800 10854 1802 10906
rect 1556 10852 1562 10854
rect 1618 10852 1642 10854
rect 1698 10852 1722 10854
rect 1778 10852 1802 10854
rect 1858 10852 1864 10854
rect 1556 10843 1864 10852
rect 2240 10826 2268 10950
rect 2332 10934 2452 10962
rect 2240 10798 2360 10826
rect 1124 10600 1176 10606
rect 1124 10542 1176 10548
rect 1952 10600 2004 10606
rect 1952 10542 2004 10548
rect 1136 10198 1164 10542
rect 1964 10266 1992 10542
rect 2332 10538 2360 10798
rect 2320 10532 2372 10538
rect 2320 10474 2372 10480
rect 1952 10260 2004 10266
rect 1952 10202 2004 10208
rect 1124 10192 1176 10198
rect 1124 10134 1176 10140
rect 2228 10056 2280 10062
rect 2228 9998 2280 10004
rect 1556 9820 1864 9829
rect 1556 9818 1562 9820
rect 1618 9818 1642 9820
rect 1698 9818 1722 9820
rect 1778 9818 1802 9820
rect 1858 9818 1864 9820
rect 1618 9766 1620 9818
rect 1800 9766 1802 9818
rect 1556 9764 1562 9766
rect 1618 9764 1642 9766
rect 1698 9764 1722 9766
rect 1778 9764 1802 9766
rect 1858 9764 1864 9766
rect 1556 9755 1864 9764
rect 2136 9376 2188 9382
rect 2136 9318 2188 9324
rect 848 8832 900 8838
rect 848 8774 900 8780
rect 860 8022 888 8774
rect 1556 8732 1864 8741
rect 1556 8730 1562 8732
rect 1618 8730 1642 8732
rect 1698 8730 1722 8732
rect 1778 8730 1802 8732
rect 1858 8730 1864 8732
rect 1618 8678 1620 8730
rect 1800 8678 1802 8730
rect 1556 8676 1562 8678
rect 1618 8676 1642 8678
rect 1698 8676 1722 8678
rect 1778 8676 1802 8678
rect 1858 8676 1864 8678
rect 1556 8667 1864 8676
rect 2148 8022 2176 9318
rect 2240 8974 2268 9998
rect 2332 9382 2360 10474
rect 2424 9518 2452 10934
rect 2792 10470 2820 11154
rect 2964 11076 3016 11082
rect 2964 11018 3016 11024
rect 3516 11076 3568 11082
rect 3516 11018 3568 11024
rect 2780 10464 2832 10470
rect 2780 10406 2832 10412
rect 2792 9994 2820 10406
rect 2872 10124 2924 10130
rect 2872 10066 2924 10072
rect 2780 9988 2832 9994
rect 2780 9930 2832 9936
rect 2412 9512 2464 9518
rect 2412 9454 2464 9460
rect 2320 9376 2372 9382
rect 2320 9318 2372 9324
rect 2320 9036 2372 9042
rect 2320 8978 2372 8984
rect 2228 8968 2280 8974
rect 2228 8910 2280 8916
rect 2332 8362 2360 8978
rect 2412 8968 2464 8974
rect 2412 8910 2464 8916
rect 2320 8356 2372 8362
rect 2320 8298 2372 8304
rect 848 8016 900 8022
rect 848 7958 900 7964
rect 2136 8016 2188 8022
rect 2136 7958 2188 7964
rect 572 7948 624 7954
rect 572 7890 624 7896
rect 584 6866 612 7890
rect 1556 7644 1864 7653
rect 1556 7642 1562 7644
rect 1618 7642 1642 7644
rect 1698 7642 1722 7644
rect 1778 7642 1802 7644
rect 1858 7642 1864 7644
rect 1618 7590 1620 7642
rect 1800 7590 1802 7642
rect 1556 7588 1562 7590
rect 1618 7588 1642 7590
rect 1698 7588 1722 7590
rect 1778 7588 1802 7590
rect 1858 7588 1864 7590
rect 1556 7579 1864 7588
rect 848 7200 900 7206
rect 848 7142 900 7148
rect 572 6860 624 6866
rect 572 6802 624 6808
rect 584 5778 612 6802
rect 860 6798 888 7142
rect 2148 6934 2176 7958
rect 2332 7886 2360 8298
rect 2320 7880 2372 7886
rect 2320 7822 2372 7828
rect 2332 7274 2360 7822
rect 2424 7410 2452 8910
rect 2792 8498 2820 9930
rect 2884 9654 2912 10066
rect 2872 9648 2924 9654
rect 2872 9590 2924 9596
rect 2976 8634 3004 11018
rect 3106 10364 3414 10373
rect 3106 10362 3112 10364
rect 3168 10362 3192 10364
rect 3248 10362 3272 10364
rect 3328 10362 3352 10364
rect 3408 10362 3414 10364
rect 3168 10310 3170 10362
rect 3350 10310 3352 10362
rect 3106 10308 3112 10310
rect 3168 10308 3192 10310
rect 3248 10308 3272 10310
rect 3328 10308 3352 10310
rect 3408 10308 3414 10310
rect 3106 10299 3414 10308
rect 3528 9518 3556 11018
rect 4080 10606 4108 11852
rect 4160 11834 4212 11840
rect 4356 11694 4384 12582
rect 4540 11830 4568 13398
rect 5448 13388 5500 13394
rect 5448 13330 5500 13336
rect 5080 13252 5132 13258
rect 5080 13194 5132 13200
rect 4988 13184 5040 13190
rect 4988 13126 5040 13132
rect 4656 13084 4964 13093
rect 4656 13082 4662 13084
rect 4718 13082 4742 13084
rect 4798 13082 4822 13084
rect 4878 13082 4902 13084
rect 4958 13082 4964 13084
rect 4718 13030 4720 13082
rect 4900 13030 4902 13082
rect 4656 13028 4662 13030
rect 4718 13028 4742 13030
rect 4798 13028 4822 13030
rect 4878 13028 4902 13030
rect 4958 13028 4964 13030
rect 4656 13019 4964 13028
rect 5000 12986 5028 13126
rect 4988 12980 5040 12986
rect 4988 12922 5040 12928
rect 5092 12782 5120 13194
rect 5460 12918 5488 13330
rect 5724 13320 5776 13326
rect 5724 13262 5776 13268
rect 6000 13320 6052 13326
rect 6000 13262 6052 13268
rect 5632 13184 5684 13190
rect 5632 13126 5684 13132
rect 5448 12912 5500 12918
rect 5448 12854 5500 12860
rect 5080 12776 5132 12782
rect 5080 12718 5132 12724
rect 5172 12232 5224 12238
rect 5172 12174 5224 12180
rect 4656 11996 4964 12005
rect 4656 11994 4662 11996
rect 4718 11994 4742 11996
rect 4798 11994 4822 11996
rect 4878 11994 4902 11996
rect 4958 11994 4964 11996
rect 4718 11942 4720 11994
rect 4900 11942 4902 11994
rect 4656 11940 4662 11942
rect 4718 11940 4742 11942
rect 4798 11940 4822 11942
rect 4878 11940 4902 11942
rect 4958 11940 4964 11942
rect 4656 11931 4964 11940
rect 4528 11824 4580 11830
rect 4528 11766 4580 11772
rect 4344 11688 4396 11694
rect 4264 11648 4344 11676
rect 4160 10736 4212 10742
rect 4160 10678 4212 10684
rect 4068 10600 4120 10606
rect 4068 10542 4120 10548
rect 3516 9512 3568 9518
rect 3516 9454 3568 9460
rect 4172 9450 4200 10678
rect 4264 9586 4292 11648
rect 4344 11630 4396 11636
rect 4540 11218 4568 11766
rect 4988 11552 5040 11558
rect 4988 11494 5040 11500
rect 4528 11212 4580 11218
rect 4528 11154 4580 11160
rect 5000 11014 5028 11494
rect 4988 11008 5040 11014
rect 4988 10950 5040 10956
rect 4656 10908 4964 10917
rect 4656 10906 4662 10908
rect 4718 10906 4742 10908
rect 4798 10906 4822 10908
rect 4878 10906 4902 10908
rect 4958 10906 4964 10908
rect 4718 10854 4720 10906
rect 4900 10854 4902 10906
rect 4656 10852 4662 10854
rect 4718 10852 4742 10854
rect 4798 10852 4822 10854
rect 4878 10852 4902 10854
rect 4958 10852 4964 10854
rect 4656 10843 4964 10852
rect 4344 10804 4396 10810
rect 4344 10746 4396 10752
rect 4356 10538 4384 10746
rect 4620 10600 4672 10606
rect 4448 10560 4620 10588
rect 4344 10532 4396 10538
rect 4344 10474 4396 10480
rect 4252 9580 4304 9586
rect 4252 9522 4304 9528
rect 4160 9444 4212 9450
rect 4160 9386 4212 9392
rect 3106 9276 3414 9285
rect 3106 9274 3112 9276
rect 3168 9274 3192 9276
rect 3248 9274 3272 9276
rect 3328 9274 3352 9276
rect 3408 9274 3414 9276
rect 3168 9222 3170 9274
rect 3350 9222 3352 9274
rect 3106 9220 3112 9222
rect 3168 9220 3192 9222
rect 3248 9220 3272 9222
rect 3328 9220 3352 9222
rect 3408 9220 3414 9222
rect 3106 9211 3414 9220
rect 3976 9036 4028 9042
rect 3976 8978 4028 8984
rect 3988 8634 4016 8978
rect 4264 8974 4292 9522
rect 4356 9042 4384 10474
rect 4448 9178 4476 10560
rect 4620 10542 4672 10548
rect 5000 10538 5028 10950
rect 4988 10532 5040 10538
rect 4988 10474 5040 10480
rect 4528 10192 4580 10198
rect 4528 10134 4580 10140
rect 4436 9172 4488 9178
rect 4436 9114 4488 9120
rect 4344 9036 4396 9042
rect 4344 8978 4396 8984
rect 4252 8968 4304 8974
rect 4252 8910 4304 8916
rect 2964 8628 3016 8634
rect 2964 8570 3016 8576
rect 3976 8628 4028 8634
rect 3976 8570 4028 8576
rect 2780 8492 2832 8498
rect 2780 8434 2832 8440
rect 2412 7404 2464 7410
rect 2412 7346 2464 7352
rect 2320 7268 2372 7274
rect 2320 7210 2372 7216
rect 2136 6928 2188 6934
rect 2136 6870 2188 6876
rect 848 6792 900 6798
rect 848 6734 900 6740
rect 1556 6556 1864 6565
rect 1556 6554 1562 6556
rect 1618 6554 1642 6556
rect 1698 6554 1722 6556
rect 1778 6554 1802 6556
rect 1858 6554 1864 6556
rect 1618 6502 1620 6554
rect 1800 6502 1802 6554
rect 1556 6500 1562 6502
rect 1618 6500 1642 6502
rect 1698 6500 1722 6502
rect 1778 6500 1802 6502
rect 1858 6500 1864 6502
rect 1556 6491 1864 6500
rect 572 5772 624 5778
rect 572 5714 624 5720
rect 584 4690 612 5714
rect 1952 5568 2004 5574
rect 1952 5510 2004 5516
rect 1556 5468 1864 5477
rect 1556 5466 1562 5468
rect 1618 5466 1642 5468
rect 1698 5466 1722 5468
rect 1778 5466 1802 5468
rect 1858 5466 1864 5468
rect 1618 5414 1620 5466
rect 1800 5414 1802 5466
rect 1556 5412 1562 5414
rect 1618 5412 1642 5414
rect 1698 5412 1722 5414
rect 1778 5412 1802 5414
rect 1858 5412 1864 5414
rect 1556 5403 1864 5412
rect 1964 5234 1992 5510
rect 1952 5228 2004 5234
rect 1952 5170 2004 5176
rect 2044 5160 2096 5166
rect 2044 5102 2096 5108
rect 572 4684 624 4690
rect 572 4626 624 4632
rect 848 4616 900 4622
rect 848 4558 900 4564
rect 860 4282 888 4558
rect 1556 4380 1864 4389
rect 1556 4378 1562 4380
rect 1618 4378 1642 4380
rect 1698 4378 1722 4380
rect 1778 4378 1802 4380
rect 1858 4378 1864 4380
rect 1618 4326 1620 4378
rect 1800 4326 1802 4378
rect 1556 4324 1562 4326
rect 1618 4324 1642 4326
rect 1698 4324 1722 4326
rect 1778 4324 1802 4326
rect 1858 4324 1864 4326
rect 1556 4315 1864 4324
rect 848 4276 900 4282
rect 848 4218 900 4224
rect 756 4072 808 4078
rect 756 4014 808 4020
rect 768 3194 796 4014
rect 2056 3738 2084 5102
rect 2148 4758 2176 6870
rect 2228 6792 2280 6798
rect 2228 6734 2280 6740
rect 2240 6458 2268 6734
rect 2424 6730 2452 7346
rect 2976 7342 3004 8570
rect 3976 8492 4028 8498
rect 3976 8434 4028 8440
rect 3106 8188 3414 8197
rect 3106 8186 3112 8188
rect 3168 8186 3192 8188
rect 3248 8186 3272 8188
rect 3328 8186 3352 8188
rect 3408 8186 3414 8188
rect 3168 8134 3170 8186
rect 3350 8134 3352 8186
rect 3106 8132 3112 8134
rect 3168 8132 3192 8134
rect 3248 8132 3272 8134
rect 3328 8132 3352 8134
rect 3408 8132 3414 8134
rect 3106 8123 3414 8132
rect 3988 7342 4016 8434
rect 4436 8424 4488 8430
rect 4436 8366 4488 8372
rect 4344 8288 4396 8294
rect 4344 8230 4396 8236
rect 4068 7744 4120 7750
rect 4068 7686 4120 7692
rect 4080 7410 4108 7686
rect 4356 7546 4384 8230
rect 4344 7540 4396 7546
rect 4344 7482 4396 7488
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 2964 7336 3016 7342
rect 2964 7278 3016 7284
rect 3976 7336 4028 7342
rect 3976 7278 4028 7284
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2792 7002 2820 7142
rect 2780 6996 2832 7002
rect 2780 6938 2832 6944
rect 2976 6934 3004 7278
rect 3106 7100 3414 7109
rect 3106 7098 3112 7100
rect 3168 7098 3192 7100
rect 3248 7098 3272 7100
rect 3328 7098 3352 7100
rect 3408 7098 3414 7100
rect 3168 7046 3170 7098
rect 3350 7046 3352 7098
rect 3106 7044 3112 7046
rect 3168 7044 3192 7046
rect 3248 7044 3272 7046
rect 3328 7044 3352 7046
rect 3408 7044 3414 7046
rect 3106 7035 3414 7044
rect 2964 6928 3016 6934
rect 2964 6870 3016 6876
rect 3516 6792 3568 6798
rect 3516 6734 3568 6740
rect 2412 6724 2464 6730
rect 2412 6666 2464 6672
rect 2228 6452 2280 6458
rect 2228 6394 2280 6400
rect 2228 6248 2280 6254
rect 2228 6190 2280 6196
rect 2136 4752 2188 4758
rect 2136 4694 2188 4700
rect 2044 3732 2096 3738
rect 2044 3674 2096 3680
rect 1400 3596 1452 3602
rect 1400 3538 1452 3544
rect 756 3188 808 3194
rect 756 3130 808 3136
rect 756 2984 808 2990
rect 756 2926 808 2932
rect 768 2650 796 2926
rect 1412 2650 1440 3538
rect 2136 3392 2188 3398
rect 2136 3334 2188 3340
rect 1556 3292 1864 3301
rect 1556 3290 1562 3292
rect 1618 3290 1642 3292
rect 1698 3290 1722 3292
rect 1778 3290 1802 3292
rect 1858 3290 1864 3292
rect 1618 3238 1620 3290
rect 1800 3238 1802 3290
rect 1556 3236 1562 3238
rect 1618 3236 1642 3238
rect 1698 3236 1722 3238
rect 1778 3236 1802 3238
rect 1858 3236 1864 3238
rect 1556 3227 1864 3236
rect 756 2644 808 2650
rect 756 2586 808 2592
rect 1400 2644 1452 2650
rect 1400 2586 1452 2592
rect 940 2508 992 2514
rect 940 2450 992 2456
rect 952 1494 980 2450
rect 2148 2446 2176 3334
rect 2240 2650 2268 6190
rect 3106 6012 3414 6021
rect 3106 6010 3112 6012
rect 3168 6010 3192 6012
rect 3248 6010 3272 6012
rect 3328 6010 3352 6012
rect 3408 6010 3414 6012
rect 3168 5958 3170 6010
rect 3350 5958 3352 6010
rect 3106 5956 3112 5958
rect 3168 5956 3192 5958
rect 3248 5956 3272 5958
rect 3328 5956 3352 5958
rect 3408 5956 3414 5958
rect 3106 5947 3414 5956
rect 3528 5846 3556 6734
rect 3516 5840 3568 5846
rect 3516 5782 3568 5788
rect 3056 5092 3108 5098
rect 2976 5052 3056 5080
rect 2976 4758 3004 5052
rect 3056 5034 3108 5040
rect 3106 4924 3414 4933
rect 3106 4922 3112 4924
rect 3168 4922 3192 4924
rect 3248 4922 3272 4924
rect 3328 4922 3352 4924
rect 3408 4922 3414 4924
rect 3168 4870 3170 4922
rect 3350 4870 3352 4922
rect 3106 4868 3112 4870
rect 3168 4868 3192 4870
rect 3248 4868 3272 4870
rect 3328 4868 3352 4870
rect 3408 4868 3414 4870
rect 3106 4859 3414 4868
rect 2964 4752 3016 4758
rect 2964 4694 3016 4700
rect 3528 4690 3556 5782
rect 3976 5024 4028 5030
rect 3976 4966 4028 4972
rect 3516 4684 3568 4690
rect 3516 4626 3568 4632
rect 2780 4616 2832 4622
rect 2780 4558 2832 4564
rect 2228 2644 2280 2650
rect 2228 2586 2280 2592
rect 1032 2440 1084 2446
rect 1032 2382 1084 2388
rect 2136 2440 2188 2446
rect 2136 2382 2188 2388
rect 1044 2106 1072 2382
rect 1556 2204 1864 2213
rect 1556 2202 1562 2204
rect 1618 2202 1642 2204
rect 1698 2202 1722 2204
rect 1778 2202 1802 2204
rect 1858 2202 1864 2204
rect 1618 2150 1620 2202
rect 1800 2150 1802 2202
rect 1556 2148 1562 2150
rect 1618 2148 1642 2150
rect 1698 2148 1722 2150
rect 1778 2148 1802 2150
rect 1858 2148 1864 2150
rect 1556 2139 1864 2148
rect 1032 2100 1084 2106
rect 1032 2042 1084 2048
rect 940 1488 992 1494
rect 2792 1442 2820 4558
rect 3148 4480 3200 4486
rect 3148 4422 3200 4428
rect 3160 4146 3188 4422
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 3528 4078 3556 4626
rect 3516 4072 3568 4078
rect 3516 4014 3568 4020
rect 3106 3836 3414 3845
rect 3106 3834 3112 3836
rect 3168 3834 3192 3836
rect 3248 3834 3272 3836
rect 3328 3834 3352 3836
rect 3408 3834 3414 3836
rect 3168 3782 3170 3834
rect 3350 3782 3352 3834
rect 3106 3780 3112 3782
rect 3168 3780 3192 3782
rect 3248 3780 3272 3782
rect 3328 3780 3352 3782
rect 3408 3780 3414 3782
rect 3106 3771 3414 3780
rect 3528 3602 3556 4014
rect 3988 3602 4016 4966
rect 3516 3596 3568 3602
rect 3516 3538 3568 3544
rect 3976 3596 4028 3602
rect 3976 3538 4028 3544
rect 3528 3398 3556 3538
rect 3516 3392 3568 3398
rect 3516 3334 3568 3340
rect 3106 2748 3414 2757
rect 3106 2746 3112 2748
rect 3168 2746 3192 2748
rect 3248 2746 3272 2748
rect 3328 2746 3352 2748
rect 3408 2746 3414 2748
rect 3168 2694 3170 2746
rect 3350 2694 3352 2746
rect 3106 2692 3112 2694
rect 3168 2692 3192 2694
rect 3248 2692 3272 2694
rect 3328 2692 3352 2694
rect 3408 2692 3414 2694
rect 3106 2683 3414 2692
rect 2872 2508 2924 2514
rect 2872 2450 2924 2456
rect 2884 2106 2912 2450
rect 2872 2100 2924 2106
rect 2872 2042 2924 2048
rect 2872 1964 2924 1970
rect 2872 1906 2924 1912
rect 2884 1494 2912 1906
rect 3988 1902 4016 3538
rect 4080 2446 4108 7346
rect 4356 7002 4384 7482
rect 4448 7274 4476 8366
rect 4540 8022 4568 10134
rect 4656 9820 4964 9829
rect 4656 9818 4662 9820
rect 4718 9818 4742 9820
rect 4798 9818 4822 9820
rect 4878 9818 4902 9820
rect 4958 9818 4964 9820
rect 4718 9766 4720 9818
rect 4900 9766 4902 9818
rect 4656 9764 4662 9766
rect 4718 9764 4742 9766
rect 4798 9764 4822 9766
rect 4878 9764 4902 9766
rect 4958 9764 4964 9766
rect 4656 9755 4964 9764
rect 5000 9382 5028 10474
rect 5184 10198 5212 12174
rect 5540 11892 5592 11898
rect 5540 11834 5592 11840
rect 5264 11756 5316 11762
rect 5264 11698 5316 11704
rect 5276 10742 5304 11698
rect 5448 11552 5500 11558
rect 5448 11494 5500 11500
rect 5460 11286 5488 11494
rect 5448 11280 5500 11286
rect 5448 11222 5500 11228
rect 5264 10736 5316 10742
rect 5264 10678 5316 10684
rect 5172 10192 5224 10198
rect 5172 10134 5224 10140
rect 5276 9674 5304 10678
rect 5092 9646 5304 9674
rect 4988 9376 5040 9382
rect 4988 9318 5040 9324
rect 5000 8974 5028 9318
rect 5092 9194 5120 9646
rect 5264 9376 5316 9382
rect 5264 9318 5316 9324
rect 5092 9166 5212 9194
rect 5080 9036 5132 9042
rect 5080 8978 5132 8984
rect 4988 8968 5040 8974
rect 4988 8910 5040 8916
rect 4656 8732 4964 8741
rect 4656 8730 4662 8732
rect 4718 8730 4742 8732
rect 4798 8730 4822 8732
rect 4878 8730 4902 8732
rect 4958 8730 4964 8732
rect 4718 8678 4720 8730
rect 4900 8678 4902 8730
rect 4656 8676 4662 8678
rect 4718 8676 4742 8678
rect 4798 8676 4822 8678
rect 4878 8676 4902 8678
rect 4958 8676 4964 8678
rect 4656 8667 4964 8676
rect 4528 8016 4580 8022
rect 4528 7958 4580 7964
rect 4656 7644 4964 7653
rect 4656 7642 4662 7644
rect 4718 7642 4742 7644
rect 4798 7642 4822 7644
rect 4878 7642 4902 7644
rect 4958 7642 4964 7644
rect 4718 7590 4720 7642
rect 4900 7590 4902 7642
rect 4656 7588 4662 7590
rect 4718 7588 4742 7590
rect 4798 7588 4822 7590
rect 4878 7588 4902 7590
rect 4958 7588 4964 7590
rect 4656 7579 4964 7588
rect 4436 7268 4488 7274
rect 4436 7210 4488 7216
rect 4344 6996 4396 7002
rect 4344 6938 4396 6944
rect 4344 6792 4396 6798
rect 4344 6734 4396 6740
rect 4252 6316 4304 6322
rect 4252 6258 4304 6264
rect 4264 5778 4292 6258
rect 4356 5914 4384 6734
rect 4656 6556 4964 6565
rect 4656 6554 4662 6556
rect 4718 6554 4742 6556
rect 4798 6554 4822 6556
rect 4878 6554 4902 6556
rect 4958 6554 4964 6556
rect 4718 6502 4720 6554
rect 4900 6502 4902 6554
rect 4656 6500 4662 6502
rect 4718 6500 4742 6502
rect 4798 6500 4822 6502
rect 4878 6500 4902 6502
rect 4958 6500 4964 6502
rect 4656 6491 4964 6500
rect 5000 6254 5028 8910
rect 5092 6254 5120 8978
rect 5184 8838 5212 9166
rect 5276 9042 5304 9318
rect 5264 9036 5316 9042
rect 5264 8978 5316 8984
rect 5172 8832 5224 8838
rect 5172 8774 5224 8780
rect 5184 8634 5212 8774
rect 5172 8628 5224 8634
rect 5172 8570 5224 8576
rect 5184 6458 5212 8570
rect 5264 8424 5316 8430
rect 5264 8366 5316 8372
rect 5276 8090 5304 8366
rect 5264 8084 5316 8090
rect 5264 8026 5316 8032
rect 5552 7886 5580 11834
rect 5644 11694 5672 13126
rect 5736 11898 5764 13262
rect 6012 12782 6040 13262
rect 6000 12776 6052 12782
rect 6000 12718 6052 12724
rect 5724 11892 5776 11898
rect 5724 11834 5776 11840
rect 6012 11694 6040 12718
rect 5632 11688 5684 11694
rect 5632 11630 5684 11636
rect 6000 11688 6052 11694
rect 6000 11630 6052 11636
rect 6104 11558 6132 13398
rect 6206 12540 6514 12549
rect 6206 12538 6212 12540
rect 6268 12538 6292 12540
rect 6348 12538 6372 12540
rect 6428 12538 6452 12540
rect 6508 12538 6514 12540
rect 6268 12486 6270 12538
rect 6450 12486 6452 12538
rect 6206 12484 6212 12486
rect 6268 12484 6292 12486
rect 6348 12484 6372 12486
rect 6428 12484 6452 12486
rect 6508 12484 6514 12486
rect 6206 12475 6514 12484
rect 6564 11762 6592 13398
rect 6656 13394 6684 14010
rect 6748 13394 6776 14486
rect 7024 14278 7052 14962
rect 7300 14804 7328 15438
rect 7484 14958 7512 16390
rect 7564 15700 7616 15706
rect 7564 15642 7616 15648
rect 7576 15026 7604 15642
rect 7668 15502 7696 16526
rect 7756 16348 8064 16357
rect 7756 16346 7762 16348
rect 7818 16346 7842 16348
rect 7898 16346 7922 16348
rect 7978 16346 8002 16348
rect 8058 16346 8064 16348
rect 7818 16294 7820 16346
rect 8000 16294 8002 16346
rect 7756 16292 7762 16294
rect 7818 16292 7842 16294
rect 7898 16292 7922 16294
rect 7978 16292 8002 16294
rect 8058 16292 8064 16294
rect 7756 16283 8064 16292
rect 7656 15496 7708 15502
rect 7656 15438 7708 15444
rect 7564 15020 7616 15026
rect 7564 14962 7616 14968
rect 7472 14952 7524 14958
rect 7472 14894 7524 14900
rect 7668 14804 7696 15438
rect 7756 15260 8064 15269
rect 7756 15258 7762 15260
rect 7818 15258 7842 15260
rect 7898 15258 7922 15260
rect 7978 15258 8002 15260
rect 8058 15258 8064 15260
rect 7818 15206 7820 15258
rect 8000 15206 8002 15258
rect 7756 15204 7762 15206
rect 7818 15204 7842 15206
rect 7898 15204 7922 15206
rect 7978 15204 8002 15206
rect 8058 15204 8064 15206
rect 7756 15195 8064 15204
rect 7840 14816 7892 14822
rect 7300 14776 7604 14804
rect 7668 14776 7840 14804
rect 7012 14272 7064 14278
rect 7012 14214 7064 14220
rect 7380 14272 7432 14278
rect 7380 14214 7432 14220
rect 7472 14272 7524 14278
rect 7472 14214 7524 14220
rect 6828 13864 6880 13870
rect 7104 13864 7156 13870
rect 6880 13824 7052 13852
rect 6828 13806 6880 13812
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 6840 13462 6868 13670
rect 6828 13456 6880 13462
rect 6828 13398 6880 13404
rect 6644 13388 6696 13394
rect 6644 13330 6696 13336
rect 6736 13388 6788 13394
rect 6736 13330 6788 13336
rect 6644 12776 6696 12782
rect 6644 12718 6696 12724
rect 6552 11756 6604 11762
rect 6552 11698 6604 11704
rect 6552 11620 6604 11626
rect 6552 11562 6604 11568
rect 6092 11552 6144 11558
rect 6092 11494 6144 11500
rect 6206 11452 6514 11461
rect 6206 11450 6212 11452
rect 6268 11450 6292 11452
rect 6348 11450 6372 11452
rect 6428 11450 6452 11452
rect 6508 11450 6514 11452
rect 6268 11398 6270 11450
rect 6450 11398 6452 11450
rect 6206 11396 6212 11398
rect 6268 11396 6292 11398
rect 6348 11396 6372 11398
rect 6428 11396 6452 11398
rect 6508 11396 6514 11398
rect 6206 11387 6514 11396
rect 5632 11008 5684 11014
rect 5632 10950 5684 10956
rect 5644 9178 5672 10950
rect 6564 10810 6592 11562
rect 6552 10804 6604 10810
rect 6552 10746 6604 10752
rect 6206 10364 6514 10373
rect 6206 10362 6212 10364
rect 6268 10362 6292 10364
rect 6348 10362 6372 10364
rect 6428 10362 6452 10364
rect 6508 10362 6514 10364
rect 6268 10310 6270 10362
rect 6450 10310 6452 10362
rect 6206 10308 6212 10310
rect 6268 10308 6292 10310
rect 6348 10308 6372 10310
rect 6428 10308 6452 10310
rect 6508 10308 6514 10310
rect 6206 10299 6514 10308
rect 6656 10266 6684 12718
rect 6748 11286 6776 13330
rect 6920 13252 6972 13258
rect 6920 13194 6972 13200
rect 6932 12782 6960 13194
rect 7024 12986 7052 13824
rect 7104 13806 7156 13812
rect 7012 12980 7064 12986
rect 7012 12922 7064 12928
rect 6920 12776 6972 12782
rect 6920 12718 6972 12724
rect 7012 12776 7064 12782
rect 7012 12718 7064 12724
rect 6920 12640 6972 12646
rect 6920 12582 6972 12588
rect 6932 11354 6960 12582
rect 6920 11348 6972 11354
rect 6920 11290 6972 11296
rect 6736 11280 6788 11286
rect 6736 11222 6788 11228
rect 7024 10266 7052 12718
rect 7116 11898 7144 13806
rect 7196 13796 7248 13802
rect 7196 13738 7248 13744
rect 7208 12782 7236 13738
rect 7288 12844 7340 12850
rect 7288 12786 7340 12792
rect 7196 12776 7248 12782
rect 7196 12718 7248 12724
rect 7196 12300 7248 12306
rect 7196 12242 7248 12248
rect 7208 11898 7236 12242
rect 7104 11892 7156 11898
rect 7104 11834 7156 11840
rect 7196 11892 7248 11898
rect 7196 11834 7248 11840
rect 6644 10260 6696 10266
rect 6644 10202 6696 10208
rect 7012 10260 7064 10266
rect 7012 10202 7064 10208
rect 7012 10124 7064 10130
rect 7012 10066 7064 10072
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 6206 9276 6514 9285
rect 6206 9274 6212 9276
rect 6268 9274 6292 9276
rect 6348 9274 6372 9276
rect 6428 9274 6452 9276
rect 6508 9274 6514 9276
rect 6268 9222 6270 9274
rect 6450 9222 6452 9274
rect 6206 9220 6212 9222
rect 6268 9220 6292 9222
rect 6348 9220 6372 9222
rect 6428 9220 6452 9222
rect 6508 9220 6514 9222
rect 6206 9211 6514 9220
rect 5632 9172 5684 9178
rect 5632 9114 5684 9120
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 5644 8634 5672 8910
rect 6840 8838 6868 9998
rect 7024 9586 7052 10066
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 5908 8832 5960 8838
rect 5908 8774 5960 8780
rect 6828 8832 6880 8838
rect 6828 8774 6880 8780
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 5632 8424 5684 8430
rect 5632 8366 5684 8372
rect 5540 7880 5592 7886
rect 5540 7822 5592 7828
rect 5264 7812 5316 7818
rect 5264 7754 5316 7760
rect 5276 7274 5304 7754
rect 5264 7268 5316 7274
rect 5264 7210 5316 7216
rect 5448 7268 5500 7274
rect 5552 7256 5580 7822
rect 5644 7546 5672 8366
rect 5816 8356 5868 8362
rect 5816 8298 5868 8304
rect 5828 7886 5856 8298
rect 5816 7880 5868 7886
rect 5816 7822 5868 7828
rect 5632 7540 5684 7546
rect 5632 7482 5684 7488
rect 5828 7410 5856 7822
rect 5816 7404 5868 7410
rect 5816 7346 5868 7352
rect 5920 7342 5948 8774
rect 6840 8430 6868 8774
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6206 8188 6514 8197
rect 6206 8186 6212 8188
rect 6268 8186 6292 8188
rect 6348 8186 6372 8188
rect 6428 8186 6452 8188
rect 6508 8186 6514 8188
rect 6268 8134 6270 8186
rect 6450 8134 6452 8186
rect 6206 8132 6212 8134
rect 6268 8132 6292 8134
rect 6348 8132 6372 8134
rect 6428 8132 6452 8134
rect 6508 8132 6514 8134
rect 6206 8123 6514 8132
rect 7300 7342 7328 12786
rect 7392 11694 7420 14214
rect 7484 13870 7512 14214
rect 7472 13864 7524 13870
rect 7472 13806 7524 13812
rect 7576 12442 7604 14776
rect 7840 14758 7892 14764
rect 7852 14482 7880 14758
rect 8496 14550 8524 18022
rect 9306 17980 9614 17989
rect 9306 17978 9312 17980
rect 9368 17978 9392 17980
rect 9448 17978 9472 17980
rect 9528 17978 9552 17980
rect 9608 17978 9614 17980
rect 9368 17926 9370 17978
rect 9550 17926 9552 17978
rect 9306 17924 9312 17926
rect 9368 17924 9392 17926
rect 9448 17924 9472 17926
rect 9528 17924 9552 17926
rect 9608 17924 9614 17926
rect 9306 17915 9614 17924
rect 9306 16892 9614 16901
rect 9306 16890 9312 16892
rect 9368 16890 9392 16892
rect 9448 16890 9472 16892
rect 9528 16890 9552 16892
rect 9608 16890 9614 16892
rect 9368 16838 9370 16890
rect 9550 16838 9552 16890
rect 9306 16836 9312 16838
rect 9368 16836 9392 16838
rect 9448 16836 9472 16838
rect 9528 16836 9552 16838
rect 9608 16836 9614 16838
rect 9306 16827 9614 16836
rect 8760 15972 8812 15978
rect 8760 15914 8812 15920
rect 8668 15360 8720 15366
rect 8668 15302 8720 15308
rect 8484 14544 8536 14550
rect 8484 14486 8536 14492
rect 7840 14476 7892 14482
rect 7840 14418 7892 14424
rect 8208 14476 8260 14482
rect 8208 14418 8260 14424
rect 8116 14408 8168 14414
rect 8116 14350 8168 14356
rect 7756 14172 8064 14181
rect 7756 14170 7762 14172
rect 7818 14170 7842 14172
rect 7898 14170 7922 14172
rect 7978 14170 8002 14172
rect 8058 14170 8064 14172
rect 7818 14118 7820 14170
rect 8000 14118 8002 14170
rect 7756 14116 7762 14118
rect 7818 14116 7842 14118
rect 7898 14116 7922 14118
rect 7978 14116 8002 14118
rect 8058 14116 8064 14118
rect 7756 14107 8064 14116
rect 8128 13546 8156 14350
rect 8220 13938 8248 14418
rect 8208 13932 8260 13938
rect 8208 13874 8260 13880
rect 8496 13802 8524 14486
rect 8680 14074 8708 15302
rect 8772 15162 8800 15914
rect 9306 15804 9614 15813
rect 9306 15802 9312 15804
rect 9368 15802 9392 15804
rect 9448 15802 9472 15804
rect 9528 15802 9552 15804
rect 9608 15802 9614 15804
rect 9368 15750 9370 15802
rect 9550 15750 9552 15802
rect 9306 15748 9312 15750
rect 9368 15748 9392 15750
rect 9448 15748 9472 15750
rect 9528 15748 9552 15750
rect 9608 15748 9614 15750
rect 9306 15739 9614 15748
rect 9692 15706 9720 18226
rect 9956 18148 10008 18154
rect 9956 18090 10008 18096
rect 9968 17746 9996 18090
rect 9956 17740 10008 17746
rect 9956 17682 10008 17688
rect 10060 17338 10088 18278
rect 11164 18222 11192 18294
rect 11152 18216 11204 18222
rect 12440 18216 12492 18222
rect 11152 18158 11204 18164
rect 12268 18164 12440 18170
rect 12268 18158 12492 18164
rect 11336 18148 11388 18154
rect 11336 18090 11388 18096
rect 11428 18148 11480 18154
rect 11428 18090 11480 18096
rect 12268 18142 12480 18158
rect 10140 18080 10192 18086
rect 10140 18022 10192 18028
rect 11244 18080 11296 18086
rect 11244 18022 11296 18028
rect 10048 17332 10100 17338
rect 10048 17274 10100 17280
rect 10152 16590 10180 18022
rect 10324 17672 10376 17678
rect 10324 17614 10376 17620
rect 10336 17270 10364 17614
rect 10856 17436 11164 17445
rect 10856 17434 10862 17436
rect 10918 17434 10942 17436
rect 10998 17434 11022 17436
rect 11078 17434 11102 17436
rect 11158 17434 11164 17436
rect 10918 17382 10920 17434
rect 11100 17382 11102 17434
rect 10856 17380 10862 17382
rect 10918 17380 10942 17382
rect 10998 17380 11022 17382
rect 11078 17380 11102 17382
rect 11158 17380 11164 17382
rect 10856 17371 11164 17380
rect 10324 17264 10376 17270
rect 10324 17206 10376 17212
rect 11256 17134 11284 18022
rect 11244 17128 11296 17134
rect 11244 17070 11296 17076
rect 10232 16720 10284 16726
rect 10284 16680 10364 16708
rect 10232 16662 10284 16668
rect 10140 16584 10192 16590
rect 10140 16526 10192 16532
rect 10152 16046 10180 16526
rect 10140 16040 10192 16046
rect 10140 15982 10192 15988
rect 9680 15700 9732 15706
rect 9680 15642 9732 15648
rect 10152 15638 10180 15982
rect 10140 15632 10192 15638
rect 10140 15574 10192 15580
rect 10140 15360 10192 15366
rect 10140 15302 10192 15308
rect 8760 15156 8812 15162
rect 8760 15098 8812 15104
rect 9036 14884 9088 14890
rect 9036 14826 9088 14832
rect 8668 14068 8720 14074
rect 8668 14010 8720 14016
rect 8484 13796 8536 13802
rect 8484 13738 8536 13744
rect 8036 13530 8156 13546
rect 8024 13524 8156 13530
rect 8076 13518 8156 13524
rect 8024 13466 8076 13472
rect 7656 13184 7708 13190
rect 7656 13126 7708 13132
rect 7564 12436 7616 12442
rect 7564 12378 7616 12384
rect 7564 12096 7616 12102
rect 7564 12038 7616 12044
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 7576 10130 7604 12038
rect 7668 11762 7696 13126
rect 7756 13084 8064 13093
rect 7756 13082 7762 13084
rect 7818 13082 7842 13084
rect 7898 13082 7922 13084
rect 7978 13082 8002 13084
rect 8058 13082 8064 13084
rect 7818 13030 7820 13082
rect 8000 13030 8002 13082
rect 7756 13028 7762 13030
rect 7818 13028 7842 13030
rect 7898 13028 7922 13030
rect 7978 13028 8002 13030
rect 8058 13028 8064 13030
rect 7756 13019 8064 13028
rect 8680 12782 8708 14010
rect 8944 13796 8996 13802
rect 8944 13738 8996 13744
rect 8852 13320 8904 13326
rect 8852 13262 8904 13268
rect 8668 12776 8720 12782
rect 8668 12718 8720 12724
rect 8668 12640 8720 12646
rect 8668 12582 8720 12588
rect 8576 12368 8628 12374
rect 8496 12316 8576 12322
rect 8496 12310 8628 12316
rect 8496 12294 8616 12310
rect 7756 11996 8064 12005
rect 7756 11994 7762 11996
rect 7818 11994 7842 11996
rect 7898 11994 7922 11996
rect 7978 11994 8002 11996
rect 8058 11994 8064 11996
rect 7818 11942 7820 11994
rect 8000 11942 8002 11994
rect 7756 11940 7762 11942
rect 7818 11940 7842 11942
rect 7898 11940 7922 11942
rect 7978 11940 8002 11942
rect 8058 11940 8064 11942
rect 7756 11931 8064 11940
rect 7656 11756 7708 11762
rect 7656 11698 7708 11704
rect 8300 11756 8352 11762
rect 8300 11698 8352 11704
rect 8312 11354 8340 11698
rect 8300 11348 8352 11354
rect 8300 11290 8352 11296
rect 7756 10908 8064 10917
rect 7756 10906 7762 10908
rect 7818 10906 7842 10908
rect 7898 10906 7922 10908
rect 7978 10906 8002 10908
rect 8058 10906 8064 10908
rect 7818 10854 7820 10906
rect 8000 10854 8002 10906
rect 7756 10852 7762 10854
rect 7818 10852 7842 10854
rect 7898 10852 7922 10854
rect 7978 10852 8002 10854
rect 8058 10852 8064 10854
rect 7756 10843 8064 10852
rect 8496 10198 8524 12294
rect 8576 12232 8628 12238
rect 8576 12174 8628 12180
rect 8484 10192 8536 10198
rect 8484 10134 8536 10140
rect 7564 10124 7616 10130
rect 7564 10066 7616 10072
rect 7576 9518 7604 10066
rect 8300 10056 8352 10062
rect 8300 9998 8352 10004
rect 7756 9820 8064 9829
rect 7756 9818 7762 9820
rect 7818 9818 7842 9820
rect 7898 9818 7922 9820
rect 7978 9818 8002 9820
rect 8058 9818 8064 9820
rect 7818 9766 7820 9818
rect 8000 9766 8002 9818
rect 7756 9764 7762 9766
rect 7818 9764 7842 9766
rect 7898 9764 7922 9766
rect 7978 9764 8002 9766
rect 8058 9764 8064 9766
rect 7756 9755 8064 9764
rect 8312 9654 8340 9998
rect 8300 9648 8352 9654
rect 8300 9590 8352 9596
rect 7564 9512 7616 9518
rect 7564 9454 7616 9460
rect 7576 7954 7604 9454
rect 8300 9444 8352 9450
rect 8300 9386 8352 9392
rect 7756 8732 8064 8741
rect 7756 8730 7762 8732
rect 7818 8730 7842 8732
rect 7898 8730 7922 8732
rect 7978 8730 8002 8732
rect 8058 8730 8064 8732
rect 7818 8678 7820 8730
rect 8000 8678 8002 8730
rect 7756 8676 7762 8678
rect 7818 8676 7842 8678
rect 7898 8676 7922 8678
rect 7978 8676 8002 8678
rect 8058 8676 8064 8678
rect 7756 8667 8064 8676
rect 7564 7948 7616 7954
rect 7564 7890 7616 7896
rect 5908 7336 5960 7342
rect 5908 7278 5960 7284
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 7288 7336 7340 7342
rect 7288 7278 7340 7284
rect 5500 7228 5580 7256
rect 5448 7210 5500 7216
rect 5172 6452 5224 6458
rect 5172 6394 5224 6400
rect 4436 6248 4488 6254
rect 4436 6190 4488 6196
rect 4988 6248 5040 6254
rect 4988 6190 5040 6196
rect 5080 6248 5132 6254
rect 5080 6190 5132 6196
rect 4448 5914 4476 6190
rect 5276 5914 5304 7210
rect 5448 6248 5500 6254
rect 5448 6190 5500 6196
rect 4344 5908 4396 5914
rect 4344 5850 4396 5856
rect 4436 5908 4488 5914
rect 4436 5850 4488 5856
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 4252 5772 4304 5778
rect 4252 5714 4304 5720
rect 4264 4758 4292 5714
rect 5080 5568 5132 5574
rect 5080 5510 5132 5516
rect 4656 5468 4964 5477
rect 4656 5466 4662 5468
rect 4718 5466 4742 5468
rect 4798 5466 4822 5468
rect 4878 5466 4902 5468
rect 4958 5466 4964 5468
rect 4718 5414 4720 5466
rect 4900 5414 4902 5466
rect 4656 5412 4662 5414
rect 4718 5412 4742 5414
rect 4798 5412 4822 5414
rect 4878 5412 4902 5414
rect 4958 5412 4964 5414
rect 4656 5403 4964 5412
rect 4528 5092 4580 5098
rect 4528 5034 4580 5040
rect 4540 4826 4568 5034
rect 4528 4820 4580 4826
rect 4528 4762 4580 4768
rect 4252 4752 4304 4758
rect 4252 4694 4304 4700
rect 4264 4010 4292 4694
rect 5092 4622 5120 5510
rect 5172 5024 5224 5030
rect 5172 4966 5224 4972
rect 4528 4616 4580 4622
rect 4528 4558 4580 4564
rect 5080 4616 5132 4622
rect 5080 4558 5132 4564
rect 4540 4282 4568 4558
rect 4656 4380 4964 4389
rect 4656 4378 4662 4380
rect 4718 4378 4742 4380
rect 4798 4378 4822 4380
rect 4878 4378 4902 4380
rect 4958 4378 4964 4380
rect 4718 4326 4720 4378
rect 4900 4326 4902 4378
rect 4656 4324 4662 4326
rect 4718 4324 4742 4326
rect 4798 4324 4822 4326
rect 4878 4324 4902 4326
rect 4958 4324 4964 4326
rect 4656 4315 4964 4324
rect 4528 4276 4580 4282
rect 4528 4218 4580 4224
rect 5092 4214 5120 4558
rect 5080 4208 5132 4214
rect 5080 4150 5132 4156
rect 5184 4146 5212 4966
rect 5264 4684 5316 4690
rect 5264 4626 5316 4632
rect 4712 4140 4764 4146
rect 4712 4082 4764 4088
rect 5172 4140 5224 4146
rect 5172 4082 5224 4088
rect 4252 4004 4304 4010
rect 4724 3992 4752 4082
rect 4252 3946 4304 3952
rect 4540 3964 4752 3992
rect 4264 3670 4292 3946
rect 4252 3664 4304 3670
rect 4252 3606 4304 3612
rect 4160 2576 4212 2582
rect 4160 2518 4212 2524
rect 4068 2440 4120 2446
rect 4068 2382 4120 2388
rect 4080 1970 4108 2382
rect 4172 2106 4200 2518
rect 4160 2100 4212 2106
rect 4160 2042 4212 2048
rect 4068 1964 4120 1970
rect 4068 1906 4120 1912
rect 3976 1896 4028 1902
rect 3976 1838 4028 1844
rect 2964 1760 3016 1766
rect 2964 1702 3016 1708
rect 940 1430 992 1436
rect 2700 1426 2820 1442
rect 2872 1488 2924 1494
rect 2872 1430 2924 1436
rect 2688 1420 2820 1426
rect 2740 1414 2820 1420
rect 2688 1362 2740 1368
rect 2792 1306 2820 1414
rect 2792 1290 2912 1306
rect 2792 1284 2924 1290
rect 2792 1278 2872 1284
rect 1556 1116 1864 1125
rect 1556 1114 1562 1116
rect 1618 1114 1642 1116
rect 1698 1114 1722 1116
rect 1778 1114 1802 1116
rect 1858 1114 1864 1116
rect 1618 1062 1620 1114
rect 1800 1062 1802 1114
rect 1556 1060 1562 1062
rect 1618 1060 1642 1062
rect 1698 1060 1722 1062
rect 1778 1060 1802 1062
rect 1858 1060 1864 1062
rect 1556 1051 1864 1060
rect 2792 882 2820 1278
rect 2872 1226 2924 1232
rect 2976 1018 3004 1702
rect 3106 1660 3414 1669
rect 3106 1658 3112 1660
rect 3168 1658 3192 1660
rect 3248 1658 3272 1660
rect 3328 1658 3352 1660
rect 3408 1658 3414 1660
rect 3168 1606 3170 1658
rect 3350 1606 3352 1658
rect 3106 1604 3112 1606
rect 3168 1604 3192 1606
rect 3248 1604 3272 1606
rect 3328 1604 3352 1606
rect 3408 1604 3414 1606
rect 3106 1595 3414 1604
rect 3988 1426 4016 1838
rect 4080 1766 4108 1906
rect 4540 1902 4568 3964
rect 5276 3738 5304 4626
rect 5460 4026 5488 6190
rect 5552 5778 5580 7228
rect 5920 5778 5948 7278
rect 6206 7100 6514 7109
rect 6206 7098 6212 7100
rect 6268 7098 6292 7100
rect 6348 7098 6372 7100
rect 6428 7098 6452 7100
rect 6508 7098 6514 7100
rect 6268 7046 6270 7098
rect 6450 7046 6452 7098
rect 6206 7044 6212 7046
rect 6268 7044 6292 7046
rect 6348 7044 6372 7046
rect 6428 7044 6452 7046
rect 6508 7044 6514 7046
rect 6206 7035 6514 7044
rect 6644 6928 6696 6934
rect 6644 6870 6696 6876
rect 6092 6452 6144 6458
rect 6092 6394 6144 6400
rect 5540 5772 5592 5778
rect 5540 5714 5592 5720
rect 5908 5772 5960 5778
rect 5908 5714 5960 5720
rect 5816 5364 5868 5370
rect 5816 5306 5868 5312
rect 5828 5098 5856 5306
rect 5816 5092 5868 5098
rect 5816 5034 5868 5040
rect 5460 3998 5580 4026
rect 5264 3732 5316 3738
rect 5264 3674 5316 3680
rect 4988 3596 5040 3602
rect 4988 3538 5040 3544
rect 4656 3292 4964 3301
rect 4656 3290 4662 3292
rect 4718 3290 4742 3292
rect 4798 3290 4822 3292
rect 4878 3290 4902 3292
rect 4958 3290 4964 3292
rect 4718 3238 4720 3290
rect 4900 3238 4902 3290
rect 4656 3236 4662 3238
rect 4718 3236 4742 3238
rect 4798 3236 4822 3238
rect 4878 3236 4902 3238
rect 4958 3236 4964 3238
rect 4656 3227 4964 3236
rect 5000 3194 5028 3538
rect 4988 3188 5040 3194
rect 4988 3130 5040 3136
rect 5552 2922 5580 3998
rect 5920 3058 5948 5714
rect 6104 3738 6132 6394
rect 6656 6186 6684 6870
rect 6840 6866 6868 7278
rect 7104 7200 7156 7206
rect 7104 7142 7156 7148
rect 7116 6934 7144 7142
rect 7104 6928 7156 6934
rect 7104 6870 7156 6876
rect 6828 6860 6880 6866
rect 6828 6802 6880 6808
rect 7300 6798 7328 7278
rect 7472 6860 7524 6866
rect 7472 6802 7524 6808
rect 7288 6792 7340 6798
rect 7288 6734 7340 6740
rect 6644 6180 6696 6186
rect 6644 6122 6696 6128
rect 6828 6180 6880 6186
rect 6828 6122 6880 6128
rect 6206 6012 6514 6021
rect 6206 6010 6212 6012
rect 6268 6010 6292 6012
rect 6348 6010 6372 6012
rect 6428 6010 6452 6012
rect 6508 6010 6514 6012
rect 6268 5958 6270 6010
rect 6450 5958 6452 6010
rect 6206 5956 6212 5958
rect 6268 5956 6292 5958
rect 6348 5956 6372 5958
rect 6428 5956 6452 5958
rect 6508 5956 6514 5958
rect 6206 5947 6514 5956
rect 6552 5704 6604 5710
rect 6552 5646 6604 5652
rect 6206 4924 6514 4933
rect 6206 4922 6212 4924
rect 6268 4922 6292 4924
rect 6348 4922 6372 4924
rect 6428 4922 6452 4924
rect 6508 4922 6514 4924
rect 6268 4870 6270 4922
rect 6450 4870 6452 4922
rect 6206 4868 6212 4870
rect 6268 4868 6292 4870
rect 6348 4868 6372 4870
rect 6428 4868 6452 4870
rect 6508 4868 6514 4870
rect 6206 4859 6514 4868
rect 6206 3836 6514 3845
rect 6206 3834 6212 3836
rect 6268 3834 6292 3836
rect 6348 3834 6372 3836
rect 6428 3834 6452 3836
rect 6508 3834 6514 3836
rect 6268 3782 6270 3834
rect 6450 3782 6452 3834
rect 6206 3780 6212 3782
rect 6268 3780 6292 3782
rect 6348 3780 6372 3782
rect 6428 3780 6452 3782
rect 6508 3780 6514 3782
rect 6206 3771 6514 3780
rect 6564 3738 6592 5646
rect 6736 5568 6788 5574
rect 6736 5510 6788 5516
rect 6644 5092 6696 5098
rect 6644 5034 6696 5040
rect 6656 4826 6684 5034
rect 6644 4820 6696 4826
rect 6644 4762 6696 4768
rect 6748 4622 6776 5510
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 6840 4486 6868 6122
rect 7288 4684 7340 4690
rect 7288 4626 7340 4632
rect 6828 4480 6880 4486
rect 6828 4422 6880 4428
rect 6092 3732 6144 3738
rect 6092 3674 6144 3680
rect 6552 3732 6604 3738
rect 6552 3674 6604 3680
rect 6644 3664 6696 3670
rect 6644 3606 6696 3612
rect 6656 3194 6684 3606
rect 6828 3596 6880 3602
rect 6828 3538 6880 3544
rect 6840 3194 6868 3538
rect 6644 3188 6696 3194
rect 6644 3130 6696 3136
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 6656 3058 6684 3130
rect 5908 3052 5960 3058
rect 5908 2994 5960 3000
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 5540 2916 5592 2922
rect 5540 2858 5592 2864
rect 5356 2848 5408 2854
rect 5356 2790 5408 2796
rect 5368 2650 5396 2790
rect 5552 2650 5580 2858
rect 6656 2774 6684 2994
rect 7300 2990 7328 4626
rect 7484 3942 7512 6802
rect 7576 5778 7604 7890
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 7756 7644 8064 7653
rect 7756 7642 7762 7644
rect 7818 7642 7842 7644
rect 7898 7642 7922 7644
rect 7978 7642 8002 7644
rect 8058 7642 8064 7644
rect 7818 7590 7820 7642
rect 8000 7590 8002 7642
rect 7756 7588 7762 7590
rect 7818 7588 7842 7590
rect 7898 7588 7922 7590
rect 7978 7588 8002 7590
rect 8058 7588 8064 7590
rect 7756 7579 8064 7588
rect 8116 7336 8168 7342
rect 8116 7278 8168 7284
rect 7656 7200 7708 7206
rect 7656 7142 7708 7148
rect 7668 6746 7696 7142
rect 7748 6792 7800 6798
rect 7668 6740 7748 6746
rect 7668 6734 7800 6740
rect 7668 6718 7788 6734
rect 7668 6254 7696 6718
rect 7756 6556 8064 6565
rect 7756 6554 7762 6556
rect 7818 6554 7842 6556
rect 7898 6554 7922 6556
rect 7978 6554 8002 6556
rect 8058 6554 8064 6556
rect 7818 6502 7820 6554
rect 8000 6502 8002 6554
rect 7756 6500 7762 6502
rect 7818 6500 7842 6502
rect 7898 6500 7922 6502
rect 7978 6500 8002 6502
rect 8058 6500 8064 6502
rect 7756 6491 8064 6500
rect 7656 6248 7708 6254
rect 7656 6190 7708 6196
rect 7668 5846 7696 6190
rect 8024 6112 8076 6118
rect 8024 6054 8076 6060
rect 8036 5846 8064 6054
rect 7656 5840 7708 5846
rect 7656 5782 7708 5788
rect 8024 5840 8076 5846
rect 8024 5782 8076 5788
rect 7564 5772 7616 5778
rect 7564 5714 7616 5720
rect 7576 5216 7604 5714
rect 7756 5468 8064 5477
rect 7756 5466 7762 5468
rect 7818 5466 7842 5468
rect 7898 5466 7922 5468
rect 7978 5466 8002 5468
rect 8058 5466 8064 5468
rect 7818 5414 7820 5466
rect 8000 5414 8002 5466
rect 7756 5412 7762 5414
rect 7818 5412 7842 5414
rect 7898 5412 7922 5414
rect 7978 5412 8002 5414
rect 8058 5412 8064 5414
rect 7756 5403 8064 5412
rect 8128 5386 8156 7278
rect 8220 7002 8248 7822
rect 8312 7342 8340 9386
rect 8496 9110 8524 10134
rect 8484 9104 8536 9110
rect 8484 9046 8536 9052
rect 8496 8022 8524 9046
rect 8484 8016 8536 8022
rect 8484 7958 8536 7964
rect 8588 7562 8616 12174
rect 8680 11626 8708 12582
rect 8668 11620 8720 11626
rect 8668 11562 8720 11568
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8404 7534 8616 7562
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 8208 6996 8260 7002
rect 8208 6938 8260 6944
rect 8312 6390 8340 7142
rect 8300 6384 8352 6390
rect 8300 6326 8352 6332
rect 8128 5358 8248 5386
rect 7656 5228 7708 5234
rect 7576 5188 7656 5216
rect 7656 5170 7708 5176
rect 8116 5228 8168 5234
rect 8116 5170 8168 5176
rect 7756 4380 8064 4389
rect 7756 4378 7762 4380
rect 7818 4378 7842 4380
rect 7898 4378 7922 4380
rect 7978 4378 8002 4380
rect 8058 4378 8064 4380
rect 7818 4326 7820 4378
rect 8000 4326 8002 4378
rect 7756 4324 7762 4326
rect 7818 4324 7842 4326
rect 7898 4324 7922 4326
rect 7978 4324 8002 4326
rect 8058 4324 8064 4326
rect 7756 4315 8064 4324
rect 7472 3936 7524 3942
rect 7472 3878 7524 3884
rect 7756 3292 8064 3301
rect 7756 3290 7762 3292
rect 7818 3290 7842 3292
rect 7898 3290 7922 3292
rect 7978 3290 8002 3292
rect 8058 3290 8064 3292
rect 7818 3238 7820 3290
rect 8000 3238 8002 3290
rect 7756 3236 7762 3238
rect 7818 3236 7842 3238
rect 7898 3236 7922 3238
rect 7978 3236 8002 3238
rect 8058 3236 8064 3238
rect 7756 3227 8064 3236
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 7288 2984 7340 2990
rect 7288 2926 7340 2932
rect 6206 2748 6514 2757
rect 6206 2746 6212 2748
rect 6268 2746 6292 2748
rect 6348 2746 6372 2748
rect 6428 2746 6452 2748
rect 6508 2746 6514 2748
rect 6268 2694 6270 2746
rect 6450 2694 6452 2746
rect 6206 2692 6212 2694
rect 6268 2692 6292 2694
rect 6348 2692 6372 2694
rect 6428 2692 6452 2694
rect 6508 2692 6514 2694
rect 6206 2683 6514 2692
rect 6564 2746 6684 2774
rect 5356 2644 5408 2650
rect 5356 2586 5408 2592
rect 5540 2644 5592 2650
rect 5540 2586 5592 2592
rect 5632 2508 5684 2514
rect 5632 2450 5684 2456
rect 4656 2204 4964 2213
rect 4656 2202 4662 2204
rect 4718 2202 4742 2204
rect 4798 2202 4822 2204
rect 4878 2202 4902 2204
rect 4958 2202 4964 2204
rect 4718 2150 4720 2202
rect 4900 2150 4902 2202
rect 4656 2148 4662 2150
rect 4718 2148 4742 2150
rect 4798 2148 4822 2150
rect 4878 2148 4902 2150
rect 4958 2148 4964 2150
rect 4656 2139 4964 2148
rect 4528 1896 4580 1902
rect 4528 1838 4580 1844
rect 5172 1896 5224 1902
rect 5172 1838 5224 1844
rect 4068 1760 4120 1766
rect 4068 1702 4120 1708
rect 3976 1420 4028 1426
rect 3976 1362 4028 1368
rect 2964 1012 3016 1018
rect 2964 954 3016 960
rect 2780 876 2832 882
rect 2780 818 2832 824
rect 3988 814 4016 1362
rect 4080 1358 4108 1702
rect 4540 1442 4568 1838
rect 4540 1414 4660 1442
rect 4632 1358 4660 1414
rect 4068 1352 4120 1358
rect 4068 1294 4120 1300
rect 4620 1352 4672 1358
rect 4620 1294 4672 1300
rect 5184 1290 5212 1838
rect 5644 1562 5672 2450
rect 6206 1660 6514 1669
rect 6206 1658 6212 1660
rect 6268 1658 6292 1660
rect 6348 1658 6372 1660
rect 6428 1658 6452 1660
rect 6508 1658 6514 1660
rect 6268 1606 6270 1658
rect 6450 1606 6452 1658
rect 6206 1604 6212 1606
rect 6268 1604 6292 1606
rect 6348 1604 6372 1606
rect 6428 1604 6452 1606
rect 6508 1604 6514 1606
rect 6206 1595 6514 1604
rect 5632 1556 5684 1562
rect 5632 1498 5684 1504
rect 6564 1494 6592 2746
rect 7300 2038 7328 2926
rect 7576 2378 7604 2994
rect 7564 2372 7616 2378
rect 7564 2314 7616 2320
rect 7288 2032 7340 2038
rect 7288 1974 7340 1980
rect 7300 1494 7328 1974
rect 7576 1766 7604 2314
rect 7756 2204 8064 2213
rect 7756 2202 7762 2204
rect 7818 2202 7842 2204
rect 7898 2202 7922 2204
rect 7978 2202 8002 2204
rect 8058 2202 8064 2204
rect 7818 2150 7820 2202
rect 8000 2150 8002 2202
rect 7756 2148 7762 2150
rect 7818 2148 7842 2150
rect 7898 2148 7922 2150
rect 7978 2148 8002 2150
rect 8058 2148 8064 2150
rect 7756 2139 8064 2148
rect 7564 1760 7616 1766
rect 7564 1702 7616 1708
rect 6552 1488 6604 1494
rect 6552 1430 6604 1436
rect 7288 1488 7340 1494
rect 7288 1430 7340 1436
rect 8128 1426 8156 5170
rect 8220 4214 8248 5358
rect 8208 4208 8260 4214
rect 8208 4150 8260 4156
rect 8208 4004 8260 4010
rect 8208 3946 8260 3952
rect 8220 2650 8248 3946
rect 8208 2644 8260 2650
rect 8208 2586 8260 2592
rect 8404 1970 8432 7534
rect 8680 7410 8708 7686
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 8588 6254 8616 6598
rect 8576 6248 8628 6254
rect 8576 6190 8628 6196
rect 8484 5840 8536 5846
rect 8484 5782 8536 5788
rect 8496 5098 8524 5782
rect 8484 5092 8536 5098
rect 8484 5034 8536 5040
rect 8484 3936 8536 3942
rect 8484 3878 8536 3884
rect 8496 3738 8524 3878
rect 8484 3732 8536 3738
rect 8484 3674 8536 3680
rect 8496 2582 8524 3674
rect 8484 2576 8536 2582
rect 8484 2518 8536 2524
rect 8576 2508 8628 2514
rect 8576 2450 8628 2456
rect 8392 1964 8444 1970
rect 8392 1906 8444 1912
rect 5264 1420 5316 1426
rect 5264 1362 5316 1368
rect 8116 1420 8168 1426
rect 8116 1362 8168 1368
rect 5172 1284 5224 1290
rect 5172 1226 5224 1232
rect 4656 1116 4964 1125
rect 4656 1114 4662 1116
rect 4718 1114 4742 1116
rect 4798 1114 4822 1116
rect 4878 1114 4902 1116
rect 4958 1114 4964 1116
rect 4718 1062 4720 1114
rect 4900 1062 4902 1114
rect 4656 1060 4662 1062
rect 4718 1060 4742 1062
rect 4798 1060 4822 1062
rect 4878 1060 4902 1062
rect 4958 1060 4964 1062
rect 4656 1051 4964 1060
rect 5184 950 5212 1226
rect 5276 1018 5304 1362
rect 5448 1352 5500 1358
rect 5448 1294 5500 1300
rect 5264 1012 5316 1018
rect 5264 954 5316 960
rect 5172 944 5224 950
rect 5172 886 5224 892
rect 5460 814 5488 1294
rect 8588 1290 8616 2450
rect 8680 1902 8708 7346
rect 8864 6730 8892 13262
rect 8956 12714 8984 13738
rect 9048 12986 9076 14826
rect 9306 14716 9614 14725
rect 9306 14714 9312 14716
rect 9368 14714 9392 14716
rect 9448 14714 9472 14716
rect 9528 14714 9552 14716
rect 9608 14714 9614 14716
rect 9368 14662 9370 14714
rect 9550 14662 9552 14714
rect 9306 14660 9312 14662
rect 9368 14660 9392 14662
rect 9448 14660 9472 14662
rect 9528 14660 9552 14662
rect 9608 14660 9614 14662
rect 9306 14651 9614 14660
rect 10152 14074 10180 15302
rect 10336 14822 10364 16680
rect 10856 16348 11164 16357
rect 10856 16346 10862 16348
rect 10918 16346 10942 16348
rect 10998 16346 11022 16348
rect 11078 16346 11102 16348
rect 11158 16346 11164 16348
rect 10918 16294 10920 16346
rect 11100 16294 11102 16346
rect 10856 16292 10862 16294
rect 10918 16292 10942 16294
rect 10998 16292 11022 16294
rect 11078 16292 11102 16294
rect 11158 16292 11164 16294
rect 10856 16283 11164 16292
rect 11348 16250 11376 18090
rect 11336 16244 11388 16250
rect 11336 16186 11388 16192
rect 11336 15496 11388 15502
rect 11336 15438 11388 15444
rect 10856 15260 11164 15269
rect 10856 15258 10862 15260
rect 10918 15258 10942 15260
rect 10998 15258 11022 15260
rect 11078 15258 11102 15260
rect 11158 15258 11164 15260
rect 10918 15206 10920 15258
rect 11100 15206 11102 15258
rect 10856 15204 10862 15206
rect 10918 15204 10942 15206
rect 10998 15204 11022 15206
rect 11078 15204 11102 15206
rect 11158 15204 11164 15206
rect 10856 15195 11164 15204
rect 11244 14952 11296 14958
rect 11244 14894 11296 14900
rect 10324 14816 10376 14822
rect 10324 14758 10376 14764
rect 11152 14816 11204 14822
rect 11152 14758 11204 14764
rect 10140 14068 10192 14074
rect 10140 14010 10192 14016
rect 9306 13628 9614 13637
rect 9306 13626 9312 13628
rect 9368 13626 9392 13628
rect 9448 13626 9472 13628
rect 9528 13626 9552 13628
rect 9608 13626 9614 13628
rect 9368 13574 9370 13626
rect 9550 13574 9552 13626
rect 9306 13572 9312 13574
rect 9368 13572 9392 13574
rect 9448 13572 9472 13574
rect 9528 13572 9552 13574
rect 9608 13572 9614 13574
rect 9306 13563 9614 13572
rect 9312 13320 9364 13326
rect 9232 13268 9312 13274
rect 9232 13262 9364 13268
rect 9232 13246 9352 13262
rect 9036 12980 9088 12986
rect 9036 12922 9088 12928
rect 9232 12850 9260 13246
rect 9220 12844 9272 12850
rect 9220 12786 9272 12792
rect 8944 12708 8996 12714
rect 8944 12650 8996 12656
rect 8956 11626 8984 12650
rect 9232 11762 9260 12786
rect 9956 12708 10008 12714
rect 9956 12650 10008 12656
rect 9306 12540 9614 12549
rect 9306 12538 9312 12540
rect 9368 12538 9392 12540
rect 9448 12538 9472 12540
rect 9528 12538 9552 12540
rect 9608 12538 9614 12540
rect 9368 12486 9370 12538
rect 9550 12486 9552 12538
rect 9306 12484 9312 12486
rect 9368 12484 9392 12486
rect 9448 12484 9472 12486
rect 9528 12484 9552 12486
rect 9608 12484 9614 12486
rect 9306 12475 9614 12484
rect 9220 11756 9272 11762
rect 9220 11698 9272 11704
rect 8944 11620 8996 11626
rect 8944 11562 8996 11568
rect 9968 11558 9996 12650
rect 9956 11552 10008 11558
rect 9956 11494 10008 11500
rect 9306 11452 9614 11461
rect 9306 11450 9312 11452
rect 9368 11450 9392 11452
rect 9448 11450 9472 11452
rect 9528 11450 9552 11452
rect 9608 11450 9614 11452
rect 9368 11398 9370 11450
rect 9550 11398 9552 11450
rect 9306 11396 9312 11398
rect 9368 11396 9392 11398
rect 9448 11396 9472 11398
rect 9528 11396 9552 11398
rect 9608 11396 9614 11398
rect 9306 11387 9614 11396
rect 10336 11286 10364 14758
rect 11164 14414 11192 14758
rect 11256 14482 11284 14894
rect 11348 14550 11376 15438
rect 11440 14618 11468 18090
rect 12268 17882 12296 18142
rect 12406 17980 12714 17989
rect 12406 17978 12412 17980
rect 12468 17978 12492 17980
rect 12548 17978 12572 17980
rect 12628 17978 12652 17980
rect 12708 17978 12714 17980
rect 12468 17926 12470 17978
rect 12650 17926 12652 17978
rect 12406 17924 12412 17926
rect 12468 17924 12492 17926
rect 12548 17924 12572 17926
rect 12628 17924 12652 17926
rect 12708 17924 12714 17926
rect 12406 17915 12714 17924
rect 12256 17876 12308 17882
rect 12256 17818 12308 17824
rect 12256 17740 12308 17746
rect 12256 17682 12308 17688
rect 11980 17536 12032 17542
rect 11980 17478 12032 17484
rect 11992 15638 12020 17478
rect 12164 16788 12216 16794
rect 12164 16730 12216 16736
rect 12072 16448 12124 16454
rect 12072 16390 12124 16396
rect 12084 16114 12112 16390
rect 12072 16108 12124 16114
rect 12072 16050 12124 16056
rect 11980 15632 12032 15638
rect 11980 15574 12032 15580
rect 11520 14952 11572 14958
rect 11520 14894 11572 14900
rect 11428 14612 11480 14618
rect 11428 14554 11480 14560
rect 11336 14544 11388 14550
rect 11336 14486 11388 14492
rect 11244 14476 11296 14482
rect 11244 14418 11296 14424
rect 11152 14408 11204 14414
rect 11152 14350 11204 14356
rect 10856 14172 11164 14181
rect 10856 14170 10862 14172
rect 10918 14170 10942 14172
rect 10998 14170 11022 14172
rect 11078 14170 11102 14172
rect 11158 14170 11164 14172
rect 10918 14118 10920 14170
rect 11100 14118 11102 14170
rect 10856 14116 10862 14118
rect 10918 14116 10942 14118
rect 10998 14116 11022 14118
rect 11078 14116 11102 14118
rect 11158 14116 11164 14118
rect 10856 14107 11164 14116
rect 11256 13530 11284 14418
rect 11348 14414 11376 14486
rect 11336 14408 11388 14414
rect 11336 14350 11388 14356
rect 11244 13524 11296 13530
rect 11244 13466 11296 13472
rect 10856 13084 11164 13093
rect 10856 13082 10862 13084
rect 10918 13082 10942 13084
rect 10998 13082 11022 13084
rect 11078 13082 11102 13084
rect 11158 13082 11164 13084
rect 10918 13030 10920 13082
rect 11100 13030 11102 13082
rect 10856 13028 10862 13030
rect 10918 13028 10942 13030
rect 10998 13028 11022 13030
rect 11078 13028 11102 13030
rect 11158 13028 11164 13030
rect 10856 13019 11164 13028
rect 11152 12776 11204 12782
rect 11152 12718 11204 12724
rect 11164 12374 11192 12718
rect 11152 12368 11204 12374
rect 11152 12310 11204 12316
rect 10600 12300 10652 12306
rect 10600 12242 10652 12248
rect 10784 12300 10836 12306
rect 10784 12242 10836 12248
rect 10612 11354 10640 12242
rect 10796 11830 10824 12242
rect 10856 11996 11164 12005
rect 10856 11994 10862 11996
rect 10918 11994 10942 11996
rect 10998 11994 11022 11996
rect 11078 11994 11102 11996
rect 11158 11994 11164 11996
rect 10918 11942 10920 11994
rect 11100 11942 11102 11994
rect 10856 11940 10862 11942
rect 10918 11940 10942 11942
rect 10998 11940 11022 11942
rect 11078 11940 11102 11942
rect 11158 11940 11164 11942
rect 10856 11931 11164 11940
rect 10784 11824 10836 11830
rect 10784 11766 10836 11772
rect 11336 11688 11388 11694
rect 11336 11630 11388 11636
rect 10600 11348 10652 11354
rect 10600 11290 10652 11296
rect 10324 11280 10376 11286
rect 10324 11222 10376 11228
rect 11348 11218 11376 11630
rect 11336 11212 11388 11218
rect 11336 11154 11388 11160
rect 10856 10908 11164 10917
rect 10856 10906 10862 10908
rect 10918 10906 10942 10908
rect 10998 10906 11022 10908
rect 11078 10906 11102 10908
rect 11158 10906 11164 10908
rect 10918 10854 10920 10906
rect 11100 10854 11102 10906
rect 10856 10852 10862 10854
rect 10918 10852 10942 10854
rect 10998 10852 11022 10854
rect 11078 10852 11102 10854
rect 11158 10852 11164 10854
rect 10856 10843 11164 10852
rect 10048 10600 10100 10606
rect 10048 10542 10100 10548
rect 9306 10364 9614 10373
rect 9306 10362 9312 10364
rect 9368 10362 9392 10364
rect 9448 10362 9472 10364
rect 9528 10362 9552 10364
rect 9608 10362 9614 10364
rect 9368 10310 9370 10362
rect 9550 10310 9552 10362
rect 9306 10308 9312 10310
rect 9368 10308 9392 10310
rect 9448 10308 9472 10310
rect 9528 10308 9552 10310
rect 9608 10308 9614 10310
rect 9306 10299 9614 10308
rect 9036 9920 9088 9926
rect 9036 9862 9088 9868
rect 9048 9518 9076 9862
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 9036 9376 9088 9382
rect 9036 9318 9088 9324
rect 9048 7478 9076 9318
rect 9306 9276 9614 9285
rect 9306 9274 9312 9276
rect 9368 9274 9392 9276
rect 9448 9274 9472 9276
rect 9528 9274 9552 9276
rect 9608 9274 9614 9276
rect 9368 9222 9370 9274
rect 9550 9222 9552 9274
rect 9306 9220 9312 9222
rect 9368 9220 9392 9222
rect 9448 9220 9472 9222
rect 9528 9220 9552 9222
rect 9608 9220 9614 9222
rect 9306 9211 9614 9220
rect 10060 8838 10088 10542
rect 10508 10532 10560 10538
rect 10508 10474 10560 10480
rect 10140 10464 10192 10470
rect 10140 10406 10192 10412
rect 10152 10130 10180 10406
rect 10520 10130 10548 10474
rect 10140 10124 10192 10130
rect 10140 10066 10192 10072
rect 10508 10124 10560 10130
rect 10508 10066 10560 10072
rect 11348 9994 11376 11154
rect 11440 10198 11468 14554
rect 11532 14074 11560 14894
rect 11888 14884 11940 14890
rect 11888 14826 11940 14832
rect 11900 14618 11928 14826
rect 11888 14612 11940 14618
rect 11888 14554 11940 14560
rect 11796 14272 11848 14278
rect 11796 14214 11848 14220
rect 11520 14068 11572 14074
rect 11520 14010 11572 14016
rect 11808 13870 11836 14214
rect 11796 13864 11848 13870
rect 11796 13806 11848 13812
rect 11520 12776 11572 12782
rect 11520 12718 11572 12724
rect 11532 12442 11560 12718
rect 11900 12714 11928 14554
rect 11992 13462 12020 15574
rect 12176 15502 12204 16730
rect 12164 15496 12216 15502
rect 12164 15438 12216 15444
rect 12176 14482 12204 15438
rect 12164 14476 12216 14482
rect 12164 14418 12216 14424
rect 12268 14006 12296 17682
rect 12406 16892 12714 16901
rect 12406 16890 12412 16892
rect 12468 16890 12492 16892
rect 12548 16890 12572 16892
rect 12628 16890 12652 16892
rect 12708 16890 12714 16892
rect 12468 16838 12470 16890
rect 12650 16838 12652 16890
rect 12406 16836 12412 16838
rect 12468 16836 12492 16838
rect 12548 16836 12572 16838
rect 12628 16836 12652 16838
rect 12708 16836 12714 16838
rect 12406 16827 12714 16836
rect 12532 16720 12584 16726
rect 12532 16662 12584 16668
rect 12544 15978 12572 16662
rect 12820 16574 12848 19200
rect 13956 18524 14264 18533
rect 13956 18522 13962 18524
rect 14018 18522 14042 18524
rect 14098 18522 14122 18524
rect 14178 18522 14202 18524
rect 14258 18522 14264 18524
rect 14018 18470 14020 18522
rect 14200 18470 14202 18522
rect 13956 18468 13962 18470
rect 14018 18468 14042 18470
rect 14098 18468 14122 18470
rect 14178 18468 14202 18470
rect 14258 18468 14264 18470
rect 13956 18459 14264 18468
rect 13452 18080 13504 18086
rect 13452 18022 13504 18028
rect 13084 17808 13136 17814
rect 13084 17750 13136 17756
rect 13096 17066 13124 17750
rect 13084 17060 13136 17066
rect 13084 17002 13136 17008
rect 13096 16726 13124 17002
rect 13084 16720 13136 16726
rect 13084 16662 13136 16668
rect 12820 16546 12940 16574
rect 12716 16448 12768 16454
rect 12716 16390 12768 16396
rect 12728 15994 12756 16390
rect 12532 15972 12584 15978
rect 12728 15966 12848 15994
rect 12532 15914 12584 15920
rect 12406 15804 12714 15813
rect 12406 15802 12412 15804
rect 12468 15802 12492 15804
rect 12548 15802 12572 15804
rect 12628 15802 12652 15804
rect 12708 15802 12714 15804
rect 12468 15750 12470 15802
rect 12650 15750 12652 15802
rect 12406 15748 12412 15750
rect 12468 15748 12492 15750
rect 12548 15748 12572 15750
rect 12628 15748 12652 15750
rect 12708 15748 12714 15750
rect 12406 15739 12714 15748
rect 12820 15706 12848 15966
rect 12912 15706 12940 16546
rect 13096 15978 13124 16662
rect 13084 15972 13136 15978
rect 13084 15914 13136 15920
rect 12808 15700 12860 15706
rect 12808 15642 12860 15648
rect 12900 15700 12952 15706
rect 12900 15642 12952 15648
rect 13096 15638 13124 15914
rect 13084 15632 13136 15638
rect 13084 15574 13136 15580
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 12406 14716 12714 14725
rect 12406 14714 12412 14716
rect 12468 14714 12492 14716
rect 12548 14714 12572 14716
rect 12628 14714 12652 14716
rect 12708 14714 12714 14716
rect 12468 14662 12470 14714
rect 12650 14662 12652 14714
rect 12406 14660 12412 14662
rect 12468 14660 12492 14662
rect 12548 14660 12572 14662
rect 12628 14660 12652 14662
rect 12708 14660 12714 14662
rect 12406 14651 12714 14660
rect 12820 14482 12848 14758
rect 13096 14550 13124 15574
rect 13464 14958 13492 18022
rect 13820 17672 13872 17678
rect 13820 17614 13872 17620
rect 14740 17672 14792 17678
rect 14740 17614 14792 17620
rect 15108 17672 15160 17678
rect 15108 17614 15160 17620
rect 13452 14952 13504 14958
rect 13452 14894 13504 14900
rect 13084 14544 13136 14550
rect 13084 14486 13136 14492
rect 12808 14476 12860 14482
rect 12808 14418 12860 14424
rect 12900 14272 12952 14278
rect 12900 14214 12952 14220
rect 12256 14000 12308 14006
rect 12256 13942 12308 13948
rect 12808 13864 12860 13870
rect 12808 13806 12860 13812
rect 12406 13628 12714 13637
rect 12406 13626 12412 13628
rect 12468 13626 12492 13628
rect 12548 13626 12572 13628
rect 12628 13626 12652 13628
rect 12708 13626 12714 13628
rect 12468 13574 12470 13626
rect 12650 13574 12652 13626
rect 12406 13572 12412 13574
rect 12468 13572 12492 13574
rect 12548 13572 12572 13574
rect 12628 13572 12652 13574
rect 12708 13572 12714 13574
rect 12406 13563 12714 13572
rect 11980 13456 12032 13462
rect 11980 13398 12032 13404
rect 12820 12986 12848 13806
rect 12808 12980 12860 12986
rect 12808 12922 12860 12928
rect 12912 12714 12940 14214
rect 13832 13802 13860 17614
rect 14280 17604 14332 17610
rect 14280 17546 14332 17552
rect 13956 17436 14264 17445
rect 13956 17434 13962 17436
rect 14018 17434 14042 17436
rect 14098 17434 14122 17436
rect 14178 17434 14202 17436
rect 14258 17434 14264 17436
rect 14018 17382 14020 17434
rect 14200 17382 14202 17434
rect 13956 17380 13962 17382
rect 14018 17380 14042 17382
rect 14098 17380 14122 17382
rect 14178 17380 14202 17382
rect 14258 17380 14264 17382
rect 13956 17371 14264 17380
rect 14292 16726 14320 17546
rect 14752 17202 14780 17614
rect 14740 17196 14792 17202
rect 14740 17138 14792 17144
rect 14280 16720 14332 16726
rect 14280 16662 14332 16668
rect 13956 16348 14264 16357
rect 13956 16346 13962 16348
rect 14018 16346 14042 16348
rect 14098 16346 14122 16348
rect 14178 16346 14202 16348
rect 14258 16346 14264 16348
rect 14018 16294 14020 16346
rect 14200 16294 14202 16346
rect 13956 16292 13962 16294
rect 14018 16292 14042 16294
rect 14098 16292 14122 16294
rect 14178 16292 14202 16294
rect 14258 16292 14264 16294
rect 13956 16283 14264 16292
rect 15120 15706 15148 17614
rect 15200 15972 15252 15978
rect 15200 15914 15252 15920
rect 14280 15700 14332 15706
rect 14280 15642 14332 15648
rect 15108 15700 15160 15706
rect 15108 15642 15160 15648
rect 13956 15260 14264 15269
rect 13956 15258 13962 15260
rect 14018 15258 14042 15260
rect 14098 15258 14122 15260
rect 14178 15258 14202 15260
rect 14258 15258 14264 15260
rect 14018 15206 14020 15258
rect 14200 15206 14202 15258
rect 13956 15204 13962 15206
rect 14018 15204 14042 15206
rect 14098 15204 14122 15206
rect 14178 15204 14202 15206
rect 14258 15204 14264 15206
rect 13956 15195 14264 15204
rect 14292 15026 14320 15642
rect 15212 15586 15240 15914
rect 15292 15904 15344 15910
rect 15292 15846 15344 15852
rect 15120 15558 15240 15586
rect 15016 15496 15068 15502
rect 15016 15438 15068 15444
rect 14280 15020 14332 15026
rect 14280 14962 14332 14968
rect 15028 14482 15056 15438
rect 15120 15366 15148 15558
rect 15108 15360 15160 15366
rect 15108 15302 15160 15308
rect 15016 14476 15068 14482
rect 15016 14418 15068 14424
rect 15120 14362 15148 15302
rect 15200 14408 15252 14414
rect 15120 14356 15200 14362
rect 15120 14350 15252 14356
rect 15120 14334 15240 14350
rect 15016 14272 15068 14278
rect 15016 14214 15068 14220
rect 13956 14172 14264 14181
rect 13956 14170 13962 14172
rect 14018 14170 14042 14172
rect 14098 14170 14122 14172
rect 14178 14170 14202 14172
rect 14258 14170 14264 14172
rect 14018 14118 14020 14170
rect 14200 14118 14202 14170
rect 13956 14116 13962 14118
rect 14018 14116 14042 14118
rect 14098 14116 14122 14118
rect 14178 14116 14202 14118
rect 14258 14116 14264 14118
rect 13956 14107 14264 14116
rect 14280 14000 14332 14006
rect 14280 13942 14332 13948
rect 13728 13796 13780 13802
rect 13728 13738 13780 13744
rect 13820 13796 13872 13802
rect 13820 13738 13872 13744
rect 13740 12782 13768 13738
rect 13832 13530 13860 13738
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 13832 12850 13860 13466
rect 13956 13084 14264 13093
rect 13956 13082 13962 13084
rect 14018 13082 14042 13084
rect 14098 13082 14122 13084
rect 14178 13082 14202 13084
rect 14258 13082 14264 13084
rect 14018 13030 14020 13082
rect 14200 13030 14202 13082
rect 13956 13028 13962 13030
rect 14018 13028 14042 13030
rect 14098 13028 14122 13030
rect 14178 13028 14202 13030
rect 14258 13028 14264 13030
rect 13956 13019 14264 13028
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13728 12776 13780 12782
rect 13728 12718 13780 12724
rect 11888 12708 11940 12714
rect 11888 12650 11940 12656
rect 12900 12708 12952 12714
rect 12900 12650 12952 12656
rect 12256 12640 12308 12646
rect 12256 12582 12308 12588
rect 12268 12442 12296 12582
rect 12406 12540 12714 12549
rect 12406 12538 12412 12540
rect 12468 12538 12492 12540
rect 12548 12538 12572 12540
rect 12628 12538 12652 12540
rect 12708 12538 12714 12540
rect 12468 12486 12470 12538
rect 12650 12486 12652 12538
rect 12406 12484 12412 12486
rect 12468 12484 12492 12486
rect 12548 12484 12572 12486
rect 12628 12484 12652 12486
rect 12708 12484 12714 12486
rect 12406 12475 12714 12484
rect 11520 12436 11572 12442
rect 11520 12378 11572 12384
rect 12256 12436 12308 12442
rect 12256 12378 12308 12384
rect 12912 12306 12940 12650
rect 12900 12300 12952 12306
rect 12900 12242 12952 12248
rect 11612 12096 11664 12102
rect 11612 12038 11664 12044
rect 11624 11694 11652 12038
rect 11704 11824 11756 11830
rect 11704 11766 11756 11772
rect 11612 11688 11664 11694
rect 11612 11630 11664 11636
rect 11624 11286 11652 11630
rect 11612 11280 11664 11286
rect 11612 11222 11664 11228
rect 11716 11150 11744 11766
rect 11796 11756 11848 11762
rect 11796 11698 11848 11704
rect 11808 11218 11836 11698
rect 12406 11452 12714 11461
rect 12406 11450 12412 11452
rect 12468 11450 12492 11452
rect 12548 11450 12572 11452
rect 12628 11450 12652 11452
rect 12708 11450 12714 11452
rect 12468 11398 12470 11450
rect 12650 11398 12652 11450
rect 12406 11396 12412 11398
rect 12468 11396 12492 11398
rect 12548 11396 12572 11398
rect 12628 11396 12652 11398
rect 12708 11396 12714 11398
rect 12406 11387 12714 11396
rect 13740 11218 13768 12718
rect 13832 12374 13860 12786
rect 13820 12368 13872 12374
rect 13820 12310 13872 12316
rect 14292 12170 14320 13942
rect 14832 13864 14884 13870
rect 14832 13806 14884 13812
rect 14924 13864 14976 13870
rect 14924 13806 14976 13812
rect 14740 13728 14792 13734
rect 14740 13670 14792 13676
rect 14648 13456 14700 13462
rect 14648 13398 14700 13404
rect 14372 13388 14424 13394
rect 14372 13330 14424 13336
rect 13820 12164 13872 12170
rect 13820 12106 13872 12112
rect 14280 12164 14332 12170
rect 14280 12106 14332 12112
rect 11796 11212 11848 11218
rect 11796 11154 11848 11160
rect 13728 11212 13780 11218
rect 13728 11154 13780 11160
rect 11704 11144 11756 11150
rect 11704 11086 11756 11092
rect 11428 10192 11480 10198
rect 11428 10134 11480 10140
rect 11336 9988 11388 9994
rect 11336 9930 11388 9936
rect 10856 9820 11164 9829
rect 10856 9818 10862 9820
rect 10918 9818 10942 9820
rect 10998 9818 11022 9820
rect 11078 9818 11102 9820
rect 11158 9818 11164 9820
rect 10918 9766 10920 9818
rect 11100 9766 11102 9818
rect 10856 9764 10862 9766
rect 10918 9764 10942 9766
rect 10998 9764 11022 9766
rect 11078 9764 11102 9766
rect 11158 9764 11164 9766
rect 10856 9755 11164 9764
rect 11244 8968 11296 8974
rect 11244 8910 11296 8916
rect 10048 8832 10100 8838
rect 10048 8774 10100 8780
rect 9306 8188 9614 8197
rect 9306 8186 9312 8188
rect 9368 8186 9392 8188
rect 9448 8186 9472 8188
rect 9528 8186 9552 8188
rect 9608 8186 9614 8188
rect 9368 8134 9370 8186
rect 9550 8134 9552 8186
rect 9306 8132 9312 8134
rect 9368 8132 9392 8134
rect 9448 8132 9472 8134
rect 9528 8132 9552 8134
rect 9608 8132 9614 8134
rect 9306 8123 9614 8132
rect 9312 7744 9364 7750
rect 9312 7686 9364 7692
rect 9036 7472 9088 7478
rect 9036 7414 9088 7420
rect 9324 7410 9352 7686
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 8944 7336 8996 7342
rect 8996 7296 9076 7324
rect 8944 7278 8996 7284
rect 8944 7200 8996 7206
rect 8944 7142 8996 7148
rect 8852 6724 8904 6730
rect 8852 6666 8904 6672
rect 8956 6662 8984 7142
rect 8944 6656 8996 6662
rect 8944 6598 8996 6604
rect 8956 6458 8984 6598
rect 8944 6452 8996 6458
rect 8944 6394 8996 6400
rect 8760 6316 8812 6322
rect 8760 6258 8812 6264
rect 8772 3942 8800 6258
rect 9048 4010 9076 7296
rect 9220 7268 9272 7274
rect 9220 7210 9272 7216
rect 9128 7200 9180 7206
rect 9128 7142 9180 7148
rect 9140 5234 9168 7142
rect 9232 6866 9260 7210
rect 9306 7100 9614 7109
rect 9306 7098 9312 7100
rect 9368 7098 9392 7100
rect 9448 7098 9472 7100
rect 9528 7098 9552 7100
rect 9608 7098 9614 7100
rect 9368 7046 9370 7098
rect 9550 7046 9552 7098
rect 9306 7044 9312 7046
rect 9368 7044 9392 7046
rect 9448 7044 9472 7046
rect 9528 7044 9552 7046
rect 9608 7044 9614 7046
rect 9306 7035 9614 7044
rect 9220 6860 9272 6866
rect 9220 6802 9272 6808
rect 9232 5574 9260 6802
rect 10060 6798 10088 8774
rect 10856 8732 11164 8741
rect 10856 8730 10862 8732
rect 10918 8730 10942 8732
rect 10998 8730 11022 8732
rect 11078 8730 11102 8732
rect 11158 8730 11164 8732
rect 10918 8678 10920 8730
rect 11100 8678 11102 8730
rect 10856 8676 10862 8678
rect 10918 8676 10942 8678
rect 10998 8676 11022 8678
rect 11078 8676 11102 8678
rect 11158 8676 11164 8678
rect 10856 8667 11164 8676
rect 11256 8634 11284 8910
rect 11244 8628 11296 8634
rect 11244 8570 11296 8576
rect 11348 8514 11376 9930
rect 11440 9382 11468 10134
rect 11428 9376 11480 9382
rect 11428 9318 11480 9324
rect 11256 8486 11376 8514
rect 11256 8022 11284 8486
rect 11336 8424 11388 8430
rect 11336 8366 11388 8372
rect 11244 8016 11296 8022
rect 11244 7958 11296 7964
rect 10784 7948 10836 7954
rect 10784 7890 10836 7896
rect 10796 7002 10824 7890
rect 11348 7818 11376 8366
rect 11336 7812 11388 7818
rect 11336 7754 11388 7760
rect 10856 7644 11164 7653
rect 10856 7642 10862 7644
rect 10918 7642 10942 7644
rect 10998 7642 11022 7644
rect 11078 7642 11102 7644
rect 11158 7642 11164 7644
rect 10918 7590 10920 7642
rect 11100 7590 11102 7642
rect 10856 7588 10862 7590
rect 10918 7588 10942 7590
rect 10998 7588 11022 7590
rect 11078 7588 11102 7590
rect 11158 7588 11164 7590
rect 10856 7579 11164 7588
rect 11348 7546 11376 7754
rect 11336 7540 11388 7546
rect 11336 7482 11388 7488
rect 11152 7200 11204 7206
rect 11152 7142 11204 7148
rect 10784 6996 10836 7002
rect 10784 6938 10836 6944
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 9306 6012 9614 6021
rect 9306 6010 9312 6012
rect 9368 6010 9392 6012
rect 9448 6010 9472 6012
rect 9528 6010 9552 6012
rect 9608 6010 9614 6012
rect 9368 5958 9370 6010
rect 9550 5958 9552 6010
rect 9306 5956 9312 5958
rect 9368 5956 9392 5958
rect 9448 5956 9472 5958
rect 9528 5956 9552 5958
rect 9608 5956 9614 5958
rect 9306 5947 9614 5956
rect 10060 5710 10088 6734
rect 10048 5704 10100 5710
rect 10048 5646 10100 5652
rect 9220 5568 9272 5574
rect 9220 5510 9272 5516
rect 9128 5228 9180 5234
rect 9128 5170 9180 5176
rect 9036 4004 9088 4010
rect 9036 3946 9088 3952
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 9048 2990 9076 3946
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 9140 3194 9168 3878
rect 9128 3188 9180 3194
rect 9128 3130 9180 3136
rect 9036 2984 9088 2990
rect 9036 2926 9088 2932
rect 9036 2848 9088 2854
rect 9036 2790 9088 2796
rect 8668 1896 8720 1902
rect 8668 1838 8720 1844
rect 8680 1290 8708 1838
rect 8760 1420 8812 1426
rect 8760 1362 8812 1368
rect 8944 1420 8996 1426
rect 8944 1362 8996 1368
rect 8576 1284 8628 1290
rect 8576 1226 8628 1232
rect 8668 1284 8720 1290
rect 8668 1226 8720 1232
rect 7756 1116 8064 1125
rect 7756 1114 7762 1116
rect 7818 1114 7842 1116
rect 7898 1114 7922 1116
rect 7978 1114 8002 1116
rect 8058 1114 8064 1116
rect 7818 1062 7820 1114
rect 8000 1062 8002 1114
rect 7756 1060 7762 1062
rect 7818 1060 7842 1062
rect 7898 1060 7922 1062
rect 7978 1060 8002 1062
rect 8058 1060 8064 1062
rect 7756 1051 8064 1060
rect 8680 950 8708 1226
rect 8668 944 8720 950
rect 8668 886 8720 892
rect 8772 814 8800 1362
rect 8956 1018 8984 1362
rect 9048 1222 9076 2790
rect 9232 2774 9260 5510
rect 10060 5166 10088 5646
rect 10048 5160 10100 5166
rect 10048 5102 10100 5108
rect 9956 5024 10008 5030
rect 9956 4966 10008 4972
rect 9306 4924 9614 4933
rect 9306 4922 9312 4924
rect 9368 4922 9392 4924
rect 9448 4922 9472 4924
rect 9528 4922 9552 4924
rect 9608 4922 9614 4924
rect 9368 4870 9370 4922
rect 9550 4870 9552 4922
rect 9306 4868 9312 4870
rect 9368 4868 9392 4870
rect 9448 4868 9472 4870
rect 9528 4868 9552 4870
rect 9608 4868 9614 4870
rect 9306 4859 9614 4868
rect 9968 4690 9996 4966
rect 9956 4684 10008 4690
rect 9956 4626 10008 4632
rect 9306 3836 9614 3845
rect 9306 3834 9312 3836
rect 9368 3834 9392 3836
rect 9448 3834 9472 3836
rect 9528 3834 9552 3836
rect 9608 3834 9614 3836
rect 9368 3782 9370 3834
rect 9550 3782 9552 3834
rect 9306 3780 9312 3782
rect 9368 3780 9392 3782
rect 9448 3780 9472 3782
rect 9528 3780 9552 3782
rect 9608 3780 9614 3782
rect 9306 3771 9614 3780
rect 10796 3466 10824 6938
rect 11164 6798 11192 7142
rect 11716 7002 11744 11086
rect 12808 11076 12860 11082
rect 12808 11018 12860 11024
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 12452 10606 12480 10950
rect 12820 10810 12848 11018
rect 13452 11008 13504 11014
rect 13452 10950 13504 10956
rect 13464 10810 13492 10950
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 13452 10804 13504 10810
rect 13452 10746 13504 10752
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 12256 10464 12308 10470
rect 12256 10406 12308 10412
rect 12268 10266 12296 10406
rect 12406 10364 12714 10373
rect 12406 10362 12412 10364
rect 12468 10362 12492 10364
rect 12548 10362 12572 10364
rect 12628 10362 12652 10364
rect 12708 10362 12714 10364
rect 12468 10310 12470 10362
rect 12650 10310 12652 10362
rect 12406 10308 12412 10310
rect 12468 10308 12492 10310
rect 12548 10308 12572 10310
rect 12628 10308 12652 10310
rect 12708 10308 12714 10310
rect 12406 10299 12714 10308
rect 12256 10260 12308 10266
rect 12256 10202 12308 10208
rect 12820 10130 12848 10746
rect 13084 10600 13136 10606
rect 13084 10542 13136 10548
rect 13096 10266 13124 10542
rect 13084 10260 13136 10266
rect 13084 10202 13136 10208
rect 12900 10192 12952 10198
rect 12900 10134 12952 10140
rect 12808 10124 12860 10130
rect 12808 10066 12860 10072
rect 12348 9920 12400 9926
rect 12348 9862 12400 9868
rect 12360 9382 12388 9862
rect 11796 9376 11848 9382
rect 11796 9318 11848 9324
rect 12348 9376 12400 9382
rect 12348 9318 12400 9324
rect 11808 9110 11836 9318
rect 12406 9276 12714 9285
rect 12406 9274 12412 9276
rect 12468 9274 12492 9276
rect 12548 9274 12572 9276
rect 12628 9274 12652 9276
rect 12708 9274 12714 9276
rect 12468 9222 12470 9274
rect 12650 9222 12652 9274
rect 12406 9220 12412 9222
rect 12468 9220 12492 9222
rect 12548 9220 12572 9222
rect 12628 9220 12652 9222
rect 12708 9220 12714 9222
rect 12406 9211 12714 9220
rect 11796 9104 11848 9110
rect 11796 9046 11848 9052
rect 11704 6996 11756 7002
rect 11704 6938 11756 6944
rect 11808 6934 11836 9046
rect 12820 9042 12848 10066
rect 12912 9110 12940 10134
rect 12900 9104 12952 9110
rect 12900 9046 12952 9052
rect 12808 9036 12860 9042
rect 12808 8978 12860 8984
rect 12808 8900 12860 8906
rect 12808 8842 12860 8848
rect 12072 8832 12124 8838
rect 12072 8774 12124 8780
rect 12084 8498 12112 8774
rect 12072 8492 12124 8498
rect 12072 8434 12124 8440
rect 12406 8188 12714 8197
rect 12406 8186 12412 8188
rect 12468 8186 12492 8188
rect 12548 8186 12572 8188
rect 12628 8186 12652 8188
rect 12708 8186 12714 8188
rect 12468 8134 12470 8186
rect 12650 8134 12652 8186
rect 12406 8132 12412 8134
rect 12468 8132 12492 8134
rect 12548 8132 12572 8134
rect 12628 8132 12652 8134
rect 12708 8132 12714 8134
rect 12406 8123 12714 8132
rect 12820 8022 12848 8842
rect 12808 8016 12860 8022
rect 12808 7958 12860 7964
rect 12440 7948 12492 7954
rect 12440 7890 12492 7896
rect 12452 7342 12480 7890
rect 12912 7410 12940 9046
rect 13728 9036 13780 9042
rect 13728 8978 13780 8984
rect 13740 8498 13768 8978
rect 13728 8492 13780 8498
rect 13728 8434 13780 8440
rect 13740 7954 13768 8434
rect 13728 7948 13780 7954
rect 13728 7890 13780 7896
rect 13740 7546 13768 7890
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 12900 7404 12952 7410
rect 12900 7346 12952 7352
rect 12164 7336 12216 7342
rect 12164 7278 12216 7284
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 11796 6928 11848 6934
rect 11796 6870 11848 6876
rect 12072 6928 12124 6934
rect 12072 6870 12124 6876
rect 11152 6792 11204 6798
rect 11152 6734 11204 6740
rect 10856 6556 11164 6565
rect 10856 6554 10862 6556
rect 10918 6554 10942 6556
rect 10998 6554 11022 6556
rect 11078 6554 11102 6556
rect 11158 6554 11164 6556
rect 10918 6502 10920 6554
rect 11100 6502 11102 6554
rect 10856 6500 10862 6502
rect 10918 6500 10942 6502
rect 10998 6500 11022 6502
rect 11078 6500 11102 6502
rect 11158 6500 11164 6502
rect 10856 6491 11164 6500
rect 12084 6118 12112 6870
rect 12176 6798 12204 7278
rect 12406 7100 12714 7109
rect 12406 7098 12412 7100
rect 12468 7098 12492 7100
rect 12548 7098 12572 7100
rect 12628 7098 12652 7100
rect 12708 7098 12714 7100
rect 12468 7046 12470 7098
rect 12650 7046 12652 7098
rect 12406 7044 12412 7046
rect 12468 7044 12492 7046
rect 12548 7044 12572 7046
rect 12628 7044 12652 7046
rect 12708 7044 12714 7046
rect 12406 7035 12714 7044
rect 12164 6792 12216 6798
rect 12164 6734 12216 6740
rect 12176 6322 12204 6734
rect 12912 6730 12940 7346
rect 13452 6792 13504 6798
rect 13452 6734 13504 6740
rect 12900 6724 12952 6730
rect 12900 6666 12952 6672
rect 12164 6316 12216 6322
rect 12164 6258 12216 6264
rect 12912 6254 12940 6666
rect 13464 6458 13492 6734
rect 13452 6452 13504 6458
rect 13452 6394 13504 6400
rect 12900 6248 12952 6254
rect 12900 6190 12952 6196
rect 12072 6112 12124 6118
rect 12072 6054 12124 6060
rect 13268 6112 13320 6118
rect 13268 6054 13320 6060
rect 12084 5846 12112 6054
rect 12406 6012 12714 6021
rect 12406 6010 12412 6012
rect 12468 6010 12492 6012
rect 12548 6010 12572 6012
rect 12628 6010 12652 6012
rect 12708 6010 12714 6012
rect 12468 5958 12470 6010
rect 12650 5958 12652 6010
rect 12406 5956 12412 5958
rect 12468 5956 12492 5958
rect 12548 5956 12572 5958
rect 12628 5956 12652 5958
rect 12708 5956 12714 5958
rect 12406 5947 12714 5956
rect 12072 5840 12124 5846
rect 12072 5782 12124 5788
rect 11336 5704 11388 5710
rect 11336 5646 11388 5652
rect 10856 5468 11164 5477
rect 10856 5466 10862 5468
rect 10918 5466 10942 5468
rect 10998 5466 11022 5468
rect 11078 5466 11102 5468
rect 11158 5466 11164 5468
rect 10918 5414 10920 5466
rect 11100 5414 11102 5466
rect 10856 5412 10862 5414
rect 10918 5412 10942 5414
rect 10998 5412 11022 5414
rect 11078 5412 11102 5414
rect 11158 5412 11164 5414
rect 10856 5403 11164 5412
rect 11348 5370 11376 5646
rect 12084 5574 12112 5782
rect 13280 5710 13308 6054
rect 13832 5778 13860 12106
rect 13956 11996 14264 12005
rect 13956 11994 13962 11996
rect 14018 11994 14042 11996
rect 14098 11994 14122 11996
rect 14178 11994 14202 11996
rect 14258 11994 14264 11996
rect 14018 11942 14020 11994
rect 14200 11942 14202 11994
rect 13956 11940 13962 11942
rect 14018 11940 14042 11942
rect 14098 11940 14122 11942
rect 14178 11940 14202 11942
rect 14258 11940 14264 11942
rect 13956 11931 14264 11940
rect 14384 11558 14412 13330
rect 14660 12238 14688 13398
rect 14752 13394 14780 13670
rect 14740 13388 14792 13394
rect 14740 13330 14792 13336
rect 14844 13326 14872 13806
rect 14936 13394 14964 13806
rect 14924 13388 14976 13394
rect 14924 13330 14976 13336
rect 14832 13320 14884 13326
rect 14832 13262 14884 13268
rect 14648 12232 14700 12238
rect 14648 12174 14700 12180
rect 14936 12186 14964 13330
rect 15028 13326 15056 14214
rect 15016 13320 15068 13326
rect 15016 13262 15068 13268
rect 15028 12306 15056 13262
rect 15120 12374 15148 14334
rect 15304 14006 15332 15846
rect 15292 14000 15344 14006
rect 15292 13942 15344 13948
rect 15200 13932 15252 13938
rect 15200 13874 15252 13880
rect 15212 13530 15240 13874
rect 15200 13524 15252 13530
rect 15200 13466 15252 13472
rect 15304 12730 15332 13942
rect 15212 12714 15332 12730
rect 15200 12708 15332 12714
rect 15252 12702 15332 12708
rect 15200 12650 15252 12656
rect 15108 12368 15160 12374
rect 15108 12310 15160 12316
rect 15212 12306 15240 12650
rect 15292 12640 15344 12646
rect 15292 12582 15344 12588
rect 15304 12306 15332 12582
rect 15016 12300 15068 12306
rect 15016 12242 15068 12248
rect 15200 12300 15252 12306
rect 15200 12242 15252 12248
rect 15292 12300 15344 12306
rect 15292 12242 15344 12248
rect 14372 11552 14424 11558
rect 14372 11494 14424 11500
rect 13956 10908 14264 10917
rect 13956 10906 13962 10908
rect 14018 10906 14042 10908
rect 14098 10906 14122 10908
rect 14178 10906 14202 10908
rect 14258 10906 14264 10908
rect 14018 10854 14020 10906
rect 14200 10854 14202 10906
rect 13956 10852 13962 10854
rect 14018 10852 14042 10854
rect 14098 10852 14122 10854
rect 14178 10852 14202 10854
rect 14258 10852 14264 10854
rect 13956 10843 14264 10852
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 13956 9820 14264 9829
rect 13956 9818 13962 9820
rect 14018 9818 14042 9820
rect 14098 9818 14122 9820
rect 14178 9818 14202 9820
rect 14258 9818 14264 9820
rect 14018 9766 14020 9818
rect 14200 9766 14202 9818
rect 13956 9764 13962 9766
rect 14018 9764 14042 9766
rect 14098 9764 14122 9766
rect 14178 9764 14202 9766
rect 14258 9764 14264 9766
rect 13956 9755 14264 9764
rect 14292 9518 14320 10610
rect 14280 9512 14332 9518
rect 14280 9454 14332 9460
rect 14292 8906 14320 9454
rect 14280 8900 14332 8906
rect 14280 8842 14332 8848
rect 13956 8732 14264 8741
rect 13956 8730 13962 8732
rect 14018 8730 14042 8732
rect 14098 8730 14122 8732
rect 14178 8730 14202 8732
rect 14258 8730 14264 8732
rect 14018 8678 14020 8730
rect 14200 8678 14202 8730
rect 13956 8676 13962 8678
rect 14018 8676 14042 8678
rect 14098 8676 14122 8678
rect 14178 8676 14202 8678
rect 14258 8676 14264 8678
rect 13956 8667 14264 8676
rect 14292 8634 14320 8842
rect 14280 8628 14332 8634
rect 14280 8570 14332 8576
rect 13912 8288 13964 8294
rect 13912 8230 13964 8236
rect 13924 8090 13952 8230
rect 13912 8084 13964 8090
rect 13912 8026 13964 8032
rect 13956 7644 14264 7653
rect 13956 7642 13962 7644
rect 14018 7642 14042 7644
rect 14098 7642 14122 7644
rect 14178 7642 14202 7644
rect 14258 7642 14264 7644
rect 14018 7590 14020 7642
rect 14200 7590 14202 7642
rect 13956 7588 13962 7590
rect 14018 7588 14042 7590
rect 14098 7588 14122 7590
rect 14178 7588 14202 7590
rect 14258 7588 14264 7590
rect 13956 7579 14264 7588
rect 13956 6556 14264 6565
rect 13956 6554 13962 6556
rect 14018 6554 14042 6556
rect 14098 6554 14122 6556
rect 14178 6554 14202 6556
rect 14258 6554 14264 6556
rect 14018 6502 14020 6554
rect 14200 6502 14202 6554
rect 13956 6500 13962 6502
rect 14018 6500 14042 6502
rect 14098 6500 14122 6502
rect 14178 6500 14202 6502
rect 14258 6500 14264 6502
rect 13956 6491 14264 6500
rect 14292 6322 14320 8570
rect 14384 8022 14412 11494
rect 14464 10600 14516 10606
rect 14464 10542 14516 10548
rect 14476 10130 14504 10542
rect 14464 10124 14516 10130
rect 14464 10066 14516 10072
rect 14476 9450 14504 10066
rect 14660 9602 14688 12174
rect 14936 12158 15332 12186
rect 15108 11688 15160 11694
rect 15108 11630 15160 11636
rect 14832 11212 14884 11218
rect 14832 11154 14884 11160
rect 14844 10742 14872 11154
rect 15120 11082 15148 11630
rect 15200 11348 15252 11354
rect 15200 11290 15252 11296
rect 15212 11150 15240 11290
rect 15200 11144 15252 11150
rect 15200 11086 15252 11092
rect 15108 11076 15160 11082
rect 15108 11018 15160 11024
rect 14832 10736 14884 10742
rect 14832 10678 14884 10684
rect 14568 9574 14688 9602
rect 14464 9444 14516 9450
rect 14464 9386 14516 9392
rect 14476 9110 14504 9386
rect 14464 9104 14516 9110
rect 14464 9046 14516 9052
rect 14476 8838 14504 9046
rect 14464 8832 14516 8838
rect 14464 8774 14516 8780
rect 14568 8566 14596 9574
rect 14648 9512 14700 9518
rect 14648 9454 14700 9460
rect 14660 9178 14688 9454
rect 15120 9382 15148 11018
rect 15108 9376 15160 9382
rect 15108 9318 15160 9324
rect 14648 9172 14700 9178
rect 14648 9114 14700 9120
rect 14660 9042 14688 9114
rect 15120 9058 15148 9318
rect 14648 9036 14700 9042
rect 14648 8978 14700 8984
rect 15028 9030 15148 9058
rect 14556 8560 14608 8566
rect 14556 8502 14608 8508
rect 14568 8022 14596 8502
rect 14372 8016 14424 8022
rect 14372 7958 14424 7964
rect 14556 8016 14608 8022
rect 14556 7958 14608 7964
rect 14372 7404 14424 7410
rect 14372 7346 14424 7352
rect 14280 6316 14332 6322
rect 14280 6258 14332 6264
rect 13820 5772 13872 5778
rect 13820 5714 13872 5720
rect 13176 5704 13228 5710
rect 13176 5646 13228 5652
rect 13268 5704 13320 5710
rect 13268 5646 13320 5652
rect 11520 5568 11572 5574
rect 11520 5510 11572 5516
rect 12072 5568 12124 5574
rect 12072 5510 12124 5516
rect 12440 5568 12492 5574
rect 12440 5510 12492 5516
rect 12716 5568 12768 5574
rect 12716 5510 12768 5516
rect 11336 5364 11388 5370
rect 11336 5306 11388 5312
rect 11532 5098 11560 5510
rect 11520 5092 11572 5098
rect 11520 5034 11572 5040
rect 11244 4616 11296 4622
rect 11244 4558 11296 4564
rect 10856 4380 11164 4389
rect 10856 4378 10862 4380
rect 10918 4378 10942 4380
rect 10998 4378 11022 4380
rect 11078 4378 11102 4380
rect 11158 4378 11164 4380
rect 10918 4326 10920 4378
rect 11100 4326 11102 4378
rect 10856 4324 10862 4326
rect 10918 4324 10942 4326
rect 10998 4324 11022 4326
rect 11078 4324 11102 4326
rect 11158 4324 11164 4326
rect 10856 4315 11164 4324
rect 11256 4282 11284 4558
rect 11244 4276 11296 4282
rect 11244 4218 11296 4224
rect 11244 4072 11296 4078
rect 11244 4014 11296 4020
rect 11256 3602 11284 4014
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 11336 3596 11388 3602
rect 11336 3538 11388 3544
rect 10784 3460 10836 3466
rect 10784 3402 10836 3408
rect 10796 2990 10824 3402
rect 10856 3292 11164 3301
rect 10856 3290 10862 3292
rect 10918 3290 10942 3292
rect 10998 3290 11022 3292
rect 11078 3290 11102 3292
rect 11158 3290 11164 3292
rect 10918 3238 10920 3290
rect 11100 3238 11102 3290
rect 10856 3236 10862 3238
rect 10918 3236 10942 3238
rect 10998 3236 11022 3238
rect 11078 3236 11102 3238
rect 11158 3236 11164 3238
rect 10856 3227 11164 3236
rect 11256 3058 11284 3538
rect 11244 3052 11296 3058
rect 11244 2994 11296 3000
rect 11348 2990 11376 3538
rect 11532 3194 11560 5034
rect 11888 5024 11940 5030
rect 11888 4966 11940 4972
rect 11612 4480 11664 4486
rect 11612 4422 11664 4428
rect 11624 4078 11652 4422
rect 11612 4072 11664 4078
rect 11612 4014 11664 4020
rect 11612 3936 11664 3942
rect 11612 3878 11664 3884
rect 11520 3188 11572 3194
rect 11520 3130 11572 3136
rect 11428 3052 11480 3058
rect 11428 2994 11480 3000
rect 10784 2984 10836 2990
rect 10784 2926 10836 2932
rect 11336 2984 11388 2990
rect 11336 2926 11388 2932
rect 9140 2746 9260 2774
rect 9306 2748 9614 2757
rect 9306 2746 9312 2748
rect 9368 2746 9392 2748
rect 9448 2746 9472 2748
rect 9528 2746 9552 2748
rect 9608 2746 9614 2748
rect 9140 1834 9168 2746
rect 9368 2694 9370 2746
rect 9550 2694 9552 2746
rect 9306 2692 9312 2694
rect 9368 2692 9392 2694
rect 9448 2692 9472 2694
rect 9528 2692 9552 2694
rect 9608 2692 9614 2694
rect 9306 2683 9614 2692
rect 10856 2204 11164 2213
rect 10856 2202 10862 2204
rect 10918 2202 10942 2204
rect 10998 2202 11022 2204
rect 11078 2202 11102 2204
rect 11158 2202 11164 2204
rect 10918 2150 10920 2202
rect 11100 2150 11102 2202
rect 10856 2148 10862 2150
rect 10918 2148 10942 2150
rect 10998 2148 11022 2150
rect 11078 2148 11102 2150
rect 11158 2148 11164 2150
rect 10856 2139 11164 2148
rect 9128 1828 9180 1834
rect 9128 1770 9180 1776
rect 9140 1562 9168 1770
rect 9306 1660 9614 1669
rect 9306 1658 9312 1660
rect 9368 1658 9392 1660
rect 9448 1658 9472 1660
rect 9528 1658 9552 1660
rect 9608 1658 9614 1660
rect 9368 1606 9370 1658
rect 9550 1606 9552 1658
rect 9306 1604 9312 1606
rect 9368 1604 9392 1606
rect 9448 1604 9472 1606
rect 9528 1604 9552 1606
rect 9608 1604 9614 1606
rect 9306 1595 9614 1604
rect 9128 1556 9180 1562
rect 9128 1498 9180 1504
rect 9588 1556 9640 1562
rect 9588 1498 9640 1504
rect 9036 1216 9088 1222
rect 9036 1158 9088 1164
rect 8944 1012 8996 1018
rect 8944 954 8996 960
rect 9140 950 9168 1498
rect 9128 944 9180 950
rect 9128 886 9180 892
rect 9600 814 9628 1498
rect 11440 1426 11468 2994
rect 11520 2848 11572 2854
rect 11520 2790 11572 2796
rect 11532 1766 11560 2790
rect 11624 2106 11652 3878
rect 11796 3188 11848 3194
rect 11796 3130 11848 3136
rect 11612 2100 11664 2106
rect 11612 2042 11664 2048
rect 11520 1760 11572 1766
rect 11520 1702 11572 1708
rect 11532 1562 11560 1702
rect 11520 1556 11572 1562
rect 11520 1498 11572 1504
rect 11808 1426 11836 3130
rect 11900 2038 11928 4966
rect 12084 4758 12112 5510
rect 12452 5302 12480 5510
rect 12440 5296 12492 5302
rect 12440 5238 12492 5244
rect 12728 5234 12756 5510
rect 12716 5228 12768 5234
rect 12716 5170 12768 5176
rect 12728 5012 12756 5170
rect 12728 4984 12848 5012
rect 12406 4924 12714 4933
rect 12406 4922 12412 4924
rect 12468 4922 12492 4924
rect 12548 4922 12572 4924
rect 12628 4922 12652 4924
rect 12708 4922 12714 4924
rect 12468 4870 12470 4922
rect 12650 4870 12652 4922
rect 12406 4868 12412 4870
rect 12468 4868 12492 4870
rect 12548 4868 12572 4870
rect 12628 4868 12652 4870
rect 12708 4868 12714 4870
rect 12406 4859 12714 4868
rect 12072 4752 12124 4758
rect 12072 4694 12124 4700
rect 12256 4480 12308 4486
rect 12256 4422 12308 4428
rect 12268 3942 12296 4422
rect 12820 4214 12848 4984
rect 12808 4208 12860 4214
rect 12808 4150 12860 4156
rect 12808 4004 12860 4010
rect 12808 3946 12860 3952
rect 12256 3936 12308 3942
rect 12256 3878 12308 3884
rect 12268 3602 12296 3878
rect 12406 3836 12714 3845
rect 12406 3834 12412 3836
rect 12468 3834 12492 3836
rect 12548 3834 12572 3836
rect 12628 3834 12652 3836
rect 12708 3834 12714 3836
rect 12468 3782 12470 3834
rect 12650 3782 12652 3834
rect 12406 3780 12412 3782
rect 12468 3780 12492 3782
rect 12548 3780 12572 3782
rect 12628 3780 12652 3782
rect 12708 3780 12714 3782
rect 12406 3771 12714 3780
rect 12256 3596 12308 3602
rect 12256 3538 12308 3544
rect 12820 3194 12848 3946
rect 12808 3188 12860 3194
rect 12808 3130 12860 3136
rect 13188 3058 13216 5646
rect 13956 5468 14264 5477
rect 13956 5466 13962 5468
rect 14018 5466 14042 5468
rect 14098 5466 14122 5468
rect 14178 5466 14202 5468
rect 14258 5466 14264 5468
rect 14018 5414 14020 5466
rect 14200 5414 14202 5466
rect 13956 5412 13962 5414
rect 14018 5412 14042 5414
rect 14098 5412 14122 5414
rect 14178 5412 14202 5414
rect 14258 5412 14264 5414
rect 13956 5403 14264 5412
rect 13268 5228 13320 5234
rect 13268 5170 13320 5176
rect 13280 4758 13308 5170
rect 13544 5160 13596 5166
rect 13544 5102 13596 5108
rect 13556 4758 13584 5102
rect 13820 5092 13872 5098
rect 13820 5034 13872 5040
rect 13832 4826 13860 5034
rect 13820 4820 13872 4826
rect 13820 4762 13872 4768
rect 13268 4752 13320 4758
rect 13268 4694 13320 4700
rect 13544 4752 13596 4758
rect 13544 4694 13596 4700
rect 13820 4616 13872 4622
rect 13820 4558 13872 4564
rect 13832 3942 13860 4558
rect 13956 4380 14264 4389
rect 13956 4378 13962 4380
rect 14018 4378 14042 4380
rect 14098 4378 14122 4380
rect 14178 4378 14202 4380
rect 14258 4378 14264 4380
rect 14018 4326 14020 4378
rect 14200 4326 14202 4378
rect 13956 4324 13962 4326
rect 14018 4324 14042 4326
rect 14098 4324 14122 4326
rect 14178 4324 14202 4326
rect 14258 4324 14264 4326
rect 13956 4315 14264 4324
rect 14384 4078 14412 7346
rect 14464 7200 14516 7206
rect 14464 7142 14516 7148
rect 14476 7002 14504 7142
rect 14464 6996 14516 7002
rect 14464 6938 14516 6944
rect 14568 6458 14596 7958
rect 15028 7886 15056 9030
rect 15108 8900 15160 8906
rect 15108 8842 15160 8848
rect 15120 8090 15148 8842
rect 15108 8084 15160 8090
rect 15108 8026 15160 8032
rect 15016 7880 15068 7886
rect 15016 7822 15068 7828
rect 15028 6934 15056 7822
rect 15212 7274 15240 11086
rect 15304 8362 15332 12158
rect 15396 11898 15424 19230
rect 15580 19122 15608 19230
rect 15658 19200 15714 20000
rect 18510 19200 18566 20000
rect 15672 19122 15700 19200
rect 15580 19094 15700 19122
rect 18418 18592 18474 18601
rect 17056 18524 17364 18533
rect 18418 18527 18474 18536
rect 17056 18522 17062 18524
rect 17118 18522 17142 18524
rect 17198 18522 17222 18524
rect 17278 18522 17302 18524
rect 17358 18522 17364 18524
rect 17118 18470 17120 18522
rect 17300 18470 17302 18522
rect 17056 18468 17062 18470
rect 17118 18468 17142 18470
rect 17198 18468 17222 18470
rect 17278 18468 17302 18470
rect 17358 18468 17364 18470
rect 17056 18459 17364 18468
rect 18432 18426 18460 18527
rect 18420 18420 18472 18426
rect 18420 18362 18472 18368
rect 16028 18284 16080 18290
rect 16028 18226 16080 18232
rect 15506 17980 15814 17989
rect 15506 17978 15512 17980
rect 15568 17978 15592 17980
rect 15648 17978 15672 17980
rect 15728 17978 15752 17980
rect 15808 17978 15814 17980
rect 15568 17926 15570 17978
rect 15750 17926 15752 17978
rect 15506 17924 15512 17926
rect 15568 17924 15592 17926
rect 15648 17924 15672 17926
rect 15728 17924 15752 17926
rect 15808 17924 15814 17926
rect 15506 17915 15814 17924
rect 15936 16992 15988 16998
rect 15936 16934 15988 16940
rect 15506 16892 15814 16901
rect 15506 16890 15512 16892
rect 15568 16890 15592 16892
rect 15648 16890 15672 16892
rect 15728 16890 15752 16892
rect 15808 16890 15814 16892
rect 15568 16838 15570 16890
rect 15750 16838 15752 16890
rect 15506 16836 15512 16838
rect 15568 16836 15592 16838
rect 15648 16836 15672 16838
rect 15728 16836 15752 16838
rect 15808 16836 15814 16838
rect 15506 16827 15814 16836
rect 15948 16574 15976 16934
rect 16040 16794 16068 18226
rect 18432 18222 18460 18362
rect 18420 18216 18472 18222
rect 18420 18158 18472 18164
rect 17500 17740 17552 17746
rect 17500 17682 17552 17688
rect 16948 17672 17000 17678
rect 16948 17614 17000 17620
rect 16856 17536 16908 17542
rect 16856 17478 16908 17484
rect 16868 17202 16896 17478
rect 16856 17196 16908 17202
rect 16856 17138 16908 17144
rect 16580 17060 16632 17066
rect 16580 17002 16632 17008
rect 16028 16788 16080 16794
rect 16028 16730 16080 16736
rect 15948 16546 16068 16574
rect 16040 16114 16068 16546
rect 16120 16244 16172 16250
rect 16120 16186 16172 16192
rect 16028 16108 16080 16114
rect 16028 16050 16080 16056
rect 15936 15904 15988 15910
rect 15936 15846 15988 15852
rect 15506 15804 15814 15813
rect 15506 15802 15512 15804
rect 15568 15802 15592 15804
rect 15648 15802 15672 15804
rect 15728 15802 15752 15804
rect 15808 15802 15814 15804
rect 15568 15750 15570 15802
rect 15750 15750 15752 15802
rect 15506 15748 15512 15750
rect 15568 15748 15592 15750
rect 15648 15748 15672 15750
rect 15728 15748 15752 15750
rect 15808 15748 15814 15750
rect 15506 15739 15814 15748
rect 15948 15638 15976 15846
rect 15936 15632 15988 15638
rect 15936 15574 15988 15580
rect 15844 15564 15896 15570
rect 15844 15506 15896 15512
rect 15856 15162 15884 15506
rect 15936 15496 15988 15502
rect 15936 15438 15988 15444
rect 15844 15156 15896 15162
rect 15844 15098 15896 15104
rect 15948 14822 15976 15438
rect 15936 14816 15988 14822
rect 15936 14758 15988 14764
rect 15506 14716 15814 14725
rect 15506 14714 15512 14716
rect 15568 14714 15592 14716
rect 15648 14714 15672 14716
rect 15728 14714 15752 14716
rect 15808 14714 15814 14716
rect 15568 14662 15570 14714
rect 15750 14662 15752 14714
rect 15506 14660 15512 14662
rect 15568 14660 15592 14662
rect 15648 14660 15672 14662
rect 15728 14660 15752 14662
rect 15808 14660 15814 14662
rect 15506 14651 15814 14660
rect 15764 14482 15976 14498
rect 15752 14476 15988 14482
rect 15804 14470 15936 14476
rect 15752 14418 15804 14424
rect 15936 14418 15988 14424
rect 16040 14414 16068 16050
rect 16132 16046 16160 16186
rect 16120 16040 16172 16046
rect 16120 15982 16172 15988
rect 16132 15026 16160 15982
rect 16304 15972 16356 15978
rect 16304 15914 16356 15920
rect 16316 15706 16344 15914
rect 16592 15706 16620 17002
rect 16960 16114 16988 17614
rect 17056 17436 17364 17445
rect 17056 17434 17062 17436
rect 17118 17434 17142 17436
rect 17198 17434 17222 17436
rect 17278 17434 17302 17436
rect 17358 17434 17364 17436
rect 17118 17382 17120 17434
rect 17300 17382 17302 17434
rect 17056 17380 17062 17382
rect 17118 17380 17142 17382
rect 17198 17380 17222 17382
rect 17278 17380 17302 17382
rect 17358 17380 17364 17382
rect 17056 17371 17364 17380
rect 17512 16794 17540 17682
rect 17684 17672 17736 17678
rect 17684 17614 17736 17620
rect 17868 17672 17920 17678
rect 17868 17614 17920 17620
rect 17696 17338 17724 17614
rect 17684 17332 17736 17338
rect 17684 17274 17736 17280
rect 17696 17082 17724 17274
rect 17604 17054 17724 17082
rect 17500 16788 17552 16794
rect 17500 16730 17552 16736
rect 17500 16652 17552 16658
rect 17500 16594 17552 16600
rect 17056 16348 17364 16357
rect 17056 16346 17062 16348
rect 17118 16346 17142 16348
rect 17198 16346 17222 16348
rect 17278 16346 17302 16348
rect 17358 16346 17364 16348
rect 17118 16294 17120 16346
rect 17300 16294 17302 16346
rect 17056 16292 17062 16294
rect 17118 16292 17142 16294
rect 17198 16292 17222 16294
rect 17278 16292 17302 16294
rect 17358 16292 17364 16294
rect 17056 16283 17364 16292
rect 16948 16108 17000 16114
rect 16948 16050 17000 16056
rect 16304 15700 16356 15706
rect 16304 15642 16356 15648
rect 16580 15700 16632 15706
rect 16580 15642 16632 15648
rect 16212 15564 16264 15570
rect 16212 15506 16264 15512
rect 16120 15020 16172 15026
rect 16120 14962 16172 14968
rect 16120 14816 16172 14822
rect 16120 14758 16172 14764
rect 16028 14408 16080 14414
rect 16028 14350 16080 14356
rect 15568 14340 15620 14346
rect 15568 14282 15620 14288
rect 15580 14006 15608 14282
rect 15568 14000 15620 14006
rect 15568 13942 15620 13948
rect 16040 13734 16068 14350
rect 16028 13728 16080 13734
rect 16028 13670 16080 13676
rect 15506 13628 15814 13637
rect 15506 13626 15512 13628
rect 15568 13626 15592 13628
rect 15648 13626 15672 13628
rect 15728 13626 15752 13628
rect 15808 13626 15814 13628
rect 15568 13574 15570 13626
rect 15750 13574 15752 13626
rect 15506 13572 15512 13574
rect 15568 13572 15592 13574
rect 15648 13572 15672 13574
rect 15728 13572 15752 13574
rect 15808 13572 15814 13574
rect 15506 13563 15814 13572
rect 16132 13410 16160 14758
rect 16224 14278 16252 15506
rect 16212 14272 16264 14278
rect 16212 14214 16264 14220
rect 16316 13870 16344 15642
rect 16960 15570 16988 16050
rect 16488 15564 16540 15570
rect 16948 15564 17000 15570
rect 16488 15506 16540 15512
rect 16868 15524 16948 15552
rect 16396 14816 16448 14822
rect 16396 14758 16448 14764
rect 16408 14618 16436 14758
rect 16396 14612 16448 14618
rect 16396 14554 16448 14560
rect 16500 14550 16528 15506
rect 16488 14544 16540 14550
rect 16488 14486 16540 14492
rect 16868 14414 16896 15524
rect 16948 15506 17000 15512
rect 17408 15564 17460 15570
rect 17408 15506 17460 15512
rect 16948 15360 17000 15366
rect 16948 15302 17000 15308
rect 16856 14408 16908 14414
rect 16856 14350 16908 14356
rect 16868 14278 16896 14350
rect 16856 14272 16908 14278
rect 16856 14214 16908 14220
rect 16960 13938 16988 15302
rect 17056 15260 17364 15269
rect 17056 15258 17062 15260
rect 17118 15258 17142 15260
rect 17198 15258 17222 15260
rect 17278 15258 17302 15260
rect 17358 15258 17364 15260
rect 17118 15206 17120 15258
rect 17300 15206 17302 15258
rect 17056 15204 17062 15206
rect 17118 15204 17142 15206
rect 17198 15204 17222 15206
rect 17278 15204 17302 15206
rect 17358 15204 17364 15206
rect 17056 15195 17364 15204
rect 17420 14822 17448 15506
rect 17512 15366 17540 16594
rect 17604 16046 17632 17054
rect 17684 16584 17736 16590
rect 17684 16526 17736 16532
rect 17776 16584 17828 16590
rect 17776 16526 17828 16532
rect 17696 16182 17724 16526
rect 17788 16250 17816 16526
rect 17776 16244 17828 16250
rect 17776 16186 17828 16192
rect 17684 16176 17736 16182
rect 17684 16118 17736 16124
rect 17592 16040 17644 16046
rect 17592 15982 17644 15988
rect 17500 15360 17552 15366
rect 17500 15302 17552 15308
rect 17604 14958 17632 15982
rect 17788 15706 17816 16186
rect 17880 15978 17908 17614
rect 18420 16652 18472 16658
rect 18420 16594 18472 16600
rect 18052 16516 18104 16522
rect 18052 16458 18104 16464
rect 17868 15972 17920 15978
rect 17868 15914 17920 15920
rect 17776 15700 17828 15706
rect 17776 15642 17828 15648
rect 17592 14952 17644 14958
rect 17592 14894 17644 14900
rect 17132 14816 17184 14822
rect 17132 14758 17184 14764
rect 17408 14816 17460 14822
rect 17408 14758 17460 14764
rect 17144 14346 17172 14758
rect 17408 14408 17460 14414
rect 17408 14350 17460 14356
rect 17132 14340 17184 14346
rect 17132 14282 17184 14288
rect 17056 14172 17364 14181
rect 17056 14170 17062 14172
rect 17118 14170 17142 14172
rect 17198 14170 17222 14172
rect 17278 14170 17302 14172
rect 17358 14170 17364 14172
rect 17118 14118 17120 14170
rect 17300 14118 17302 14170
rect 17056 14116 17062 14118
rect 17118 14116 17142 14118
rect 17198 14116 17222 14118
rect 17278 14116 17302 14118
rect 17358 14116 17364 14118
rect 17056 14107 17364 14116
rect 16948 13932 17000 13938
rect 16948 13874 17000 13880
rect 17420 13870 17448 14350
rect 17604 14278 17632 14894
rect 17880 14482 17908 15914
rect 17960 14884 18012 14890
rect 17960 14826 18012 14832
rect 17972 14482 18000 14826
rect 17868 14476 17920 14482
rect 17868 14418 17920 14424
rect 17960 14476 18012 14482
rect 17960 14418 18012 14424
rect 17592 14272 17644 14278
rect 17592 14214 17644 14220
rect 16304 13864 16356 13870
rect 16304 13806 16356 13812
rect 17408 13864 17460 13870
rect 17408 13806 17460 13812
rect 16212 13796 16264 13802
rect 16212 13738 16264 13744
rect 16040 13382 16160 13410
rect 16224 13394 16252 13738
rect 16856 13728 16908 13734
rect 16856 13670 16908 13676
rect 16212 13388 16264 13394
rect 15506 12540 15814 12549
rect 15506 12538 15512 12540
rect 15568 12538 15592 12540
rect 15648 12538 15672 12540
rect 15728 12538 15752 12540
rect 15808 12538 15814 12540
rect 15568 12486 15570 12538
rect 15750 12486 15752 12538
rect 15506 12484 15512 12486
rect 15568 12484 15592 12486
rect 15648 12484 15672 12486
rect 15728 12484 15752 12486
rect 15808 12484 15814 12486
rect 15506 12475 15814 12484
rect 15384 11892 15436 11898
rect 15384 11834 15436 11840
rect 15506 11452 15814 11461
rect 15506 11450 15512 11452
rect 15568 11450 15592 11452
rect 15648 11450 15672 11452
rect 15728 11450 15752 11452
rect 15808 11450 15814 11452
rect 15568 11398 15570 11450
rect 15750 11398 15752 11450
rect 15506 11396 15512 11398
rect 15568 11396 15592 11398
rect 15648 11396 15672 11398
rect 15728 11396 15752 11398
rect 15808 11396 15814 11398
rect 15506 11387 15814 11396
rect 16040 11354 16068 13382
rect 16212 13330 16264 13336
rect 16304 13320 16356 13326
rect 16304 13262 16356 13268
rect 16212 13184 16264 13190
rect 16212 13126 16264 13132
rect 16120 12776 16172 12782
rect 16120 12718 16172 12724
rect 16132 11762 16160 12718
rect 16224 12646 16252 13126
rect 16212 12640 16264 12646
rect 16212 12582 16264 12588
rect 16120 11756 16172 11762
rect 16120 11698 16172 11704
rect 16028 11348 16080 11354
rect 16028 11290 16080 11296
rect 15936 11076 15988 11082
rect 15936 11018 15988 11024
rect 15948 10810 15976 11018
rect 15936 10804 15988 10810
rect 15936 10746 15988 10752
rect 15506 10364 15814 10373
rect 15506 10362 15512 10364
rect 15568 10362 15592 10364
rect 15648 10362 15672 10364
rect 15728 10362 15752 10364
rect 15808 10362 15814 10364
rect 15568 10310 15570 10362
rect 15750 10310 15752 10362
rect 15506 10308 15512 10310
rect 15568 10308 15592 10310
rect 15648 10308 15672 10310
rect 15728 10308 15752 10310
rect 15808 10308 15814 10310
rect 15506 10299 15814 10308
rect 15506 9276 15814 9285
rect 15506 9274 15512 9276
rect 15568 9274 15592 9276
rect 15648 9274 15672 9276
rect 15728 9274 15752 9276
rect 15808 9274 15814 9276
rect 15568 9222 15570 9274
rect 15750 9222 15752 9274
rect 15506 9220 15512 9222
rect 15568 9220 15592 9222
rect 15648 9220 15672 9222
rect 15728 9220 15752 9222
rect 15808 9220 15814 9222
rect 15506 9211 15814 9220
rect 15568 8832 15620 8838
rect 15568 8774 15620 8780
rect 15580 8634 15608 8774
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 15292 8356 15344 8362
rect 15292 8298 15344 8304
rect 15304 7342 15332 8298
rect 15506 8188 15814 8197
rect 15506 8186 15512 8188
rect 15568 8186 15592 8188
rect 15648 8186 15672 8188
rect 15728 8186 15752 8188
rect 15808 8186 15814 8188
rect 15568 8134 15570 8186
rect 15750 8134 15752 8186
rect 15506 8132 15512 8134
rect 15568 8132 15592 8134
rect 15648 8132 15672 8134
rect 15728 8132 15752 8134
rect 15808 8132 15814 8134
rect 15506 8123 15814 8132
rect 15384 7404 15436 7410
rect 15384 7346 15436 7352
rect 15292 7336 15344 7342
rect 15292 7278 15344 7284
rect 15200 7268 15252 7274
rect 15200 7210 15252 7216
rect 15212 7002 15240 7210
rect 15200 6996 15252 7002
rect 15200 6938 15252 6944
rect 15016 6928 15068 6934
rect 15304 6882 15332 7278
rect 15016 6870 15068 6876
rect 15108 6860 15160 6866
rect 15108 6802 15160 6808
rect 15212 6854 15332 6882
rect 15396 6866 15424 7346
rect 15506 7100 15814 7109
rect 15506 7098 15512 7100
rect 15568 7098 15592 7100
rect 15648 7098 15672 7100
rect 15728 7098 15752 7100
rect 15808 7098 15814 7100
rect 15568 7046 15570 7098
rect 15750 7046 15752 7098
rect 15506 7044 15512 7046
rect 15568 7044 15592 7046
rect 15648 7044 15672 7046
rect 15728 7044 15752 7046
rect 15808 7044 15814 7046
rect 15506 7035 15814 7044
rect 15384 6860 15436 6866
rect 15120 6458 15148 6802
rect 15212 6798 15240 6854
rect 15384 6802 15436 6808
rect 15200 6792 15252 6798
rect 15200 6734 15252 6740
rect 14556 6452 14608 6458
rect 14556 6394 14608 6400
rect 15108 6452 15160 6458
rect 15108 6394 15160 6400
rect 14568 6118 14596 6394
rect 14556 6112 14608 6118
rect 14556 6054 14608 6060
rect 14372 4072 14424 4078
rect 14372 4014 14424 4020
rect 14188 4004 14240 4010
rect 14188 3946 14240 3952
rect 13820 3936 13872 3942
rect 13820 3878 13872 3884
rect 14200 3738 14228 3946
rect 14568 3738 14596 6054
rect 15212 5846 15240 6734
rect 15506 6012 15814 6021
rect 15506 6010 15512 6012
rect 15568 6010 15592 6012
rect 15648 6010 15672 6012
rect 15728 6010 15752 6012
rect 15808 6010 15814 6012
rect 15568 5958 15570 6010
rect 15750 5958 15752 6010
rect 15506 5956 15512 5958
rect 15568 5956 15592 5958
rect 15648 5956 15672 5958
rect 15728 5956 15752 5958
rect 15808 5956 15814 5958
rect 15506 5947 15814 5956
rect 15200 5840 15252 5846
rect 15200 5782 15252 5788
rect 14924 5636 14976 5642
rect 14924 5578 14976 5584
rect 14936 4690 14964 5578
rect 15212 5556 15240 5782
rect 15660 5772 15712 5778
rect 15660 5714 15712 5720
rect 15844 5772 15896 5778
rect 15844 5714 15896 5720
rect 15120 5528 15240 5556
rect 14924 4684 14976 4690
rect 14924 4626 14976 4632
rect 14740 4616 14792 4622
rect 14740 4558 14792 4564
rect 14752 4282 14780 4558
rect 14740 4276 14792 4282
rect 14740 4218 14792 4224
rect 14832 4140 14884 4146
rect 14832 4082 14884 4088
rect 14188 3732 14240 3738
rect 14188 3674 14240 3680
rect 14556 3732 14608 3738
rect 14556 3674 14608 3680
rect 14372 3664 14424 3670
rect 14372 3606 14424 3612
rect 13956 3292 14264 3301
rect 13956 3290 13962 3292
rect 14018 3290 14042 3292
rect 14098 3290 14122 3292
rect 14178 3290 14202 3292
rect 14258 3290 14264 3292
rect 14018 3238 14020 3290
rect 14200 3238 14202 3290
rect 13956 3236 13962 3238
rect 14018 3236 14042 3238
rect 14098 3236 14122 3238
rect 14178 3236 14202 3238
rect 14258 3236 14264 3238
rect 13956 3227 14264 3236
rect 12808 3052 12860 3058
rect 12808 2994 12860 3000
rect 13176 3052 13228 3058
rect 13176 2994 13228 3000
rect 12406 2748 12714 2757
rect 12406 2746 12412 2748
rect 12468 2746 12492 2748
rect 12548 2746 12572 2748
rect 12628 2746 12652 2748
rect 12708 2746 12714 2748
rect 12468 2694 12470 2746
rect 12650 2694 12652 2746
rect 12406 2692 12412 2694
rect 12468 2692 12492 2694
rect 12548 2692 12572 2694
rect 12628 2692 12652 2694
rect 12708 2692 12714 2694
rect 12406 2683 12714 2692
rect 11888 2032 11940 2038
rect 12820 1986 12848 2994
rect 13176 2848 13228 2854
rect 13176 2790 13228 2796
rect 13728 2848 13780 2854
rect 13728 2790 13780 2796
rect 11888 1974 11940 1980
rect 12544 1970 12848 1986
rect 12532 1964 12848 1970
rect 12584 1958 12716 1964
rect 12532 1906 12584 1912
rect 12768 1958 12848 1964
rect 12716 1906 12768 1912
rect 12808 1760 12860 1766
rect 12808 1702 12860 1708
rect 12406 1660 12714 1669
rect 12406 1658 12412 1660
rect 12468 1658 12492 1660
rect 12548 1658 12572 1660
rect 12628 1658 12652 1660
rect 12708 1658 12714 1660
rect 12468 1606 12470 1658
rect 12650 1606 12652 1658
rect 12406 1604 12412 1606
rect 12468 1604 12492 1606
rect 12548 1604 12572 1606
rect 12628 1604 12652 1606
rect 12708 1604 12714 1606
rect 12406 1595 12714 1604
rect 11428 1420 11480 1426
rect 11428 1362 11480 1368
rect 11796 1420 11848 1426
rect 11796 1362 11848 1368
rect 12820 1290 12848 1702
rect 13188 1562 13216 2790
rect 13740 2514 13768 2790
rect 14384 2650 14412 3606
rect 14464 3596 14516 3602
rect 14464 3538 14516 3544
rect 14372 2644 14424 2650
rect 14372 2586 14424 2592
rect 14384 2514 14412 2586
rect 13728 2508 13780 2514
rect 13728 2450 13780 2456
rect 14372 2508 14424 2514
rect 14372 2450 14424 2456
rect 14384 2378 14412 2450
rect 14476 2446 14504 3538
rect 14844 3194 14872 4082
rect 15120 3602 15148 5528
rect 15672 5370 15700 5714
rect 15660 5364 15712 5370
rect 15660 5306 15712 5312
rect 15856 5098 15884 5714
rect 15948 5642 15976 10746
rect 16132 10674 16160 11698
rect 16120 10668 16172 10674
rect 16120 10610 16172 10616
rect 16224 10470 16252 12582
rect 16028 10464 16080 10470
rect 16028 10406 16080 10412
rect 16212 10464 16264 10470
rect 16212 10406 16264 10412
rect 16040 9926 16068 10406
rect 16028 9920 16080 9926
rect 16028 9862 16080 9868
rect 16316 9194 16344 13262
rect 16868 12850 16896 13670
rect 17056 13084 17364 13093
rect 17056 13082 17062 13084
rect 17118 13082 17142 13084
rect 17198 13082 17222 13084
rect 17278 13082 17302 13084
rect 17358 13082 17364 13084
rect 17118 13030 17120 13082
rect 17300 13030 17302 13082
rect 17056 13028 17062 13030
rect 17118 13028 17142 13030
rect 17198 13028 17222 13030
rect 17278 13028 17302 13030
rect 17358 13028 17364 13030
rect 17056 13019 17364 13028
rect 17972 12986 18000 14418
rect 17960 12980 18012 12986
rect 17960 12922 18012 12928
rect 16856 12844 16908 12850
rect 16856 12786 16908 12792
rect 16856 12436 16908 12442
rect 16856 12378 16908 12384
rect 17960 12436 18012 12442
rect 17960 12378 18012 12384
rect 16580 12232 16632 12238
rect 16580 12174 16632 12180
rect 16488 11688 16540 11694
rect 16488 11630 16540 11636
rect 16500 11354 16528 11630
rect 16488 11348 16540 11354
rect 16488 11290 16540 11296
rect 16488 10532 16540 10538
rect 16488 10474 16540 10480
rect 16500 10266 16528 10474
rect 16488 10260 16540 10266
rect 16488 10202 16540 10208
rect 16592 9994 16620 12174
rect 16868 11626 16896 12378
rect 16948 12096 17000 12102
rect 16948 12038 17000 12044
rect 16856 11620 16908 11626
rect 16856 11562 16908 11568
rect 16672 11348 16724 11354
rect 16672 11290 16724 11296
rect 16684 10810 16712 11290
rect 16764 11280 16816 11286
rect 16764 11222 16816 11228
rect 16776 11014 16804 11222
rect 16764 11008 16816 11014
rect 16764 10950 16816 10956
rect 16672 10804 16724 10810
rect 16672 10746 16724 10752
rect 16960 10198 16988 12038
rect 17056 11996 17364 12005
rect 17056 11994 17062 11996
rect 17118 11994 17142 11996
rect 17198 11994 17222 11996
rect 17278 11994 17302 11996
rect 17358 11994 17364 11996
rect 17118 11942 17120 11994
rect 17300 11942 17302 11994
rect 17056 11940 17062 11942
rect 17118 11940 17142 11942
rect 17198 11940 17222 11942
rect 17278 11940 17302 11942
rect 17358 11940 17364 11942
rect 17056 11931 17364 11940
rect 17972 11762 18000 12378
rect 17960 11756 18012 11762
rect 17960 11698 18012 11704
rect 17316 11552 17368 11558
rect 17316 11494 17368 11500
rect 17328 11218 17356 11494
rect 18064 11354 18092 16458
rect 18432 16250 18460 16594
rect 18420 16244 18472 16250
rect 18420 16186 18472 16192
rect 18432 16153 18460 16186
rect 18418 16144 18474 16153
rect 18418 16079 18474 16088
rect 18236 14272 18288 14278
rect 18236 14214 18288 14220
rect 18144 14000 18196 14006
rect 18144 13942 18196 13948
rect 18052 11348 18104 11354
rect 18052 11290 18104 11296
rect 17316 11212 17368 11218
rect 17316 11154 17368 11160
rect 17500 11212 17552 11218
rect 17500 11154 17552 11160
rect 17056 10908 17364 10917
rect 17056 10906 17062 10908
rect 17118 10906 17142 10908
rect 17198 10906 17222 10908
rect 17278 10906 17302 10908
rect 17358 10906 17364 10908
rect 17118 10854 17120 10906
rect 17300 10854 17302 10906
rect 17056 10852 17062 10854
rect 17118 10852 17142 10854
rect 17198 10852 17222 10854
rect 17278 10852 17302 10854
rect 17358 10852 17364 10854
rect 17056 10843 17364 10852
rect 17512 10810 17540 11154
rect 17500 10804 17552 10810
rect 17500 10746 17552 10752
rect 17684 10804 17736 10810
rect 17684 10746 17736 10752
rect 16948 10192 17000 10198
rect 16948 10134 17000 10140
rect 17696 10130 17724 10746
rect 17316 10124 17368 10130
rect 17316 10066 17368 10072
rect 17684 10124 17736 10130
rect 17684 10066 17736 10072
rect 16580 9988 16632 9994
rect 16580 9930 16632 9936
rect 17328 9908 17356 10066
rect 17592 9988 17644 9994
rect 17592 9930 17644 9936
rect 17328 9880 17448 9908
rect 17056 9820 17364 9829
rect 17056 9818 17062 9820
rect 17118 9818 17142 9820
rect 17198 9818 17222 9820
rect 17278 9818 17302 9820
rect 17358 9818 17364 9820
rect 17118 9766 17120 9818
rect 17300 9766 17302 9818
rect 17056 9764 17062 9766
rect 17118 9764 17142 9766
rect 17198 9764 17222 9766
rect 17278 9764 17302 9766
rect 17358 9764 17364 9766
rect 17056 9755 17364 9764
rect 16224 9166 16344 9194
rect 17420 9178 17448 9880
rect 17408 9172 17460 9178
rect 16224 8498 16252 9166
rect 17408 9114 17460 9120
rect 17500 9104 17552 9110
rect 17500 9046 17552 9052
rect 16304 9036 16356 9042
rect 16304 8978 16356 8984
rect 16316 8566 16344 8978
rect 17056 8732 17364 8741
rect 17056 8730 17062 8732
rect 17118 8730 17142 8732
rect 17198 8730 17222 8732
rect 17278 8730 17302 8732
rect 17358 8730 17364 8732
rect 17118 8678 17120 8730
rect 17300 8678 17302 8730
rect 17056 8676 17062 8678
rect 17118 8676 17142 8678
rect 17198 8676 17222 8678
rect 17278 8676 17302 8678
rect 17358 8676 17364 8678
rect 17056 8667 17364 8676
rect 16304 8560 16356 8566
rect 16304 8502 16356 8508
rect 16212 8492 16264 8498
rect 16212 8434 16264 8440
rect 16396 8424 16448 8430
rect 16396 8366 16448 8372
rect 17224 8424 17276 8430
rect 17224 8366 17276 8372
rect 16408 7410 16436 8366
rect 16672 8356 16724 8362
rect 16672 8298 16724 8304
rect 16684 7954 16712 8298
rect 17236 7954 17264 8366
rect 17512 8090 17540 9046
rect 17500 8084 17552 8090
rect 17500 8026 17552 8032
rect 16672 7948 16724 7954
rect 16672 7890 16724 7896
rect 17224 7948 17276 7954
rect 17224 7890 17276 7896
rect 16684 7546 16712 7890
rect 17056 7644 17364 7653
rect 17056 7642 17062 7644
rect 17118 7642 17142 7644
rect 17198 7642 17222 7644
rect 17278 7642 17302 7644
rect 17358 7642 17364 7644
rect 17118 7590 17120 7642
rect 17300 7590 17302 7642
rect 17056 7588 17062 7590
rect 17118 7588 17142 7590
rect 17198 7588 17222 7590
rect 17278 7588 17302 7590
rect 17358 7588 17364 7590
rect 17056 7579 17364 7588
rect 16672 7540 16724 7546
rect 16672 7482 16724 7488
rect 16396 7404 16448 7410
rect 16396 7346 16448 7352
rect 16304 7268 16356 7274
rect 16304 7210 16356 7216
rect 16028 6180 16080 6186
rect 16028 6122 16080 6128
rect 15936 5636 15988 5642
rect 15936 5578 15988 5584
rect 16040 5166 16068 6122
rect 16316 5794 16344 7210
rect 16408 6322 16436 7346
rect 16764 6656 16816 6662
rect 16764 6598 16816 6604
rect 16396 6316 16448 6322
rect 16396 6258 16448 6264
rect 16224 5778 16344 5794
rect 16224 5772 16356 5778
rect 16224 5766 16304 5772
rect 16028 5160 16080 5166
rect 16028 5102 16080 5108
rect 15844 5092 15896 5098
rect 15844 5034 15896 5040
rect 15506 4924 15814 4933
rect 15506 4922 15512 4924
rect 15568 4922 15592 4924
rect 15648 4922 15672 4924
rect 15728 4922 15752 4924
rect 15808 4922 15814 4924
rect 15568 4870 15570 4922
rect 15750 4870 15752 4922
rect 15506 4868 15512 4870
rect 15568 4868 15592 4870
rect 15648 4868 15672 4870
rect 15728 4868 15752 4870
rect 15808 4868 15814 4870
rect 15506 4859 15814 4868
rect 15384 4684 15436 4690
rect 15384 4626 15436 4632
rect 15108 3596 15160 3602
rect 15108 3538 15160 3544
rect 14832 3188 14884 3194
rect 14832 3130 14884 3136
rect 15120 2990 15148 3538
rect 15108 2984 15160 2990
rect 15108 2926 15160 2932
rect 15120 2582 15148 2926
rect 15200 2848 15252 2854
rect 15200 2790 15252 2796
rect 15212 2650 15240 2790
rect 15396 2650 15424 4626
rect 15506 3836 15814 3845
rect 15506 3834 15512 3836
rect 15568 3834 15592 3836
rect 15648 3834 15672 3836
rect 15728 3834 15752 3836
rect 15808 3834 15814 3836
rect 15568 3782 15570 3834
rect 15750 3782 15752 3834
rect 15506 3780 15512 3782
rect 15568 3780 15592 3782
rect 15648 3780 15672 3782
rect 15728 3780 15752 3782
rect 15808 3780 15814 3782
rect 15506 3771 15814 3780
rect 15506 2748 15814 2757
rect 15506 2746 15512 2748
rect 15568 2746 15592 2748
rect 15648 2746 15672 2748
rect 15728 2746 15752 2748
rect 15808 2746 15814 2748
rect 15568 2694 15570 2746
rect 15750 2694 15752 2746
rect 15506 2692 15512 2694
rect 15568 2692 15592 2694
rect 15648 2692 15672 2694
rect 15728 2692 15752 2694
rect 15808 2692 15814 2694
rect 15506 2683 15814 2692
rect 15200 2644 15252 2650
rect 15200 2586 15252 2592
rect 15384 2644 15436 2650
rect 15384 2586 15436 2592
rect 15108 2576 15160 2582
rect 15108 2518 15160 2524
rect 14464 2440 14516 2446
rect 14464 2382 14516 2388
rect 13268 2372 13320 2378
rect 13268 2314 13320 2320
rect 14372 2372 14424 2378
rect 14372 2314 14424 2320
rect 13280 1970 13308 2314
rect 13728 2304 13780 2310
rect 13728 2246 13780 2252
rect 13740 2038 13768 2246
rect 13956 2204 14264 2213
rect 13956 2202 13962 2204
rect 14018 2202 14042 2204
rect 14098 2202 14122 2204
rect 14178 2202 14202 2204
rect 14258 2202 14264 2204
rect 14018 2150 14020 2202
rect 14200 2150 14202 2202
rect 13956 2148 13962 2150
rect 14018 2148 14042 2150
rect 14098 2148 14122 2150
rect 14178 2148 14202 2150
rect 14258 2148 14264 2150
rect 13956 2139 14264 2148
rect 13728 2032 13780 2038
rect 13728 1974 13780 1980
rect 13268 1964 13320 1970
rect 13268 1906 13320 1912
rect 14004 1964 14056 1970
rect 14004 1906 14056 1912
rect 13728 1896 13780 1902
rect 13728 1838 13780 1844
rect 13176 1556 13228 1562
rect 13176 1498 13228 1504
rect 13740 1358 13768 1838
rect 14016 1426 14044 1906
rect 14384 1562 14412 2314
rect 14476 1970 14504 2382
rect 14464 1964 14516 1970
rect 14464 1906 14516 1912
rect 15396 1902 15424 2586
rect 15568 2440 15620 2446
rect 15568 2382 15620 2388
rect 15580 1902 15608 2382
rect 15108 1896 15160 1902
rect 15108 1838 15160 1844
rect 15384 1896 15436 1902
rect 15384 1838 15436 1844
rect 15568 1896 15620 1902
rect 15568 1838 15620 1844
rect 14372 1556 14424 1562
rect 14372 1498 14424 1504
rect 15120 1426 15148 1838
rect 15396 1494 15424 1838
rect 15506 1660 15814 1669
rect 15506 1658 15512 1660
rect 15568 1658 15592 1660
rect 15648 1658 15672 1660
rect 15728 1658 15752 1660
rect 15808 1658 15814 1660
rect 15568 1606 15570 1658
rect 15750 1606 15752 1658
rect 15506 1604 15512 1606
rect 15568 1604 15592 1606
rect 15648 1604 15672 1606
rect 15728 1604 15752 1606
rect 15808 1604 15814 1606
rect 15506 1595 15814 1604
rect 15384 1488 15436 1494
rect 15384 1430 15436 1436
rect 15856 1426 15884 5034
rect 16040 4826 16068 5102
rect 16028 4820 16080 4826
rect 16028 4762 16080 4768
rect 16224 4078 16252 5766
rect 16304 5714 16356 5720
rect 16304 5636 16356 5642
rect 16304 5578 16356 5584
rect 16212 4072 16264 4078
rect 16212 4014 16264 4020
rect 16120 3936 16172 3942
rect 16120 3878 16172 3884
rect 16132 3602 16160 3878
rect 16120 3596 16172 3602
rect 16120 3538 16172 3544
rect 16224 3466 16252 4014
rect 16316 3738 16344 5578
rect 16408 5234 16436 6258
rect 16488 6248 16540 6254
rect 16488 6190 16540 6196
rect 16500 5914 16528 6190
rect 16488 5908 16540 5914
rect 16488 5850 16540 5856
rect 16776 5794 16804 6598
rect 17056 6556 17364 6565
rect 17056 6554 17062 6556
rect 17118 6554 17142 6556
rect 17198 6554 17222 6556
rect 17278 6554 17302 6556
rect 17358 6554 17364 6556
rect 17118 6502 17120 6554
rect 17300 6502 17302 6554
rect 17056 6500 17062 6502
rect 17118 6500 17142 6502
rect 17198 6500 17222 6502
rect 17278 6500 17302 6502
rect 17358 6500 17364 6502
rect 17056 6491 17364 6500
rect 17604 6338 17632 9930
rect 17960 9036 18012 9042
rect 17960 8978 18012 8984
rect 17972 8634 18000 8978
rect 17960 8628 18012 8634
rect 17960 8570 18012 8576
rect 17420 6310 17632 6338
rect 16948 6112 17000 6118
rect 16948 6054 17000 6060
rect 16960 5846 16988 6054
rect 16500 5778 16804 5794
rect 16948 5840 17000 5846
rect 16948 5782 17000 5788
rect 17420 5778 17448 6310
rect 17500 6180 17552 6186
rect 17500 6122 17552 6128
rect 17960 6180 18012 6186
rect 17960 6122 18012 6128
rect 16500 5772 16816 5778
rect 16500 5766 16764 5772
rect 16396 5228 16448 5234
rect 16396 5170 16448 5176
rect 16408 4758 16436 5170
rect 16396 4752 16448 4758
rect 16396 4694 16448 4700
rect 16500 4146 16528 5766
rect 16764 5714 16816 5720
rect 17408 5772 17460 5778
rect 17408 5714 17460 5720
rect 17056 5468 17364 5477
rect 17056 5466 17062 5468
rect 17118 5466 17142 5468
rect 17198 5466 17222 5468
rect 17278 5466 17302 5468
rect 17358 5466 17364 5468
rect 17118 5414 17120 5466
rect 17300 5414 17302 5466
rect 17056 5412 17062 5414
rect 17118 5412 17142 5414
rect 17198 5412 17222 5414
rect 17278 5412 17302 5414
rect 17358 5412 17364 5414
rect 17056 5403 17364 5412
rect 16672 5092 16724 5098
rect 16672 5034 16724 5040
rect 16684 4146 16712 5034
rect 17056 4380 17364 4389
rect 17056 4378 17062 4380
rect 17118 4378 17142 4380
rect 17198 4378 17222 4380
rect 17278 4378 17302 4380
rect 17358 4378 17364 4380
rect 17118 4326 17120 4378
rect 17300 4326 17302 4378
rect 17056 4324 17062 4326
rect 17118 4324 17142 4326
rect 17198 4324 17222 4326
rect 17278 4324 17302 4326
rect 17358 4324 17364 4326
rect 17056 4315 17364 4324
rect 16856 4208 16908 4214
rect 16856 4150 16908 4156
rect 16488 4140 16540 4146
rect 16488 4082 16540 4088
rect 16672 4140 16724 4146
rect 16672 4082 16724 4088
rect 16304 3732 16356 3738
rect 16304 3674 16356 3680
rect 16500 3602 16528 4082
rect 16672 4004 16724 4010
rect 16672 3946 16724 3952
rect 16580 3936 16632 3942
rect 16580 3878 16632 3884
rect 16592 3738 16620 3878
rect 16580 3732 16632 3738
rect 16580 3674 16632 3680
rect 16488 3596 16540 3602
rect 16488 3538 16540 3544
rect 16212 3460 16264 3466
rect 16212 3402 16264 3408
rect 16224 2106 16252 3402
rect 16500 3058 16528 3538
rect 16488 3052 16540 3058
rect 16488 2994 16540 3000
rect 16304 2440 16356 2446
rect 16304 2382 16356 2388
rect 16212 2100 16264 2106
rect 16212 2042 16264 2048
rect 16224 1766 16252 2042
rect 16316 1970 16344 2382
rect 16684 2106 16712 3946
rect 16672 2100 16724 2106
rect 16672 2042 16724 2048
rect 16304 1964 16356 1970
rect 16304 1906 16356 1912
rect 16868 1902 16896 4150
rect 17420 4146 17448 5714
rect 17512 5166 17540 6122
rect 17972 5710 18000 6122
rect 17960 5704 18012 5710
rect 17960 5646 18012 5652
rect 17592 5364 17644 5370
rect 17592 5306 17644 5312
rect 17500 5160 17552 5166
rect 17500 5102 17552 5108
rect 17512 4826 17540 5102
rect 17500 4820 17552 4826
rect 17500 4762 17552 4768
rect 17604 4214 17632 5306
rect 17592 4208 17644 4214
rect 17592 4150 17644 4156
rect 17408 4140 17460 4146
rect 17408 4082 17460 4088
rect 17420 3942 17448 4082
rect 17500 4072 17552 4078
rect 17500 4014 17552 4020
rect 17408 3936 17460 3942
rect 17408 3878 17460 3884
rect 17420 3602 17448 3878
rect 17512 3738 17540 4014
rect 17500 3732 17552 3738
rect 17500 3674 17552 3680
rect 17408 3596 17460 3602
rect 17408 3538 17460 3544
rect 16948 3392 17000 3398
rect 16948 3334 17000 3340
rect 16960 3194 16988 3334
rect 17056 3292 17364 3301
rect 17056 3290 17062 3292
rect 17118 3290 17142 3292
rect 17198 3290 17222 3292
rect 17278 3290 17302 3292
rect 17358 3290 17364 3292
rect 17118 3238 17120 3290
rect 17300 3238 17302 3290
rect 17056 3236 17062 3238
rect 17118 3236 17142 3238
rect 17198 3236 17222 3238
rect 17278 3236 17302 3238
rect 17358 3236 17364 3238
rect 17056 3227 17364 3236
rect 16948 3188 17000 3194
rect 16948 3130 17000 3136
rect 17592 2916 17644 2922
rect 17592 2858 17644 2864
rect 17500 2848 17552 2854
rect 17500 2790 17552 2796
rect 17512 2650 17540 2790
rect 17604 2650 17632 2858
rect 17500 2644 17552 2650
rect 17500 2586 17552 2592
rect 17592 2644 17644 2650
rect 17592 2586 17644 2592
rect 17592 2508 17644 2514
rect 17592 2450 17644 2456
rect 17056 2204 17364 2213
rect 17056 2202 17062 2204
rect 17118 2202 17142 2204
rect 17198 2202 17222 2204
rect 17278 2202 17302 2204
rect 17358 2202 17364 2204
rect 17118 2150 17120 2202
rect 17300 2150 17302 2202
rect 17056 2148 17062 2150
rect 17118 2148 17142 2150
rect 17198 2148 17222 2150
rect 17278 2148 17302 2150
rect 17358 2148 17364 2150
rect 17056 2139 17364 2148
rect 16856 1896 16908 1902
rect 16856 1838 16908 1844
rect 16212 1760 16264 1766
rect 16212 1702 16264 1708
rect 16304 1760 16356 1766
rect 16304 1702 16356 1708
rect 16316 1562 16344 1702
rect 16304 1556 16356 1562
rect 16304 1498 16356 1504
rect 14004 1420 14056 1426
rect 14004 1362 14056 1368
rect 15108 1420 15160 1426
rect 15108 1362 15160 1368
rect 15844 1420 15896 1426
rect 15844 1362 15896 1368
rect 13728 1352 13780 1358
rect 13728 1294 13780 1300
rect 12808 1284 12860 1290
rect 12808 1226 12860 1232
rect 10856 1116 11164 1125
rect 10856 1114 10862 1116
rect 10918 1114 10942 1116
rect 10998 1114 11022 1116
rect 11078 1114 11102 1116
rect 11158 1114 11164 1116
rect 10918 1062 10920 1114
rect 11100 1062 11102 1114
rect 10856 1060 10862 1062
rect 10918 1060 10942 1062
rect 10998 1060 11022 1062
rect 11078 1060 11102 1062
rect 11158 1060 11164 1062
rect 10856 1051 11164 1060
rect 13956 1116 14264 1125
rect 13956 1114 13962 1116
rect 14018 1114 14042 1116
rect 14098 1114 14122 1116
rect 14178 1114 14202 1116
rect 14258 1114 14264 1116
rect 14018 1062 14020 1114
rect 14200 1062 14202 1114
rect 13956 1060 13962 1062
rect 14018 1060 14042 1062
rect 14098 1060 14122 1062
rect 14178 1060 14202 1062
rect 14258 1060 14264 1062
rect 13956 1051 14264 1060
rect 15856 950 15884 1362
rect 16868 1358 16896 1838
rect 17604 1562 17632 2450
rect 17972 2038 18000 5646
rect 18156 3738 18184 13942
rect 18248 13938 18276 14214
rect 18236 13932 18288 13938
rect 18236 13874 18288 13880
rect 18524 12442 18552 19200
rect 18606 17980 18914 17989
rect 18606 17978 18612 17980
rect 18668 17978 18692 17980
rect 18748 17978 18772 17980
rect 18828 17978 18852 17980
rect 18908 17978 18914 17980
rect 18668 17926 18670 17978
rect 18850 17926 18852 17978
rect 18606 17924 18612 17926
rect 18668 17924 18692 17926
rect 18748 17924 18772 17926
rect 18828 17924 18852 17926
rect 18908 17924 18914 17926
rect 18606 17915 18914 17924
rect 18606 16892 18914 16901
rect 18606 16890 18612 16892
rect 18668 16890 18692 16892
rect 18748 16890 18772 16892
rect 18828 16890 18852 16892
rect 18908 16890 18914 16892
rect 18668 16838 18670 16890
rect 18850 16838 18852 16890
rect 18606 16836 18612 16838
rect 18668 16836 18692 16838
rect 18748 16836 18772 16838
rect 18828 16836 18852 16838
rect 18908 16836 18914 16838
rect 18606 16827 18914 16836
rect 18606 15804 18914 15813
rect 18606 15802 18612 15804
rect 18668 15802 18692 15804
rect 18748 15802 18772 15804
rect 18828 15802 18852 15804
rect 18908 15802 18914 15804
rect 18668 15750 18670 15802
rect 18850 15750 18852 15802
rect 18606 15748 18612 15750
rect 18668 15748 18692 15750
rect 18748 15748 18772 15750
rect 18828 15748 18852 15750
rect 18908 15748 18914 15750
rect 18606 15739 18914 15748
rect 18606 14716 18914 14725
rect 18606 14714 18612 14716
rect 18668 14714 18692 14716
rect 18748 14714 18772 14716
rect 18828 14714 18852 14716
rect 18908 14714 18914 14716
rect 18668 14662 18670 14714
rect 18850 14662 18852 14714
rect 18606 14660 18612 14662
rect 18668 14660 18692 14662
rect 18748 14660 18772 14662
rect 18828 14660 18852 14662
rect 18908 14660 18914 14662
rect 18606 14651 18914 14660
rect 19064 13864 19116 13870
rect 19064 13806 19116 13812
rect 19076 13705 19104 13806
rect 19062 13696 19118 13705
rect 18606 13628 18914 13637
rect 19062 13631 19118 13640
rect 18606 13626 18612 13628
rect 18668 13626 18692 13628
rect 18748 13626 18772 13628
rect 18828 13626 18852 13628
rect 18908 13626 18914 13628
rect 18668 13574 18670 13626
rect 18850 13574 18852 13626
rect 18606 13572 18612 13574
rect 18668 13572 18692 13574
rect 18748 13572 18772 13574
rect 18828 13572 18852 13574
rect 18908 13572 18914 13574
rect 18606 13563 18914 13572
rect 18606 12540 18914 12549
rect 18606 12538 18612 12540
rect 18668 12538 18692 12540
rect 18748 12538 18772 12540
rect 18828 12538 18852 12540
rect 18908 12538 18914 12540
rect 18668 12486 18670 12538
rect 18850 12486 18852 12538
rect 18606 12484 18612 12486
rect 18668 12484 18692 12486
rect 18748 12484 18772 12486
rect 18828 12484 18852 12486
rect 18908 12484 18914 12486
rect 18606 12475 18914 12484
rect 18512 12436 18564 12442
rect 18512 12378 18564 12384
rect 18236 11892 18288 11898
rect 18236 11834 18288 11840
rect 18248 9178 18276 11834
rect 18606 11452 18914 11461
rect 18606 11450 18612 11452
rect 18668 11450 18692 11452
rect 18748 11450 18772 11452
rect 18828 11450 18852 11452
rect 18908 11450 18914 11452
rect 18668 11398 18670 11450
rect 18850 11398 18852 11450
rect 18606 11396 18612 11398
rect 18668 11396 18692 11398
rect 18748 11396 18772 11398
rect 18828 11396 18852 11398
rect 18908 11396 18914 11398
rect 18606 11387 18914 11396
rect 18418 11248 18474 11257
rect 18418 11183 18420 11192
rect 18472 11183 18474 11192
rect 18420 11154 18472 11160
rect 18606 10364 18914 10373
rect 18606 10362 18612 10364
rect 18668 10362 18692 10364
rect 18748 10362 18772 10364
rect 18828 10362 18852 10364
rect 18908 10362 18914 10364
rect 18668 10310 18670 10362
rect 18850 10310 18852 10362
rect 18606 10308 18612 10310
rect 18668 10308 18692 10310
rect 18748 10308 18772 10310
rect 18828 10308 18852 10310
rect 18908 10308 18914 10310
rect 18606 10299 18914 10308
rect 18606 9276 18914 9285
rect 18606 9274 18612 9276
rect 18668 9274 18692 9276
rect 18748 9274 18772 9276
rect 18828 9274 18852 9276
rect 18908 9274 18914 9276
rect 18668 9222 18670 9274
rect 18850 9222 18852 9274
rect 18606 9220 18612 9222
rect 18668 9220 18692 9222
rect 18748 9220 18772 9222
rect 18828 9220 18852 9222
rect 18908 9220 18914 9222
rect 18606 9211 18914 9220
rect 18236 9172 18288 9178
rect 18236 9114 18288 9120
rect 18420 9036 18472 9042
rect 18420 8978 18472 8984
rect 18432 8906 18460 8978
rect 18420 8900 18472 8906
rect 18420 8842 18472 8848
rect 18432 8809 18460 8842
rect 18418 8800 18474 8809
rect 18418 8735 18474 8744
rect 18606 8188 18914 8197
rect 18606 8186 18612 8188
rect 18668 8186 18692 8188
rect 18748 8186 18772 8188
rect 18828 8186 18852 8188
rect 18908 8186 18914 8188
rect 18668 8134 18670 8186
rect 18850 8134 18852 8186
rect 18606 8132 18612 8134
rect 18668 8132 18692 8134
rect 18748 8132 18772 8134
rect 18828 8132 18852 8134
rect 18908 8132 18914 8134
rect 18606 8123 18914 8132
rect 18606 7100 18914 7109
rect 18606 7098 18612 7100
rect 18668 7098 18692 7100
rect 18748 7098 18772 7100
rect 18828 7098 18852 7100
rect 18908 7098 18914 7100
rect 18668 7046 18670 7098
rect 18850 7046 18852 7098
rect 18606 7044 18612 7046
rect 18668 7044 18692 7046
rect 18748 7044 18772 7046
rect 18828 7044 18852 7046
rect 18908 7044 18914 7046
rect 18606 7035 18914 7044
rect 18420 6860 18472 6866
rect 18420 6802 18472 6808
rect 18432 6361 18460 6802
rect 18418 6352 18474 6361
rect 18418 6287 18474 6296
rect 18606 6012 18914 6021
rect 18606 6010 18612 6012
rect 18668 6010 18692 6012
rect 18748 6010 18772 6012
rect 18828 6010 18852 6012
rect 18908 6010 18914 6012
rect 18668 5958 18670 6010
rect 18850 5958 18852 6010
rect 18606 5956 18612 5958
rect 18668 5956 18692 5958
rect 18748 5956 18772 5958
rect 18828 5956 18852 5958
rect 18908 5956 18914 5958
rect 18606 5947 18914 5956
rect 18606 4924 18914 4933
rect 18606 4922 18612 4924
rect 18668 4922 18692 4924
rect 18748 4922 18772 4924
rect 18828 4922 18852 4924
rect 18908 4922 18914 4924
rect 18668 4870 18670 4922
rect 18850 4870 18852 4922
rect 18606 4868 18612 4870
rect 18668 4868 18692 4870
rect 18748 4868 18772 4870
rect 18828 4868 18852 4870
rect 18908 4868 18914 4870
rect 18606 4859 18914 4868
rect 19062 3904 19118 3913
rect 18606 3836 18914 3845
rect 19062 3839 19118 3848
rect 18606 3834 18612 3836
rect 18668 3834 18692 3836
rect 18748 3834 18772 3836
rect 18828 3834 18852 3836
rect 18908 3834 18914 3836
rect 18668 3782 18670 3834
rect 18850 3782 18852 3834
rect 18606 3780 18612 3782
rect 18668 3780 18692 3782
rect 18748 3780 18772 3782
rect 18828 3780 18852 3782
rect 18908 3780 18914 3782
rect 18606 3771 18914 3780
rect 18144 3732 18196 3738
rect 18144 3674 18196 3680
rect 19076 3602 19104 3839
rect 18420 3596 18472 3602
rect 18420 3538 18472 3544
rect 19064 3596 19116 3602
rect 19064 3538 19116 3544
rect 18432 3194 18460 3538
rect 18420 3188 18472 3194
rect 18420 3130 18472 3136
rect 18606 2748 18914 2757
rect 18606 2746 18612 2748
rect 18668 2746 18692 2748
rect 18748 2746 18772 2748
rect 18828 2746 18852 2748
rect 18908 2746 18914 2748
rect 18668 2694 18670 2746
rect 18850 2694 18852 2746
rect 18606 2692 18612 2694
rect 18668 2692 18692 2694
rect 18748 2692 18772 2694
rect 18828 2692 18852 2694
rect 18908 2692 18914 2694
rect 18606 2683 18914 2692
rect 17960 2032 18012 2038
rect 17960 1974 18012 1980
rect 17592 1556 17644 1562
rect 17592 1498 17644 1504
rect 17500 1420 17552 1426
rect 17500 1362 17552 1368
rect 16856 1352 16908 1358
rect 16856 1294 16908 1300
rect 17408 1352 17460 1358
rect 17408 1294 17460 1300
rect 17056 1116 17364 1125
rect 17056 1114 17062 1116
rect 17118 1114 17142 1116
rect 17198 1114 17222 1116
rect 17278 1114 17302 1116
rect 17358 1114 17364 1116
rect 17118 1062 17120 1114
rect 17300 1062 17302 1114
rect 17056 1060 17062 1062
rect 17118 1060 17142 1062
rect 17198 1060 17222 1062
rect 17278 1060 17302 1062
rect 17358 1060 17364 1062
rect 17056 1051 17364 1060
rect 15844 944 15896 950
rect 15844 886 15896 892
rect 17420 882 17448 1294
rect 17512 1018 17540 1362
rect 17972 1358 18000 1974
rect 18420 1760 18472 1766
rect 18420 1702 18472 1708
rect 18432 1465 18460 1702
rect 18606 1660 18914 1669
rect 18606 1658 18612 1660
rect 18668 1658 18692 1660
rect 18748 1658 18772 1660
rect 18828 1658 18852 1660
rect 18908 1658 18914 1660
rect 18668 1606 18670 1658
rect 18850 1606 18852 1658
rect 18606 1604 18612 1606
rect 18668 1604 18692 1606
rect 18748 1604 18772 1606
rect 18828 1604 18852 1606
rect 18908 1604 18914 1606
rect 18606 1595 18914 1604
rect 18418 1456 18474 1465
rect 18418 1391 18474 1400
rect 17960 1352 18012 1358
rect 17960 1294 18012 1300
rect 17592 1284 17644 1290
rect 17592 1226 17644 1232
rect 17604 1018 17632 1226
rect 17500 1012 17552 1018
rect 17500 954 17552 960
rect 17592 1012 17644 1018
rect 17592 954 17644 960
rect 17408 876 17460 882
rect 17408 818 17460 824
rect 17972 814 18000 1294
rect 3976 808 4028 814
rect 3976 750 4028 756
rect 5448 808 5500 814
rect 5448 750 5500 756
rect 8760 808 8812 814
rect 8760 750 8812 756
rect 9588 808 9640 814
rect 9588 750 9640 756
rect 17960 808 18012 814
rect 17960 750 18012 756
rect 3106 572 3414 581
rect 3106 570 3112 572
rect 3168 570 3192 572
rect 3248 570 3272 572
rect 3328 570 3352 572
rect 3408 570 3414 572
rect 3168 518 3170 570
rect 3350 518 3352 570
rect 3106 516 3112 518
rect 3168 516 3192 518
rect 3248 516 3272 518
rect 3328 516 3352 518
rect 3408 516 3414 518
rect 3106 507 3414 516
rect 6206 572 6514 581
rect 6206 570 6212 572
rect 6268 570 6292 572
rect 6348 570 6372 572
rect 6428 570 6452 572
rect 6508 570 6514 572
rect 6268 518 6270 570
rect 6450 518 6452 570
rect 6206 516 6212 518
rect 6268 516 6292 518
rect 6348 516 6372 518
rect 6428 516 6452 518
rect 6508 516 6514 518
rect 6206 507 6514 516
rect 9306 572 9614 581
rect 9306 570 9312 572
rect 9368 570 9392 572
rect 9448 570 9472 572
rect 9528 570 9552 572
rect 9608 570 9614 572
rect 9368 518 9370 570
rect 9550 518 9552 570
rect 9306 516 9312 518
rect 9368 516 9392 518
rect 9448 516 9472 518
rect 9528 516 9552 518
rect 9608 516 9614 518
rect 9306 507 9614 516
rect 12406 572 12714 581
rect 12406 570 12412 572
rect 12468 570 12492 572
rect 12548 570 12572 572
rect 12628 570 12652 572
rect 12708 570 12714 572
rect 12468 518 12470 570
rect 12650 518 12652 570
rect 12406 516 12412 518
rect 12468 516 12492 518
rect 12548 516 12572 518
rect 12628 516 12652 518
rect 12708 516 12714 518
rect 12406 507 12714 516
rect 15506 572 15814 581
rect 15506 570 15512 572
rect 15568 570 15592 572
rect 15648 570 15672 572
rect 15728 570 15752 572
rect 15808 570 15814 572
rect 15568 518 15570 570
rect 15750 518 15752 570
rect 15506 516 15512 518
rect 15568 516 15592 518
rect 15648 516 15672 518
rect 15728 516 15752 518
rect 15808 516 15814 518
rect 15506 507 15814 516
rect 18606 572 18914 581
rect 18606 570 18612 572
rect 18668 570 18692 572
rect 18748 570 18772 572
rect 18828 570 18852 572
rect 18908 570 18914 572
rect 18668 518 18670 570
rect 18850 518 18852 570
rect 18606 516 18612 518
rect 18668 516 18692 518
rect 18748 516 18772 518
rect 18828 516 18852 518
rect 18908 516 18914 518
rect 18606 507 18914 516
<< via2 >>
rect 1562 18522 1618 18524
rect 1642 18522 1698 18524
rect 1722 18522 1778 18524
rect 1802 18522 1858 18524
rect 1562 18470 1608 18522
rect 1608 18470 1618 18522
rect 1642 18470 1672 18522
rect 1672 18470 1684 18522
rect 1684 18470 1698 18522
rect 1722 18470 1736 18522
rect 1736 18470 1748 18522
rect 1748 18470 1778 18522
rect 1802 18470 1812 18522
rect 1812 18470 1858 18522
rect 1562 18468 1618 18470
rect 1642 18468 1698 18470
rect 1722 18468 1778 18470
rect 1802 18468 1858 18470
rect 1562 17434 1618 17436
rect 1642 17434 1698 17436
rect 1722 17434 1778 17436
rect 1802 17434 1858 17436
rect 1562 17382 1608 17434
rect 1608 17382 1618 17434
rect 1642 17382 1672 17434
rect 1672 17382 1684 17434
rect 1684 17382 1698 17434
rect 1722 17382 1736 17434
rect 1736 17382 1748 17434
rect 1748 17382 1778 17434
rect 1802 17382 1812 17434
rect 1812 17382 1858 17434
rect 1562 17380 1618 17382
rect 1642 17380 1698 17382
rect 1722 17380 1778 17382
rect 1802 17380 1858 17382
rect 1562 16346 1618 16348
rect 1642 16346 1698 16348
rect 1722 16346 1778 16348
rect 1802 16346 1858 16348
rect 1562 16294 1608 16346
rect 1608 16294 1618 16346
rect 1642 16294 1672 16346
rect 1672 16294 1684 16346
rect 1684 16294 1698 16346
rect 1722 16294 1736 16346
rect 1736 16294 1748 16346
rect 1748 16294 1778 16346
rect 1802 16294 1812 16346
rect 1812 16294 1858 16346
rect 1562 16292 1618 16294
rect 1642 16292 1698 16294
rect 1722 16292 1778 16294
rect 1802 16292 1858 16294
rect 1562 15258 1618 15260
rect 1642 15258 1698 15260
rect 1722 15258 1778 15260
rect 1802 15258 1858 15260
rect 1562 15206 1608 15258
rect 1608 15206 1618 15258
rect 1642 15206 1672 15258
rect 1672 15206 1684 15258
rect 1684 15206 1698 15258
rect 1722 15206 1736 15258
rect 1736 15206 1748 15258
rect 1748 15206 1778 15258
rect 1802 15206 1812 15258
rect 1812 15206 1858 15258
rect 1562 15204 1618 15206
rect 1642 15204 1698 15206
rect 1722 15204 1778 15206
rect 1802 15204 1858 15206
rect 1562 14170 1618 14172
rect 1642 14170 1698 14172
rect 1722 14170 1778 14172
rect 1802 14170 1858 14172
rect 1562 14118 1608 14170
rect 1608 14118 1618 14170
rect 1642 14118 1672 14170
rect 1672 14118 1684 14170
rect 1684 14118 1698 14170
rect 1722 14118 1736 14170
rect 1736 14118 1748 14170
rect 1748 14118 1778 14170
rect 1802 14118 1812 14170
rect 1812 14118 1858 14170
rect 1562 14116 1618 14118
rect 1642 14116 1698 14118
rect 1722 14116 1778 14118
rect 1802 14116 1858 14118
rect 1562 13082 1618 13084
rect 1642 13082 1698 13084
rect 1722 13082 1778 13084
rect 1802 13082 1858 13084
rect 1562 13030 1608 13082
rect 1608 13030 1618 13082
rect 1642 13030 1672 13082
rect 1672 13030 1684 13082
rect 1684 13030 1698 13082
rect 1722 13030 1736 13082
rect 1736 13030 1748 13082
rect 1748 13030 1778 13082
rect 1802 13030 1812 13082
rect 1812 13030 1858 13082
rect 1562 13028 1618 13030
rect 1642 13028 1698 13030
rect 1722 13028 1778 13030
rect 1802 13028 1858 13030
rect 1562 11994 1618 11996
rect 1642 11994 1698 11996
rect 1722 11994 1778 11996
rect 1802 11994 1858 11996
rect 1562 11942 1608 11994
rect 1608 11942 1618 11994
rect 1642 11942 1672 11994
rect 1672 11942 1684 11994
rect 1684 11942 1698 11994
rect 1722 11942 1736 11994
rect 1736 11942 1748 11994
rect 1748 11942 1778 11994
rect 1802 11942 1812 11994
rect 1812 11942 1858 11994
rect 1562 11940 1618 11942
rect 1642 11940 1698 11942
rect 1722 11940 1778 11942
rect 1802 11940 1858 11942
rect 3112 17978 3168 17980
rect 3192 17978 3248 17980
rect 3272 17978 3328 17980
rect 3352 17978 3408 17980
rect 3112 17926 3158 17978
rect 3158 17926 3168 17978
rect 3192 17926 3222 17978
rect 3222 17926 3234 17978
rect 3234 17926 3248 17978
rect 3272 17926 3286 17978
rect 3286 17926 3298 17978
rect 3298 17926 3328 17978
rect 3352 17926 3362 17978
rect 3362 17926 3408 17978
rect 3112 17924 3168 17926
rect 3192 17924 3248 17926
rect 3272 17924 3328 17926
rect 3352 17924 3408 17926
rect 3112 16890 3168 16892
rect 3192 16890 3248 16892
rect 3272 16890 3328 16892
rect 3352 16890 3408 16892
rect 3112 16838 3158 16890
rect 3158 16838 3168 16890
rect 3192 16838 3222 16890
rect 3222 16838 3234 16890
rect 3234 16838 3248 16890
rect 3272 16838 3286 16890
rect 3286 16838 3298 16890
rect 3298 16838 3328 16890
rect 3352 16838 3362 16890
rect 3362 16838 3408 16890
rect 3112 16836 3168 16838
rect 3192 16836 3248 16838
rect 3272 16836 3328 16838
rect 3352 16836 3408 16838
rect 4662 18522 4718 18524
rect 4742 18522 4798 18524
rect 4822 18522 4878 18524
rect 4902 18522 4958 18524
rect 4662 18470 4708 18522
rect 4708 18470 4718 18522
rect 4742 18470 4772 18522
rect 4772 18470 4784 18522
rect 4784 18470 4798 18522
rect 4822 18470 4836 18522
rect 4836 18470 4848 18522
rect 4848 18470 4878 18522
rect 4902 18470 4912 18522
rect 4912 18470 4958 18522
rect 4662 18468 4718 18470
rect 4742 18468 4798 18470
rect 4822 18468 4878 18470
rect 4902 18468 4958 18470
rect 3112 15802 3168 15804
rect 3192 15802 3248 15804
rect 3272 15802 3328 15804
rect 3352 15802 3408 15804
rect 3112 15750 3158 15802
rect 3158 15750 3168 15802
rect 3192 15750 3222 15802
rect 3222 15750 3234 15802
rect 3234 15750 3248 15802
rect 3272 15750 3286 15802
rect 3286 15750 3298 15802
rect 3298 15750 3328 15802
rect 3352 15750 3362 15802
rect 3362 15750 3408 15802
rect 3112 15748 3168 15750
rect 3192 15748 3248 15750
rect 3272 15748 3328 15750
rect 3352 15748 3408 15750
rect 4662 17434 4718 17436
rect 4742 17434 4798 17436
rect 4822 17434 4878 17436
rect 4902 17434 4958 17436
rect 4662 17382 4708 17434
rect 4708 17382 4718 17434
rect 4742 17382 4772 17434
rect 4772 17382 4784 17434
rect 4784 17382 4798 17434
rect 4822 17382 4836 17434
rect 4836 17382 4848 17434
rect 4848 17382 4878 17434
rect 4902 17382 4912 17434
rect 4912 17382 4958 17434
rect 4662 17380 4718 17382
rect 4742 17380 4798 17382
rect 4822 17380 4878 17382
rect 4902 17380 4958 17382
rect 4662 16346 4718 16348
rect 4742 16346 4798 16348
rect 4822 16346 4878 16348
rect 4902 16346 4958 16348
rect 4662 16294 4708 16346
rect 4708 16294 4718 16346
rect 4742 16294 4772 16346
rect 4772 16294 4784 16346
rect 4784 16294 4798 16346
rect 4822 16294 4836 16346
rect 4836 16294 4848 16346
rect 4848 16294 4878 16346
rect 4902 16294 4912 16346
rect 4912 16294 4958 16346
rect 4662 16292 4718 16294
rect 4742 16292 4798 16294
rect 4822 16292 4878 16294
rect 4902 16292 4958 16294
rect 3112 14714 3168 14716
rect 3192 14714 3248 14716
rect 3272 14714 3328 14716
rect 3352 14714 3408 14716
rect 3112 14662 3158 14714
rect 3158 14662 3168 14714
rect 3192 14662 3222 14714
rect 3222 14662 3234 14714
rect 3234 14662 3248 14714
rect 3272 14662 3286 14714
rect 3286 14662 3298 14714
rect 3298 14662 3328 14714
rect 3352 14662 3362 14714
rect 3362 14662 3408 14714
rect 3112 14660 3168 14662
rect 3192 14660 3248 14662
rect 3272 14660 3328 14662
rect 3352 14660 3408 14662
rect 3112 13626 3168 13628
rect 3192 13626 3248 13628
rect 3272 13626 3328 13628
rect 3352 13626 3408 13628
rect 3112 13574 3158 13626
rect 3158 13574 3168 13626
rect 3192 13574 3222 13626
rect 3222 13574 3234 13626
rect 3234 13574 3248 13626
rect 3272 13574 3286 13626
rect 3286 13574 3298 13626
rect 3298 13574 3328 13626
rect 3352 13574 3362 13626
rect 3362 13574 3408 13626
rect 3112 13572 3168 13574
rect 3192 13572 3248 13574
rect 3272 13572 3328 13574
rect 3352 13572 3408 13574
rect 7762 18522 7818 18524
rect 7842 18522 7898 18524
rect 7922 18522 7978 18524
rect 8002 18522 8058 18524
rect 7762 18470 7808 18522
rect 7808 18470 7818 18522
rect 7842 18470 7872 18522
rect 7872 18470 7884 18522
rect 7884 18470 7898 18522
rect 7922 18470 7936 18522
rect 7936 18470 7948 18522
rect 7948 18470 7978 18522
rect 8002 18470 8012 18522
rect 8012 18470 8058 18522
rect 7762 18468 7818 18470
rect 7842 18468 7898 18470
rect 7922 18468 7978 18470
rect 8002 18468 8058 18470
rect 10862 18522 10918 18524
rect 10942 18522 10998 18524
rect 11022 18522 11078 18524
rect 11102 18522 11158 18524
rect 10862 18470 10908 18522
rect 10908 18470 10918 18522
rect 10942 18470 10972 18522
rect 10972 18470 10984 18522
rect 10984 18470 10998 18522
rect 11022 18470 11036 18522
rect 11036 18470 11048 18522
rect 11048 18470 11078 18522
rect 11102 18470 11112 18522
rect 11112 18470 11158 18522
rect 10862 18468 10918 18470
rect 10942 18468 10998 18470
rect 11022 18468 11078 18470
rect 11102 18468 11158 18470
rect 6212 17978 6268 17980
rect 6292 17978 6348 17980
rect 6372 17978 6428 17980
rect 6452 17978 6508 17980
rect 6212 17926 6258 17978
rect 6258 17926 6268 17978
rect 6292 17926 6322 17978
rect 6322 17926 6334 17978
rect 6334 17926 6348 17978
rect 6372 17926 6386 17978
rect 6386 17926 6398 17978
rect 6398 17926 6428 17978
rect 6452 17926 6462 17978
rect 6462 17926 6508 17978
rect 6212 17924 6268 17926
rect 6292 17924 6348 17926
rect 6372 17924 6428 17926
rect 6452 17924 6508 17926
rect 6212 16890 6268 16892
rect 6292 16890 6348 16892
rect 6372 16890 6428 16892
rect 6452 16890 6508 16892
rect 6212 16838 6258 16890
rect 6258 16838 6268 16890
rect 6292 16838 6322 16890
rect 6322 16838 6334 16890
rect 6334 16838 6348 16890
rect 6372 16838 6386 16890
rect 6386 16838 6398 16890
rect 6398 16838 6428 16890
rect 6452 16838 6462 16890
rect 6462 16838 6508 16890
rect 6212 16836 6268 16838
rect 6292 16836 6348 16838
rect 6372 16836 6428 16838
rect 6452 16836 6508 16838
rect 6212 15802 6268 15804
rect 6292 15802 6348 15804
rect 6372 15802 6428 15804
rect 6452 15802 6508 15804
rect 6212 15750 6258 15802
rect 6258 15750 6268 15802
rect 6292 15750 6322 15802
rect 6322 15750 6334 15802
rect 6334 15750 6348 15802
rect 6372 15750 6386 15802
rect 6386 15750 6398 15802
rect 6398 15750 6428 15802
rect 6452 15750 6462 15802
rect 6462 15750 6508 15802
rect 6212 15748 6268 15750
rect 6292 15748 6348 15750
rect 6372 15748 6428 15750
rect 6452 15748 6508 15750
rect 4662 15258 4718 15260
rect 4742 15258 4798 15260
rect 4822 15258 4878 15260
rect 4902 15258 4958 15260
rect 4662 15206 4708 15258
rect 4708 15206 4718 15258
rect 4742 15206 4772 15258
rect 4772 15206 4784 15258
rect 4784 15206 4798 15258
rect 4822 15206 4836 15258
rect 4836 15206 4848 15258
rect 4848 15206 4878 15258
rect 4902 15206 4912 15258
rect 4912 15206 4958 15258
rect 4662 15204 4718 15206
rect 4742 15204 4798 15206
rect 4822 15204 4878 15206
rect 4902 15204 4958 15206
rect 3112 12538 3168 12540
rect 3192 12538 3248 12540
rect 3272 12538 3328 12540
rect 3352 12538 3408 12540
rect 3112 12486 3158 12538
rect 3158 12486 3168 12538
rect 3192 12486 3222 12538
rect 3222 12486 3234 12538
rect 3234 12486 3248 12538
rect 3272 12486 3286 12538
rect 3286 12486 3298 12538
rect 3298 12486 3328 12538
rect 3352 12486 3362 12538
rect 3362 12486 3408 12538
rect 3112 12484 3168 12486
rect 3192 12484 3248 12486
rect 3272 12484 3328 12486
rect 3352 12484 3408 12486
rect 4662 14170 4718 14172
rect 4742 14170 4798 14172
rect 4822 14170 4878 14172
rect 4902 14170 4958 14172
rect 4662 14118 4708 14170
rect 4708 14118 4718 14170
rect 4742 14118 4772 14170
rect 4772 14118 4784 14170
rect 4784 14118 4798 14170
rect 4822 14118 4836 14170
rect 4836 14118 4848 14170
rect 4848 14118 4878 14170
rect 4902 14118 4912 14170
rect 4912 14118 4958 14170
rect 4662 14116 4718 14118
rect 4742 14116 4798 14118
rect 4822 14116 4878 14118
rect 4902 14116 4958 14118
rect 7762 17434 7818 17436
rect 7842 17434 7898 17436
rect 7922 17434 7978 17436
rect 8002 17434 8058 17436
rect 7762 17382 7808 17434
rect 7808 17382 7818 17434
rect 7842 17382 7872 17434
rect 7872 17382 7884 17434
rect 7884 17382 7898 17434
rect 7922 17382 7936 17434
rect 7936 17382 7948 17434
rect 7948 17382 7978 17434
rect 8002 17382 8012 17434
rect 8012 17382 8058 17434
rect 7762 17380 7818 17382
rect 7842 17380 7898 17382
rect 7922 17380 7978 17382
rect 8002 17380 8058 17382
rect 6212 14714 6268 14716
rect 6292 14714 6348 14716
rect 6372 14714 6428 14716
rect 6452 14714 6508 14716
rect 6212 14662 6258 14714
rect 6258 14662 6268 14714
rect 6292 14662 6322 14714
rect 6322 14662 6334 14714
rect 6334 14662 6348 14714
rect 6372 14662 6386 14714
rect 6386 14662 6398 14714
rect 6398 14662 6428 14714
rect 6452 14662 6462 14714
rect 6462 14662 6508 14714
rect 6212 14660 6268 14662
rect 6292 14660 6348 14662
rect 6372 14660 6428 14662
rect 6452 14660 6508 14662
rect 6212 13626 6268 13628
rect 6292 13626 6348 13628
rect 6372 13626 6428 13628
rect 6452 13626 6508 13628
rect 6212 13574 6258 13626
rect 6258 13574 6268 13626
rect 6292 13574 6322 13626
rect 6322 13574 6334 13626
rect 6334 13574 6348 13626
rect 6372 13574 6386 13626
rect 6386 13574 6398 13626
rect 6398 13574 6428 13626
rect 6452 13574 6462 13626
rect 6462 13574 6508 13626
rect 6212 13572 6268 13574
rect 6292 13572 6348 13574
rect 6372 13572 6428 13574
rect 6452 13572 6508 13574
rect 3112 11450 3168 11452
rect 3192 11450 3248 11452
rect 3272 11450 3328 11452
rect 3352 11450 3408 11452
rect 3112 11398 3158 11450
rect 3158 11398 3168 11450
rect 3192 11398 3222 11450
rect 3222 11398 3234 11450
rect 3234 11398 3248 11450
rect 3272 11398 3286 11450
rect 3286 11398 3298 11450
rect 3298 11398 3328 11450
rect 3352 11398 3362 11450
rect 3362 11398 3408 11450
rect 3112 11396 3168 11398
rect 3192 11396 3248 11398
rect 3272 11396 3328 11398
rect 3352 11396 3408 11398
rect 1562 10906 1618 10908
rect 1642 10906 1698 10908
rect 1722 10906 1778 10908
rect 1802 10906 1858 10908
rect 1562 10854 1608 10906
rect 1608 10854 1618 10906
rect 1642 10854 1672 10906
rect 1672 10854 1684 10906
rect 1684 10854 1698 10906
rect 1722 10854 1736 10906
rect 1736 10854 1748 10906
rect 1748 10854 1778 10906
rect 1802 10854 1812 10906
rect 1812 10854 1858 10906
rect 1562 10852 1618 10854
rect 1642 10852 1698 10854
rect 1722 10852 1778 10854
rect 1802 10852 1858 10854
rect 1562 9818 1618 9820
rect 1642 9818 1698 9820
rect 1722 9818 1778 9820
rect 1802 9818 1858 9820
rect 1562 9766 1608 9818
rect 1608 9766 1618 9818
rect 1642 9766 1672 9818
rect 1672 9766 1684 9818
rect 1684 9766 1698 9818
rect 1722 9766 1736 9818
rect 1736 9766 1748 9818
rect 1748 9766 1778 9818
rect 1802 9766 1812 9818
rect 1812 9766 1858 9818
rect 1562 9764 1618 9766
rect 1642 9764 1698 9766
rect 1722 9764 1778 9766
rect 1802 9764 1858 9766
rect 1562 8730 1618 8732
rect 1642 8730 1698 8732
rect 1722 8730 1778 8732
rect 1802 8730 1858 8732
rect 1562 8678 1608 8730
rect 1608 8678 1618 8730
rect 1642 8678 1672 8730
rect 1672 8678 1684 8730
rect 1684 8678 1698 8730
rect 1722 8678 1736 8730
rect 1736 8678 1748 8730
rect 1748 8678 1778 8730
rect 1802 8678 1812 8730
rect 1812 8678 1858 8730
rect 1562 8676 1618 8678
rect 1642 8676 1698 8678
rect 1722 8676 1778 8678
rect 1802 8676 1858 8678
rect 1562 7642 1618 7644
rect 1642 7642 1698 7644
rect 1722 7642 1778 7644
rect 1802 7642 1858 7644
rect 1562 7590 1608 7642
rect 1608 7590 1618 7642
rect 1642 7590 1672 7642
rect 1672 7590 1684 7642
rect 1684 7590 1698 7642
rect 1722 7590 1736 7642
rect 1736 7590 1748 7642
rect 1748 7590 1778 7642
rect 1802 7590 1812 7642
rect 1812 7590 1858 7642
rect 1562 7588 1618 7590
rect 1642 7588 1698 7590
rect 1722 7588 1778 7590
rect 1802 7588 1858 7590
rect 3112 10362 3168 10364
rect 3192 10362 3248 10364
rect 3272 10362 3328 10364
rect 3352 10362 3408 10364
rect 3112 10310 3158 10362
rect 3158 10310 3168 10362
rect 3192 10310 3222 10362
rect 3222 10310 3234 10362
rect 3234 10310 3248 10362
rect 3272 10310 3286 10362
rect 3286 10310 3298 10362
rect 3298 10310 3328 10362
rect 3352 10310 3362 10362
rect 3362 10310 3408 10362
rect 3112 10308 3168 10310
rect 3192 10308 3248 10310
rect 3272 10308 3328 10310
rect 3352 10308 3408 10310
rect 4662 13082 4718 13084
rect 4742 13082 4798 13084
rect 4822 13082 4878 13084
rect 4902 13082 4958 13084
rect 4662 13030 4708 13082
rect 4708 13030 4718 13082
rect 4742 13030 4772 13082
rect 4772 13030 4784 13082
rect 4784 13030 4798 13082
rect 4822 13030 4836 13082
rect 4836 13030 4848 13082
rect 4848 13030 4878 13082
rect 4902 13030 4912 13082
rect 4912 13030 4958 13082
rect 4662 13028 4718 13030
rect 4742 13028 4798 13030
rect 4822 13028 4878 13030
rect 4902 13028 4958 13030
rect 4662 11994 4718 11996
rect 4742 11994 4798 11996
rect 4822 11994 4878 11996
rect 4902 11994 4958 11996
rect 4662 11942 4708 11994
rect 4708 11942 4718 11994
rect 4742 11942 4772 11994
rect 4772 11942 4784 11994
rect 4784 11942 4798 11994
rect 4822 11942 4836 11994
rect 4836 11942 4848 11994
rect 4848 11942 4878 11994
rect 4902 11942 4912 11994
rect 4912 11942 4958 11994
rect 4662 11940 4718 11942
rect 4742 11940 4798 11942
rect 4822 11940 4878 11942
rect 4902 11940 4958 11942
rect 4662 10906 4718 10908
rect 4742 10906 4798 10908
rect 4822 10906 4878 10908
rect 4902 10906 4958 10908
rect 4662 10854 4708 10906
rect 4708 10854 4718 10906
rect 4742 10854 4772 10906
rect 4772 10854 4784 10906
rect 4784 10854 4798 10906
rect 4822 10854 4836 10906
rect 4836 10854 4848 10906
rect 4848 10854 4878 10906
rect 4902 10854 4912 10906
rect 4912 10854 4958 10906
rect 4662 10852 4718 10854
rect 4742 10852 4798 10854
rect 4822 10852 4878 10854
rect 4902 10852 4958 10854
rect 3112 9274 3168 9276
rect 3192 9274 3248 9276
rect 3272 9274 3328 9276
rect 3352 9274 3408 9276
rect 3112 9222 3158 9274
rect 3158 9222 3168 9274
rect 3192 9222 3222 9274
rect 3222 9222 3234 9274
rect 3234 9222 3248 9274
rect 3272 9222 3286 9274
rect 3286 9222 3298 9274
rect 3298 9222 3328 9274
rect 3352 9222 3362 9274
rect 3362 9222 3408 9274
rect 3112 9220 3168 9222
rect 3192 9220 3248 9222
rect 3272 9220 3328 9222
rect 3352 9220 3408 9222
rect 1562 6554 1618 6556
rect 1642 6554 1698 6556
rect 1722 6554 1778 6556
rect 1802 6554 1858 6556
rect 1562 6502 1608 6554
rect 1608 6502 1618 6554
rect 1642 6502 1672 6554
rect 1672 6502 1684 6554
rect 1684 6502 1698 6554
rect 1722 6502 1736 6554
rect 1736 6502 1748 6554
rect 1748 6502 1778 6554
rect 1802 6502 1812 6554
rect 1812 6502 1858 6554
rect 1562 6500 1618 6502
rect 1642 6500 1698 6502
rect 1722 6500 1778 6502
rect 1802 6500 1858 6502
rect 1562 5466 1618 5468
rect 1642 5466 1698 5468
rect 1722 5466 1778 5468
rect 1802 5466 1858 5468
rect 1562 5414 1608 5466
rect 1608 5414 1618 5466
rect 1642 5414 1672 5466
rect 1672 5414 1684 5466
rect 1684 5414 1698 5466
rect 1722 5414 1736 5466
rect 1736 5414 1748 5466
rect 1748 5414 1778 5466
rect 1802 5414 1812 5466
rect 1812 5414 1858 5466
rect 1562 5412 1618 5414
rect 1642 5412 1698 5414
rect 1722 5412 1778 5414
rect 1802 5412 1858 5414
rect 1562 4378 1618 4380
rect 1642 4378 1698 4380
rect 1722 4378 1778 4380
rect 1802 4378 1858 4380
rect 1562 4326 1608 4378
rect 1608 4326 1618 4378
rect 1642 4326 1672 4378
rect 1672 4326 1684 4378
rect 1684 4326 1698 4378
rect 1722 4326 1736 4378
rect 1736 4326 1748 4378
rect 1748 4326 1778 4378
rect 1802 4326 1812 4378
rect 1812 4326 1858 4378
rect 1562 4324 1618 4326
rect 1642 4324 1698 4326
rect 1722 4324 1778 4326
rect 1802 4324 1858 4326
rect 3112 8186 3168 8188
rect 3192 8186 3248 8188
rect 3272 8186 3328 8188
rect 3352 8186 3408 8188
rect 3112 8134 3158 8186
rect 3158 8134 3168 8186
rect 3192 8134 3222 8186
rect 3222 8134 3234 8186
rect 3234 8134 3248 8186
rect 3272 8134 3286 8186
rect 3286 8134 3298 8186
rect 3298 8134 3328 8186
rect 3352 8134 3362 8186
rect 3362 8134 3408 8186
rect 3112 8132 3168 8134
rect 3192 8132 3248 8134
rect 3272 8132 3328 8134
rect 3352 8132 3408 8134
rect 3112 7098 3168 7100
rect 3192 7098 3248 7100
rect 3272 7098 3328 7100
rect 3352 7098 3408 7100
rect 3112 7046 3158 7098
rect 3158 7046 3168 7098
rect 3192 7046 3222 7098
rect 3222 7046 3234 7098
rect 3234 7046 3248 7098
rect 3272 7046 3286 7098
rect 3286 7046 3298 7098
rect 3298 7046 3328 7098
rect 3352 7046 3362 7098
rect 3362 7046 3408 7098
rect 3112 7044 3168 7046
rect 3192 7044 3248 7046
rect 3272 7044 3328 7046
rect 3352 7044 3408 7046
rect 1562 3290 1618 3292
rect 1642 3290 1698 3292
rect 1722 3290 1778 3292
rect 1802 3290 1858 3292
rect 1562 3238 1608 3290
rect 1608 3238 1618 3290
rect 1642 3238 1672 3290
rect 1672 3238 1684 3290
rect 1684 3238 1698 3290
rect 1722 3238 1736 3290
rect 1736 3238 1748 3290
rect 1748 3238 1778 3290
rect 1802 3238 1812 3290
rect 1812 3238 1858 3290
rect 1562 3236 1618 3238
rect 1642 3236 1698 3238
rect 1722 3236 1778 3238
rect 1802 3236 1858 3238
rect 3112 6010 3168 6012
rect 3192 6010 3248 6012
rect 3272 6010 3328 6012
rect 3352 6010 3408 6012
rect 3112 5958 3158 6010
rect 3158 5958 3168 6010
rect 3192 5958 3222 6010
rect 3222 5958 3234 6010
rect 3234 5958 3248 6010
rect 3272 5958 3286 6010
rect 3286 5958 3298 6010
rect 3298 5958 3328 6010
rect 3352 5958 3362 6010
rect 3362 5958 3408 6010
rect 3112 5956 3168 5958
rect 3192 5956 3248 5958
rect 3272 5956 3328 5958
rect 3352 5956 3408 5958
rect 3112 4922 3168 4924
rect 3192 4922 3248 4924
rect 3272 4922 3328 4924
rect 3352 4922 3408 4924
rect 3112 4870 3158 4922
rect 3158 4870 3168 4922
rect 3192 4870 3222 4922
rect 3222 4870 3234 4922
rect 3234 4870 3248 4922
rect 3272 4870 3286 4922
rect 3286 4870 3298 4922
rect 3298 4870 3328 4922
rect 3352 4870 3362 4922
rect 3362 4870 3408 4922
rect 3112 4868 3168 4870
rect 3192 4868 3248 4870
rect 3272 4868 3328 4870
rect 3352 4868 3408 4870
rect 1562 2202 1618 2204
rect 1642 2202 1698 2204
rect 1722 2202 1778 2204
rect 1802 2202 1858 2204
rect 1562 2150 1608 2202
rect 1608 2150 1618 2202
rect 1642 2150 1672 2202
rect 1672 2150 1684 2202
rect 1684 2150 1698 2202
rect 1722 2150 1736 2202
rect 1736 2150 1748 2202
rect 1748 2150 1778 2202
rect 1802 2150 1812 2202
rect 1812 2150 1858 2202
rect 1562 2148 1618 2150
rect 1642 2148 1698 2150
rect 1722 2148 1778 2150
rect 1802 2148 1858 2150
rect 3112 3834 3168 3836
rect 3192 3834 3248 3836
rect 3272 3834 3328 3836
rect 3352 3834 3408 3836
rect 3112 3782 3158 3834
rect 3158 3782 3168 3834
rect 3192 3782 3222 3834
rect 3222 3782 3234 3834
rect 3234 3782 3248 3834
rect 3272 3782 3286 3834
rect 3286 3782 3298 3834
rect 3298 3782 3328 3834
rect 3352 3782 3362 3834
rect 3362 3782 3408 3834
rect 3112 3780 3168 3782
rect 3192 3780 3248 3782
rect 3272 3780 3328 3782
rect 3352 3780 3408 3782
rect 3112 2746 3168 2748
rect 3192 2746 3248 2748
rect 3272 2746 3328 2748
rect 3352 2746 3408 2748
rect 3112 2694 3158 2746
rect 3158 2694 3168 2746
rect 3192 2694 3222 2746
rect 3222 2694 3234 2746
rect 3234 2694 3248 2746
rect 3272 2694 3286 2746
rect 3286 2694 3298 2746
rect 3298 2694 3328 2746
rect 3352 2694 3362 2746
rect 3362 2694 3408 2746
rect 3112 2692 3168 2694
rect 3192 2692 3248 2694
rect 3272 2692 3328 2694
rect 3352 2692 3408 2694
rect 4662 9818 4718 9820
rect 4742 9818 4798 9820
rect 4822 9818 4878 9820
rect 4902 9818 4958 9820
rect 4662 9766 4708 9818
rect 4708 9766 4718 9818
rect 4742 9766 4772 9818
rect 4772 9766 4784 9818
rect 4784 9766 4798 9818
rect 4822 9766 4836 9818
rect 4836 9766 4848 9818
rect 4848 9766 4878 9818
rect 4902 9766 4912 9818
rect 4912 9766 4958 9818
rect 4662 9764 4718 9766
rect 4742 9764 4798 9766
rect 4822 9764 4878 9766
rect 4902 9764 4958 9766
rect 4662 8730 4718 8732
rect 4742 8730 4798 8732
rect 4822 8730 4878 8732
rect 4902 8730 4958 8732
rect 4662 8678 4708 8730
rect 4708 8678 4718 8730
rect 4742 8678 4772 8730
rect 4772 8678 4784 8730
rect 4784 8678 4798 8730
rect 4822 8678 4836 8730
rect 4836 8678 4848 8730
rect 4848 8678 4878 8730
rect 4902 8678 4912 8730
rect 4912 8678 4958 8730
rect 4662 8676 4718 8678
rect 4742 8676 4798 8678
rect 4822 8676 4878 8678
rect 4902 8676 4958 8678
rect 4662 7642 4718 7644
rect 4742 7642 4798 7644
rect 4822 7642 4878 7644
rect 4902 7642 4958 7644
rect 4662 7590 4708 7642
rect 4708 7590 4718 7642
rect 4742 7590 4772 7642
rect 4772 7590 4784 7642
rect 4784 7590 4798 7642
rect 4822 7590 4836 7642
rect 4836 7590 4848 7642
rect 4848 7590 4878 7642
rect 4902 7590 4912 7642
rect 4912 7590 4958 7642
rect 4662 7588 4718 7590
rect 4742 7588 4798 7590
rect 4822 7588 4878 7590
rect 4902 7588 4958 7590
rect 4662 6554 4718 6556
rect 4742 6554 4798 6556
rect 4822 6554 4878 6556
rect 4902 6554 4958 6556
rect 4662 6502 4708 6554
rect 4708 6502 4718 6554
rect 4742 6502 4772 6554
rect 4772 6502 4784 6554
rect 4784 6502 4798 6554
rect 4822 6502 4836 6554
rect 4836 6502 4848 6554
rect 4848 6502 4878 6554
rect 4902 6502 4912 6554
rect 4912 6502 4958 6554
rect 4662 6500 4718 6502
rect 4742 6500 4798 6502
rect 4822 6500 4878 6502
rect 4902 6500 4958 6502
rect 6212 12538 6268 12540
rect 6292 12538 6348 12540
rect 6372 12538 6428 12540
rect 6452 12538 6508 12540
rect 6212 12486 6258 12538
rect 6258 12486 6268 12538
rect 6292 12486 6322 12538
rect 6322 12486 6334 12538
rect 6334 12486 6348 12538
rect 6372 12486 6386 12538
rect 6386 12486 6398 12538
rect 6398 12486 6428 12538
rect 6452 12486 6462 12538
rect 6462 12486 6508 12538
rect 6212 12484 6268 12486
rect 6292 12484 6348 12486
rect 6372 12484 6428 12486
rect 6452 12484 6508 12486
rect 7762 16346 7818 16348
rect 7842 16346 7898 16348
rect 7922 16346 7978 16348
rect 8002 16346 8058 16348
rect 7762 16294 7808 16346
rect 7808 16294 7818 16346
rect 7842 16294 7872 16346
rect 7872 16294 7884 16346
rect 7884 16294 7898 16346
rect 7922 16294 7936 16346
rect 7936 16294 7948 16346
rect 7948 16294 7978 16346
rect 8002 16294 8012 16346
rect 8012 16294 8058 16346
rect 7762 16292 7818 16294
rect 7842 16292 7898 16294
rect 7922 16292 7978 16294
rect 8002 16292 8058 16294
rect 7762 15258 7818 15260
rect 7842 15258 7898 15260
rect 7922 15258 7978 15260
rect 8002 15258 8058 15260
rect 7762 15206 7808 15258
rect 7808 15206 7818 15258
rect 7842 15206 7872 15258
rect 7872 15206 7884 15258
rect 7884 15206 7898 15258
rect 7922 15206 7936 15258
rect 7936 15206 7948 15258
rect 7948 15206 7978 15258
rect 8002 15206 8012 15258
rect 8012 15206 8058 15258
rect 7762 15204 7818 15206
rect 7842 15204 7898 15206
rect 7922 15204 7978 15206
rect 8002 15204 8058 15206
rect 6212 11450 6268 11452
rect 6292 11450 6348 11452
rect 6372 11450 6428 11452
rect 6452 11450 6508 11452
rect 6212 11398 6258 11450
rect 6258 11398 6268 11450
rect 6292 11398 6322 11450
rect 6322 11398 6334 11450
rect 6334 11398 6348 11450
rect 6372 11398 6386 11450
rect 6386 11398 6398 11450
rect 6398 11398 6428 11450
rect 6452 11398 6462 11450
rect 6462 11398 6508 11450
rect 6212 11396 6268 11398
rect 6292 11396 6348 11398
rect 6372 11396 6428 11398
rect 6452 11396 6508 11398
rect 6212 10362 6268 10364
rect 6292 10362 6348 10364
rect 6372 10362 6428 10364
rect 6452 10362 6508 10364
rect 6212 10310 6258 10362
rect 6258 10310 6268 10362
rect 6292 10310 6322 10362
rect 6322 10310 6334 10362
rect 6334 10310 6348 10362
rect 6372 10310 6386 10362
rect 6386 10310 6398 10362
rect 6398 10310 6428 10362
rect 6452 10310 6462 10362
rect 6462 10310 6508 10362
rect 6212 10308 6268 10310
rect 6292 10308 6348 10310
rect 6372 10308 6428 10310
rect 6452 10308 6508 10310
rect 6212 9274 6268 9276
rect 6292 9274 6348 9276
rect 6372 9274 6428 9276
rect 6452 9274 6508 9276
rect 6212 9222 6258 9274
rect 6258 9222 6268 9274
rect 6292 9222 6322 9274
rect 6322 9222 6334 9274
rect 6334 9222 6348 9274
rect 6372 9222 6386 9274
rect 6386 9222 6398 9274
rect 6398 9222 6428 9274
rect 6452 9222 6462 9274
rect 6462 9222 6508 9274
rect 6212 9220 6268 9222
rect 6292 9220 6348 9222
rect 6372 9220 6428 9222
rect 6452 9220 6508 9222
rect 6212 8186 6268 8188
rect 6292 8186 6348 8188
rect 6372 8186 6428 8188
rect 6452 8186 6508 8188
rect 6212 8134 6258 8186
rect 6258 8134 6268 8186
rect 6292 8134 6322 8186
rect 6322 8134 6334 8186
rect 6334 8134 6348 8186
rect 6372 8134 6386 8186
rect 6386 8134 6398 8186
rect 6398 8134 6428 8186
rect 6452 8134 6462 8186
rect 6462 8134 6508 8186
rect 6212 8132 6268 8134
rect 6292 8132 6348 8134
rect 6372 8132 6428 8134
rect 6452 8132 6508 8134
rect 9312 17978 9368 17980
rect 9392 17978 9448 17980
rect 9472 17978 9528 17980
rect 9552 17978 9608 17980
rect 9312 17926 9358 17978
rect 9358 17926 9368 17978
rect 9392 17926 9422 17978
rect 9422 17926 9434 17978
rect 9434 17926 9448 17978
rect 9472 17926 9486 17978
rect 9486 17926 9498 17978
rect 9498 17926 9528 17978
rect 9552 17926 9562 17978
rect 9562 17926 9608 17978
rect 9312 17924 9368 17926
rect 9392 17924 9448 17926
rect 9472 17924 9528 17926
rect 9552 17924 9608 17926
rect 9312 16890 9368 16892
rect 9392 16890 9448 16892
rect 9472 16890 9528 16892
rect 9552 16890 9608 16892
rect 9312 16838 9358 16890
rect 9358 16838 9368 16890
rect 9392 16838 9422 16890
rect 9422 16838 9434 16890
rect 9434 16838 9448 16890
rect 9472 16838 9486 16890
rect 9486 16838 9498 16890
rect 9498 16838 9528 16890
rect 9552 16838 9562 16890
rect 9562 16838 9608 16890
rect 9312 16836 9368 16838
rect 9392 16836 9448 16838
rect 9472 16836 9528 16838
rect 9552 16836 9608 16838
rect 7762 14170 7818 14172
rect 7842 14170 7898 14172
rect 7922 14170 7978 14172
rect 8002 14170 8058 14172
rect 7762 14118 7808 14170
rect 7808 14118 7818 14170
rect 7842 14118 7872 14170
rect 7872 14118 7884 14170
rect 7884 14118 7898 14170
rect 7922 14118 7936 14170
rect 7936 14118 7948 14170
rect 7948 14118 7978 14170
rect 8002 14118 8012 14170
rect 8012 14118 8058 14170
rect 7762 14116 7818 14118
rect 7842 14116 7898 14118
rect 7922 14116 7978 14118
rect 8002 14116 8058 14118
rect 9312 15802 9368 15804
rect 9392 15802 9448 15804
rect 9472 15802 9528 15804
rect 9552 15802 9608 15804
rect 9312 15750 9358 15802
rect 9358 15750 9368 15802
rect 9392 15750 9422 15802
rect 9422 15750 9434 15802
rect 9434 15750 9448 15802
rect 9472 15750 9486 15802
rect 9486 15750 9498 15802
rect 9498 15750 9528 15802
rect 9552 15750 9562 15802
rect 9562 15750 9608 15802
rect 9312 15748 9368 15750
rect 9392 15748 9448 15750
rect 9472 15748 9528 15750
rect 9552 15748 9608 15750
rect 10862 17434 10918 17436
rect 10942 17434 10998 17436
rect 11022 17434 11078 17436
rect 11102 17434 11158 17436
rect 10862 17382 10908 17434
rect 10908 17382 10918 17434
rect 10942 17382 10972 17434
rect 10972 17382 10984 17434
rect 10984 17382 10998 17434
rect 11022 17382 11036 17434
rect 11036 17382 11048 17434
rect 11048 17382 11078 17434
rect 11102 17382 11112 17434
rect 11112 17382 11158 17434
rect 10862 17380 10918 17382
rect 10942 17380 10998 17382
rect 11022 17380 11078 17382
rect 11102 17380 11158 17382
rect 7762 13082 7818 13084
rect 7842 13082 7898 13084
rect 7922 13082 7978 13084
rect 8002 13082 8058 13084
rect 7762 13030 7808 13082
rect 7808 13030 7818 13082
rect 7842 13030 7872 13082
rect 7872 13030 7884 13082
rect 7884 13030 7898 13082
rect 7922 13030 7936 13082
rect 7936 13030 7948 13082
rect 7948 13030 7978 13082
rect 8002 13030 8012 13082
rect 8012 13030 8058 13082
rect 7762 13028 7818 13030
rect 7842 13028 7898 13030
rect 7922 13028 7978 13030
rect 8002 13028 8058 13030
rect 7762 11994 7818 11996
rect 7842 11994 7898 11996
rect 7922 11994 7978 11996
rect 8002 11994 8058 11996
rect 7762 11942 7808 11994
rect 7808 11942 7818 11994
rect 7842 11942 7872 11994
rect 7872 11942 7884 11994
rect 7884 11942 7898 11994
rect 7922 11942 7936 11994
rect 7936 11942 7948 11994
rect 7948 11942 7978 11994
rect 8002 11942 8012 11994
rect 8012 11942 8058 11994
rect 7762 11940 7818 11942
rect 7842 11940 7898 11942
rect 7922 11940 7978 11942
rect 8002 11940 8058 11942
rect 7762 10906 7818 10908
rect 7842 10906 7898 10908
rect 7922 10906 7978 10908
rect 8002 10906 8058 10908
rect 7762 10854 7808 10906
rect 7808 10854 7818 10906
rect 7842 10854 7872 10906
rect 7872 10854 7884 10906
rect 7884 10854 7898 10906
rect 7922 10854 7936 10906
rect 7936 10854 7948 10906
rect 7948 10854 7978 10906
rect 8002 10854 8012 10906
rect 8012 10854 8058 10906
rect 7762 10852 7818 10854
rect 7842 10852 7898 10854
rect 7922 10852 7978 10854
rect 8002 10852 8058 10854
rect 7762 9818 7818 9820
rect 7842 9818 7898 9820
rect 7922 9818 7978 9820
rect 8002 9818 8058 9820
rect 7762 9766 7808 9818
rect 7808 9766 7818 9818
rect 7842 9766 7872 9818
rect 7872 9766 7884 9818
rect 7884 9766 7898 9818
rect 7922 9766 7936 9818
rect 7936 9766 7948 9818
rect 7948 9766 7978 9818
rect 8002 9766 8012 9818
rect 8012 9766 8058 9818
rect 7762 9764 7818 9766
rect 7842 9764 7898 9766
rect 7922 9764 7978 9766
rect 8002 9764 8058 9766
rect 7762 8730 7818 8732
rect 7842 8730 7898 8732
rect 7922 8730 7978 8732
rect 8002 8730 8058 8732
rect 7762 8678 7808 8730
rect 7808 8678 7818 8730
rect 7842 8678 7872 8730
rect 7872 8678 7884 8730
rect 7884 8678 7898 8730
rect 7922 8678 7936 8730
rect 7936 8678 7948 8730
rect 7948 8678 7978 8730
rect 8002 8678 8012 8730
rect 8012 8678 8058 8730
rect 7762 8676 7818 8678
rect 7842 8676 7898 8678
rect 7922 8676 7978 8678
rect 8002 8676 8058 8678
rect 4662 5466 4718 5468
rect 4742 5466 4798 5468
rect 4822 5466 4878 5468
rect 4902 5466 4958 5468
rect 4662 5414 4708 5466
rect 4708 5414 4718 5466
rect 4742 5414 4772 5466
rect 4772 5414 4784 5466
rect 4784 5414 4798 5466
rect 4822 5414 4836 5466
rect 4836 5414 4848 5466
rect 4848 5414 4878 5466
rect 4902 5414 4912 5466
rect 4912 5414 4958 5466
rect 4662 5412 4718 5414
rect 4742 5412 4798 5414
rect 4822 5412 4878 5414
rect 4902 5412 4958 5414
rect 4662 4378 4718 4380
rect 4742 4378 4798 4380
rect 4822 4378 4878 4380
rect 4902 4378 4958 4380
rect 4662 4326 4708 4378
rect 4708 4326 4718 4378
rect 4742 4326 4772 4378
rect 4772 4326 4784 4378
rect 4784 4326 4798 4378
rect 4822 4326 4836 4378
rect 4836 4326 4848 4378
rect 4848 4326 4878 4378
rect 4902 4326 4912 4378
rect 4912 4326 4958 4378
rect 4662 4324 4718 4326
rect 4742 4324 4798 4326
rect 4822 4324 4878 4326
rect 4902 4324 4958 4326
rect 1562 1114 1618 1116
rect 1642 1114 1698 1116
rect 1722 1114 1778 1116
rect 1802 1114 1858 1116
rect 1562 1062 1608 1114
rect 1608 1062 1618 1114
rect 1642 1062 1672 1114
rect 1672 1062 1684 1114
rect 1684 1062 1698 1114
rect 1722 1062 1736 1114
rect 1736 1062 1748 1114
rect 1748 1062 1778 1114
rect 1802 1062 1812 1114
rect 1812 1062 1858 1114
rect 1562 1060 1618 1062
rect 1642 1060 1698 1062
rect 1722 1060 1778 1062
rect 1802 1060 1858 1062
rect 3112 1658 3168 1660
rect 3192 1658 3248 1660
rect 3272 1658 3328 1660
rect 3352 1658 3408 1660
rect 3112 1606 3158 1658
rect 3158 1606 3168 1658
rect 3192 1606 3222 1658
rect 3222 1606 3234 1658
rect 3234 1606 3248 1658
rect 3272 1606 3286 1658
rect 3286 1606 3298 1658
rect 3298 1606 3328 1658
rect 3352 1606 3362 1658
rect 3362 1606 3408 1658
rect 3112 1604 3168 1606
rect 3192 1604 3248 1606
rect 3272 1604 3328 1606
rect 3352 1604 3408 1606
rect 6212 7098 6268 7100
rect 6292 7098 6348 7100
rect 6372 7098 6428 7100
rect 6452 7098 6508 7100
rect 6212 7046 6258 7098
rect 6258 7046 6268 7098
rect 6292 7046 6322 7098
rect 6322 7046 6334 7098
rect 6334 7046 6348 7098
rect 6372 7046 6386 7098
rect 6386 7046 6398 7098
rect 6398 7046 6428 7098
rect 6452 7046 6462 7098
rect 6462 7046 6508 7098
rect 6212 7044 6268 7046
rect 6292 7044 6348 7046
rect 6372 7044 6428 7046
rect 6452 7044 6508 7046
rect 4662 3290 4718 3292
rect 4742 3290 4798 3292
rect 4822 3290 4878 3292
rect 4902 3290 4958 3292
rect 4662 3238 4708 3290
rect 4708 3238 4718 3290
rect 4742 3238 4772 3290
rect 4772 3238 4784 3290
rect 4784 3238 4798 3290
rect 4822 3238 4836 3290
rect 4836 3238 4848 3290
rect 4848 3238 4878 3290
rect 4902 3238 4912 3290
rect 4912 3238 4958 3290
rect 4662 3236 4718 3238
rect 4742 3236 4798 3238
rect 4822 3236 4878 3238
rect 4902 3236 4958 3238
rect 6212 6010 6268 6012
rect 6292 6010 6348 6012
rect 6372 6010 6428 6012
rect 6452 6010 6508 6012
rect 6212 5958 6258 6010
rect 6258 5958 6268 6010
rect 6292 5958 6322 6010
rect 6322 5958 6334 6010
rect 6334 5958 6348 6010
rect 6372 5958 6386 6010
rect 6386 5958 6398 6010
rect 6398 5958 6428 6010
rect 6452 5958 6462 6010
rect 6462 5958 6508 6010
rect 6212 5956 6268 5958
rect 6292 5956 6348 5958
rect 6372 5956 6428 5958
rect 6452 5956 6508 5958
rect 6212 4922 6268 4924
rect 6292 4922 6348 4924
rect 6372 4922 6428 4924
rect 6452 4922 6508 4924
rect 6212 4870 6258 4922
rect 6258 4870 6268 4922
rect 6292 4870 6322 4922
rect 6322 4870 6334 4922
rect 6334 4870 6348 4922
rect 6372 4870 6386 4922
rect 6386 4870 6398 4922
rect 6398 4870 6428 4922
rect 6452 4870 6462 4922
rect 6462 4870 6508 4922
rect 6212 4868 6268 4870
rect 6292 4868 6348 4870
rect 6372 4868 6428 4870
rect 6452 4868 6508 4870
rect 6212 3834 6268 3836
rect 6292 3834 6348 3836
rect 6372 3834 6428 3836
rect 6452 3834 6508 3836
rect 6212 3782 6258 3834
rect 6258 3782 6268 3834
rect 6292 3782 6322 3834
rect 6322 3782 6334 3834
rect 6334 3782 6348 3834
rect 6372 3782 6386 3834
rect 6386 3782 6398 3834
rect 6398 3782 6428 3834
rect 6452 3782 6462 3834
rect 6462 3782 6508 3834
rect 6212 3780 6268 3782
rect 6292 3780 6348 3782
rect 6372 3780 6428 3782
rect 6452 3780 6508 3782
rect 7762 7642 7818 7644
rect 7842 7642 7898 7644
rect 7922 7642 7978 7644
rect 8002 7642 8058 7644
rect 7762 7590 7808 7642
rect 7808 7590 7818 7642
rect 7842 7590 7872 7642
rect 7872 7590 7884 7642
rect 7884 7590 7898 7642
rect 7922 7590 7936 7642
rect 7936 7590 7948 7642
rect 7948 7590 7978 7642
rect 8002 7590 8012 7642
rect 8012 7590 8058 7642
rect 7762 7588 7818 7590
rect 7842 7588 7898 7590
rect 7922 7588 7978 7590
rect 8002 7588 8058 7590
rect 7762 6554 7818 6556
rect 7842 6554 7898 6556
rect 7922 6554 7978 6556
rect 8002 6554 8058 6556
rect 7762 6502 7808 6554
rect 7808 6502 7818 6554
rect 7842 6502 7872 6554
rect 7872 6502 7884 6554
rect 7884 6502 7898 6554
rect 7922 6502 7936 6554
rect 7936 6502 7948 6554
rect 7948 6502 7978 6554
rect 8002 6502 8012 6554
rect 8012 6502 8058 6554
rect 7762 6500 7818 6502
rect 7842 6500 7898 6502
rect 7922 6500 7978 6502
rect 8002 6500 8058 6502
rect 7762 5466 7818 5468
rect 7842 5466 7898 5468
rect 7922 5466 7978 5468
rect 8002 5466 8058 5468
rect 7762 5414 7808 5466
rect 7808 5414 7818 5466
rect 7842 5414 7872 5466
rect 7872 5414 7884 5466
rect 7884 5414 7898 5466
rect 7922 5414 7936 5466
rect 7936 5414 7948 5466
rect 7948 5414 7978 5466
rect 8002 5414 8012 5466
rect 8012 5414 8058 5466
rect 7762 5412 7818 5414
rect 7842 5412 7898 5414
rect 7922 5412 7978 5414
rect 8002 5412 8058 5414
rect 7762 4378 7818 4380
rect 7842 4378 7898 4380
rect 7922 4378 7978 4380
rect 8002 4378 8058 4380
rect 7762 4326 7808 4378
rect 7808 4326 7818 4378
rect 7842 4326 7872 4378
rect 7872 4326 7884 4378
rect 7884 4326 7898 4378
rect 7922 4326 7936 4378
rect 7936 4326 7948 4378
rect 7948 4326 7978 4378
rect 8002 4326 8012 4378
rect 8012 4326 8058 4378
rect 7762 4324 7818 4326
rect 7842 4324 7898 4326
rect 7922 4324 7978 4326
rect 8002 4324 8058 4326
rect 7762 3290 7818 3292
rect 7842 3290 7898 3292
rect 7922 3290 7978 3292
rect 8002 3290 8058 3292
rect 7762 3238 7808 3290
rect 7808 3238 7818 3290
rect 7842 3238 7872 3290
rect 7872 3238 7884 3290
rect 7884 3238 7898 3290
rect 7922 3238 7936 3290
rect 7936 3238 7948 3290
rect 7948 3238 7978 3290
rect 8002 3238 8012 3290
rect 8012 3238 8058 3290
rect 7762 3236 7818 3238
rect 7842 3236 7898 3238
rect 7922 3236 7978 3238
rect 8002 3236 8058 3238
rect 6212 2746 6268 2748
rect 6292 2746 6348 2748
rect 6372 2746 6428 2748
rect 6452 2746 6508 2748
rect 6212 2694 6258 2746
rect 6258 2694 6268 2746
rect 6292 2694 6322 2746
rect 6322 2694 6334 2746
rect 6334 2694 6348 2746
rect 6372 2694 6386 2746
rect 6386 2694 6398 2746
rect 6398 2694 6428 2746
rect 6452 2694 6462 2746
rect 6462 2694 6508 2746
rect 6212 2692 6268 2694
rect 6292 2692 6348 2694
rect 6372 2692 6428 2694
rect 6452 2692 6508 2694
rect 4662 2202 4718 2204
rect 4742 2202 4798 2204
rect 4822 2202 4878 2204
rect 4902 2202 4958 2204
rect 4662 2150 4708 2202
rect 4708 2150 4718 2202
rect 4742 2150 4772 2202
rect 4772 2150 4784 2202
rect 4784 2150 4798 2202
rect 4822 2150 4836 2202
rect 4836 2150 4848 2202
rect 4848 2150 4878 2202
rect 4902 2150 4912 2202
rect 4912 2150 4958 2202
rect 4662 2148 4718 2150
rect 4742 2148 4798 2150
rect 4822 2148 4878 2150
rect 4902 2148 4958 2150
rect 6212 1658 6268 1660
rect 6292 1658 6348 1660
rect 6372 1658 6428 1660
rect 6452 1658 6508 1660
rect 6212 1606 6258 1658
rect 6258 1606 6268 1658
rect 6292 1606 6322 1658
rect 6322 1606 6334 1658
rect 6334 1606 6348 1658
rect 6372 1606 6386 1658
rect 6386 1606 6398 1658
rect 6398 1606 6428 1658
rect 6452 1606 6462 1658
rect 6462 1606 6508 1658
rect 6212 1604 6268 1606
rect 6292 1604 6348 1606
rect 6372 1604 6428 1606
rect 6452 1604 6508 1606
rect 7762 2202 7818 2204
rect 7842 2202 7898 2204
rect 7922 2202 7978 2204
rect 8002 2202 8058 2204
rect 7762 2150 7808 2202
rect 7808 2150 7818 2202
rect 7842 2150 7872 2202
rect 7872 2150 7884 2202
rect 7884 2150 7898 2202
rect 7922 2150 7936 2202
rect 7936 2150 7948 2202
rect 7948 2150 7978 2202
rect 8002 2150 8012 2202
rect 8012 2150 8058 2202
rect 7762 2148 7818 2150
rect 7842 2148 7898 2150
rect 7922 2148 7978 2150
rect 8002 2148 8058 2150
rect 4662 1114 4718 1116
rect 4742 1114 4798 1116
rect 4822 1114 4878 1116
rect 4902 1114 4958 1116
rect 4662 1062 4708 1114
rect 4708 1062 4718 1114
rect 4742 1062 4772 1114
rect 4772 1062 4784 1114
rect 4784 1062 4798 1114
rect 4822 1062 4836 1114
rect 4836 1062 4848 1114
rect 4848 1062 4878 1114
rect 4902 1062 4912 1114
rect 4912 1062 4958 1114
rect 4662 1060 4718 1062
rect 4742 1060 4798 1062
rect 4822 1060 4878 1062
rect 4902 1060 4958 1062
rect 9312 14714 9368 14716
rect 9392 14714 9448 14716
rect 9472 14714 9528 14716
rect 9552 14714 9608 14716
rect 9312 14662 9358 14714
rect 9358 14662 9368 14714
rect 9392 14662 9422 14714
rect 9422 14662 9434 14714
rect 9434 14662 9448 14714
rect 9472 14662 9486 14714
rect 9486 14662 9498 14714
rect 9498 14662 9528 14714
rect 9552 14662 9562 14714
rect 9562 14662 9608 14714
rect 9312 14660 9368 14662
rect 9392 14660 9448 14662
rect 9472 14660 9528 14662
rect 9552 14660 9608 14662
rect 10862 16346 10918 16348
rect 10942 16346 10998 16348
rect 11022 16346 11078 16348
rect 11102 16346 11158 16348
rect 10862 16294 10908 16346
rect 10908 16294 10918 16346
rect 10942 16294 10972 16346
rect 10972 16294 10984 16346
rect 10984 16294 10998 16346
rect 11022 16294 11036 16346
rect 11036 16294 11048 16346
rect 11048 16294 11078 16346
rect 11102 16294 11112 16346
rect 11112 16294 11158 16346
rect 10862 16292 10918 16294
rect 10942 16292 10998 16294
rect 11022 16292 11078 16294
rect 11102 16292 11158 16294
rect 10862 15258 10918 15260
rect 10942 15258 10998 15260
rect 11022 15258 11078 15260
rect 11102 15258 11158 15260
rect 10862 15206 10908 15258
rect 10908 15206 10918 15258
rect 10942 15206 10972 15258
rect 10972 15206 10984 15258
rect 10984 15206 10998 15258
rect 11022 15206 11036 15258
rect 11036 15206 11048 15258
rect 11048 15206 11078 15258
rect 11102 15206 11112 15258
rect 11112 15206 11158 15258
rect 10862 15204 10918 15206
rect 10942 15204 10998 15206
rect 11022 15204 11078 15206
rect 11102 15204 11158 15206
rect 9312 13626 9368 13628
rect 9392 13626 9448 13628
rect 9472 13626 9528 13628
rect 9552 13626 9608 13628
rect 9312 13574 9358 13626
rect 9358 13574 9368 13626
rect 9392 13574 9422 13626
rect 9422 13574 9434 13626
rect 9434 13574 9448 13626
rect 9472 13574 9486 13626
rect 9486 13574 9498 13626
rect 9498 13574 9528 13626
rect 9552 13574 9562 13626
rect 9562 13574 9608 13626
rect 9312 13572 9368 13574
rect 9392 13572 9448 13574
rect 9472 13572 9528 13574
rect 9552 13572 9608 13574
rect 9312 12538 9368 12540
rect 9392 12538 9448 12540
rect 9472 12538 9528 12540
rect 9552 12538 9608 12540
rect 9312 12486 9358 12538
rect 9358 12486 9368 12538
rect 9392 12486 9422 12538
rect 9422 12486 9434 12538
rect 9434 12486 9448 12538
rect 9472 12486 9486 12538
rect 9486 12486 9498 12538
rect 9498 12486 9528 12538
rect 9552 12486 9562 12538
rect 9562 12486 9608 12538
rect 9312 12484 9368 12486
rect 9392 12484 9448 12486
rect 9472 12484 9528 12486
rect 9552 12484 9608 12486
rect 9312 11450 9368 11452
rect 9392 11450 9448 11452
rect 9472 11450 9528 11452
rect 9552 11450 9608 11452
rect 9312 11398 9358 11450
rect 9358 11398 9368 11450
rect 9392 11398 9422 11450
rect 9422 11398 9434 11450
rect 9434 11398 9448 11450
rect 9472 11398 9486 11450
rect 9486 11398 9498 11450
rect 9498 11398 9528 11450
rect 9552 11398 9562 11450
rect 9562 11398 9608 11450
rect 9312 11396 9368 11398
rect 9392 11396 9448 11398
rect 9472 11396 9528 11398
rect 9552 11396 9608 11398
rect 12412 17978 12468 17980
rect 12492 17978 12548 17980
rect 12572 17978 12628 17980
rect 12652 17978 12708 17980
rect 12412 17926 12458 17978
rect 12458 17926 12468 17978
rect 12492 17926 12522 17978
rect 12522 17926 12534 17978
rect 12534 17926 12548 17978
rect 12572 17926 12586 17978
rect 12586 17926 12598 17978
rect 12598 17926 12628 17978
rect 12652 17926 12662 17978
rect 12662 17926 12708 17978
rect 12412 17924 12468 17926
rect 12492 17924 12548 17926
rect 12572 17924 12628 17926
rect 12652 17924 12708 17926
rect 10862 14170 10918 14172
rect 10942 14170 10998 14172
rect 11022 14170 11078 14172
rect 11102 14170 11158 14172
rect 10862 14118 10908 14170
rect 10908 14118 10918 14170
rect 10942 14118 10972 14170
rect 10972 14118 10984 14170
rect 10984 14118 10998 14170
rect 11022 14118 11036 14170
rect 11036 14118 11048 14170
rect 11048 14118 11078 14170
rect 11102 14118 11112 14170
rect 11112 14118 11158 14170
rect 10862 14116 10918 14118
rect 10942 14116 10998 14118
rect 11022 14116 11078 14118
rect 11102 14116 11158 14118
rect 10862 13082 10918 13084
rect 10942 13082 10998 13084
rect 11022 13082 11078 13084
rect 11102 13082 11158 13084
rect 10862 13030 10908 13082
rect 10908 13030 10918 13082
rect 10942 13030 10972 13082
rect 10972 13030 10984 13082
rect 10984 13030 10998 13082
rect 11022 13030 11036 13082
rect 11036 13030 11048 13082
rect 11048 13030 11078 13082
rect 11102 13030 11112 13082
rect 11112 13030 11158 13082
rect 10862 13028 10918 13030
rect 10942 13028 10998 13030
rect 11022 13028 11078 13030
rect 11102 13028 11158 13030
rect 10862 11994 10918 11996
rect 10942 11994 10998 11996
rect 11022 11994 11078 11996
rect 11102 11994 11158 11996
rect 10862 11942 10908 11994
rect 10908 11942 10918 11994
rect 10942 11942 10972 11994
rect 10972 11942 10984 11994
rect 10984 11942 10998 11994
rect 11022 11942 11036 11994
rect 11036 11942 11048 11994
rect 11048 11942 11078 11994
rect 11102 11942 11112 11994
rect 11112 11942 11158 11994
rect 10862 11940 10918 11942
rect 10942 11940 10998 11942
rect 11022 11940 11078 11942
rect 11102 11940 11158 11942
rect 10862 10906 10918 10908
rect 10942 10906 10998 10908
rect 11022 10906 11078 10908
rect 11102 10906 11158 10908
rect 10862 10854 10908 10906
rect 10908 10854 10918 10906
rect 10942 10854 10972 10906
rect 10972 10854 10984 10906
rect 10984 10854 10998 10906
rect 11022 10854 11036 10906
rect 11036 10854 11048 10906
rect 11048 10854 11078 10906
rect 11102 10854 11112 10906
rect 11112 10854 11158 10906
rect 10862 10852 10918 10854
rect 10942 10852 10998 10854
rect 11022 10852 11078 10854
rect 11102 10852 11158 10854
rect 9312 10362 9368 10364
rect 9392 10362 9448 10364
rect 9472 10362 9528 10364
rect 9552 10362 9608 10364
rect 9312 10310 9358 10362
rect 9358 10310 9368 10362
rect 9392 10310 9422 10362
rect 9422 10310 9434 10362
rect 9434 10310 9448 10362
rect 9472 10310 9486 10362
rect 9486 10310 9498 10362
rect 9498 10310 9528 10362
rect 9552 10310 9562 10362
rect 9562 10310 9608 10362
rect 9312 10308 9368 10310
rect 9392 10308 9448 10310
rect 9472 10308 9528 10310
rect 9552 10308 9608 10310
rect 9312 9274 9368 9276
rect 9392 9274 9448 9276
rect 9472 9274 9528 9276
rect 9552 9274 9608 9276
rect 9312 9222 9358 9274
rect 9358 9222 9368 9274
rect 9392 9222 9422 9274
rect 9422 9222 9434 9274
rect 9434 9222 9448 9274
rect 9472 9222 9486 9274
rect 9486 9222 9498 9274
rect 9498 9222 9528 9274
rect 9552 9222 9562 9274
rect 9562 9222 9608 9274
rect 9312 9220 9368 9222
rect 9392 9220 9448 9222
rect 9472 9220 9528 9222
rect 9552 9220 9608 9222
rect 12412 16890 12468 16892
rect 12492 16890 12548 16892
rect 12572 16890 12628 16892
rect 12652 16890 12708 16892
rect 12412 16838 12458 16890
rect 12458 16838 12468 16890
rect 12492 16838 12522 16890
rect 12522 16838 12534 16890
rect 12534 16838 12548 16890
rect 12572 16838 12586 16890
rect 12586 16838 12598 16890
rect 12598 16838 12628 16890
rect 12652 16838 12662 16890
rect 12662 16838 12708 16890
rect 12412 16836 12468 16838
rect 12492 16836 12548 16838
rect 12572 16836 12628 16838
rect 12652 16836 12708 16838
rect 13962 18522 14018 18524
rect 14042 18522 14098 18524
rect 14122 18522 14178 18524
rect 14202 18522 14258 18524
rect 13962 18470 14008 18522
rect 14008 18470 14018 18522
rect 14042 18470 14072 18522
rect 14072 18470 14084 18522
rect 14084 18470 14098 18522
rect 14122 18470 14136 18522
rect 14136 18470 14148 18522
rect 14148 18470 14178 18522
rect 14202 18470 14212 18522
rect 14212 18470 14258 18522
rect 13962 18468 14018 18470
rect 14042 18468 14098 18470
rect 14122 18468 14178 18470
rect 14202 18468 14258 18470
rect 12412 15802 12468 15804
rect 12492 15802 12548 15804
rect 12572 15802 12628 15804
rect 12652 15802 12708 15804
rect 12412 15750 12458 15802
rect 12458 15750 12468 15802
rect 12492 15750 12522 15802
rect 12522 15750 12534 15802
rect 12534 15750 12548 15802
rect 12572 15750 12586 15802
rect 12586 15750 12598 15802
rect 12598 15750 12628 15802
rect 12652 15750 12662 15802
rect 12662 15750 12708 15802
rect 12412 15748 12468 15750
rect 12492 15748 12548 15750
rect 12572 15748 12628 15750
rect 12652 15748 12708 15750
rect 12412 14714 12468 14716
rect 12492 14714 12548 14716
rect 12572 14714 12628 14716
rect 12652 14714 12708 14716
rect 12412 14662 12458 14714
rect 12458 14662 12468 14714
rect 12492 14662 12522 14714
rect 12522 14662 12534 14714
rect 12534 14662 12548 14714
rect 12572 14662 12586 14714
rect 12586 14662 12598 14714
rect 12598 14662 12628 14714
rect 12652 14662 12662 14714
rect 12662 14662 12708 14714
rect 12412 14660 12468 14662
rect 12492 14660 12548 14662
rect 12572 14660 12628 14662
rect 12652 14660 12708 14662
rect 12412 13626 12468 13628
rect 12492 13626 12548 13628
rect 12572 13626 12628 13628
rect 12652 13626 12708 13628
rect 12412 13574 12458 13626
rect 12458 13574 12468 13626
rect 12492 13574 12522 13626
rect 12522 13574 12534 13626
rect 12534 13574 12548 13626
rect 12572 13574 12586 13626
rect 12586 13574 12598 13626
rect 12598 13574 12628 13626
rect 12652 13574 12662 13626
rect 12662 13574 12708 13626
rect 12412 13572 12468 13574
rect 12492 13572 12548 13574
rect 12572 13572 12628 13574
rect 12652 13572 12708 13574
rect 13962 17434 14018 17436
rect 14042 17434 14098 17436
rect 14122 17434 14178 17436
rect 14202 17434 14258 17436
rect 13962 17382 14008 17434
rect 14008 17382 14018 17434
rect 14042 17382 14072 17434
rect 14072 17382 14084 17434
rect 14084 17382 14098 17434
rect 14122 17382 14136 17434
rect 14136 17382 14148 17434
rect 14148 17382 14178 17434
rect 14202 17382 14212 17434
rect 14212 17382 14258 17434
rect 13962 17380 14018 17382
rect 14042 17380 14098 17382
rect 14122 17380 14178 17382
rect 14202 17380 14258 17382
rect 13962 16346 14018 16348
rect 14042 16346 14098 16348
rect 14122 16346 14178 16348
rect 14202 16346 14258 16348
rect 13962 16294 14008 16346
rect 14008 16294 14018 16346
rect 14042 16294 14072 16346
rect 14072 16294 14084 16346
rect 14084 16294 14098 16346
rect 14122 16294 14136 16346
rect 14136 16294 14148 16346
rect 14148 16294 14178 16346
rect 14202 16294 14212 16346
rect 14212 16294 14258 16346
rect 13962 16292 14018 16294
rect 14042 16292 14098 16294
rect 14122 16292 14178 16294
rect 14202 16292 14258 16294
rect 13962 15258 14018 15260
rect 14042 15258 14098 15260
rect 14122 15258 14178 15260
rect 14202 15258 14258 15260
rect 13962 15206 14008 15258
rect 14008 15206 14018 15258
rect 14042 15206 14072 15258
rect 14072 15206 14084 15258
rect 14084 15206 14098 15258
rect 14122 15206 14136 15258
rect 14136 15206 14148 15258
rect 14148 15206 14178 15258
rect 14202 15206 14212 15258
rect 14212 15206 14258 15258
rect 13962 15204 14018 15206
rect 14042 15204 14098 15206
rect 14122 15204 14178 15206
rect 14202 15204 14258 15206
rect 13962 14170 14018 14172
rect 14042 14170 14098 14172
rect 14122 14170 14178 14172
rect 14202 14170 14258 14172
rect 13962 14118 14008 14170
rect 14008 14118 14018 14170
rect 14042 14118 14072 14170
rect 14072 14118 14084 14170
rect 14084 14118 14098 14170
rect 14122 14118 14136 14170
rect 14136 14118 14148 14170
rect 14148 14118 14178 14170
rect 14202 14118 14212 14170
rect 14212 14118 14258 14170
rect 13962 14116 14018 14118
rect 14042 14116 14098 14118
rect 14122 14116 14178 14118
rect 14202 14116 14258 14118
rect 13962 13082 14018 13084
rect 14042 13082 14098 13084
rect 14122 13082 14178 13084
rect 14202 13082 14258 13084
rect 13962 13030 14008 13082
rect 14008 13030 14018 13082
rect 14042 13030 14072 13082
rect 14072 13030 14084 13082
rect 14084 13030 14098 13082
rect 14122 13030 14136 13082
rect 14136 13030 14148 13082
rect 14148 13030 14178 13082
rect 14202 13030 14212 13082
rect 14212 13030 14258 13082
rect 13962 13028 14018 13030
rect 14042 13028 14098 13030
rect 14122 13028 14178 13030
rect 14202 13028 14258 13030
rect 12412 12538 12468 12540
rect 12492 12538 12548 12540
rect 12572 12538 12628 12540
rect 12652 12538 12708 12540
rect 12412 12486 12458 12538
rect 12458 12486 12468 12538
rect 12492 12486 12522 12538
rect 12522 12486 12534 12538
rect 12534 12486 12548 12538
rect 12572 12486 12586 12538
rect 12586 12486 12598 12538
rect 12598 12486 12628 12538
rect 12652 12486 12662 12538
rect 12662 12486 12708 12538
rect 12412 12484 12468 12486
rect 12492 12484 12548 12486
rect 12572 12484 12628 12486
rect 12652 12484 12708 12486
rect 12412 11450 12468 11452
rect 12492 11450 12548 11452
rect 12572 11450 12628 11452
rect 12652 11450 12708 11452
rect 12412 11398 12458 11450
rect 12458 11398 12468 11450
rect 12492 11398 12522 11450
rect 12522 11398 12534 11450
rect 12534 11398 12548 11450
rect 12572 11398 12586 11450
rect 12586 11398 12598 11450
rect 12598 11398 12628 11450
rect 12652 11398 12662 11450
rect 12662 11398 12708 11450
rect 12412 11396 12468 11398
rect 12492 11396 12548 11398
rect 12572 11396 12628 11398
rect 12652 11396 12708 11398
rect 10862 9818 10918 9820
rect 10942 9818 10998 9820
rect 11022 9818 11078 9820
rect 11102 9818 11158 9820
rect 10862 9766 10908 9818
rect 10908 9766 10918 9818
rect 10942 9766 10972 9818
rect 10972 9766 10984 9818
rect 10984 9766 10998 9818
rect 11022 9766 11036 9818
rect 11036 9766 11048 9818
rect 11048 9766 11078 9818
rect 11102 9766 11112 9818
rect 11112 9766 11158 9818
rect 10862 9764 10918 9766
rect 10942 9764 10998 9766
rect 11022 9764 11078 9766
rect 11102 9764 11158 9766
rect 9312 8186 9368 8188
rect 9392 8186 9448 8188
rect 9472 8186 9528 8188
rect 9552 8186 9608 8188
rect 9312 8134 9358 8186
rect 9358 8134 9368 8186
rect 9392 8134 9422 8186
rect 9422 8134 9434 8186
rect 9434 8134 9448 8186
rect 9472 8134 9486 8186
rect 9486 8134 9498 8186
rect 9498 8134 9528 8186
rect 9552 8134 9562 8186
rect 9562 8134 9608 8186
rect 9312 8132 9368 8134
rect 9392 8132 9448 8134
rect 9472 8132 9528 8134
rect 9552 8132 9608 8134
rect 9312 7098 9368 7100
rect 9392 7098 9448 7100
rect 9472 7098 9528 7100
rect 9552 7098 9608 7100
rect 9312 7046 9358 7098
rect 9358 7046 9368 7098
rect 9392 7046 9422 7098
rect 9422 7046 9434 7098
rect 9434 7046 9448 7098
rect 9472 7046 9486 7098
rect 9486 7046 9498 7098
rect 9498 7046 9528 7098
rect 9552 7046 9562 7098
rect 9562 7046 9608 7098
rect 9312 7044 9368 7046
rect 9392 7044 9448 7046
rect 9472 7044 9528 7046
rect 9552 7044 9608 7046
rect 10862 8730 10918 8732
rect 10942 8730 10998 8732
rect 11022 8730 11078 8732
rect 11102 8730 11158 8732
rect 10862 8678 10908 8730
rect 10908 8678 10918 8730
rect 10942 8678 10972 8730
rect 10972 8678 10984 8730
rect 10984 8678 10998 8730
rect 11022 8678 11036 8730
rect 11036 8678 11048 8730
rect 11048 8678 11078 8730
rect 11102 8678 11112 8730
rect 11112 8678 11158 8730
rect 10862 8676 10918 8678
rect 10942 8676 10998 8678
rect 11022 8676 11078 8678
rect 11102 8676 11158 8678
rect 10862 7642 10918 7644
rect 10942 7642 10998 7644
rect 11022 7642 11078 7644
rect 11102 7642 11158 7644
rect 10862 7590 10908 7642
rect 10908 7590 10918 7642
rect 10942 7590 10972 7642
rect 10972 7590 10984 7642
rect 10984 7590 10998 7642
rect 11022 7590 11036 7642
rect 11036 7590 11048 7642
rect 11048 7590 11078 7642
rect 11102 7590 11112 7642
rect 11112 7590 11158 7642
rect 10862 7588 10918 7590
rect 10942 7588 10998 7590
rect 11022 7588 11078 7590
rect 11102 7588 11158 7590
rect 9312 6010 9368 6012
rect 9392 6010 9448 6012
rect 9472 6010 9528 6012
rect 9552 6010 9608 6012
rect 9312 5958 9358 6010
rect 9358 5958 9368 6010
rect 9392 5958 9422 6010
rect 9422 5958 9434 6010
rect 9434 5958 9448 6010
rect 9472 5958 9486 6010
rect 9486 5958 9498 6010
rect 9498 5958 9528 6010
rect 9552 5958 9562 6010
rect 9562 5958 9608 6010
rect 9312 5956 9368 5958
rect 9392 5956 9448 5958
rect 9472 5956 9528 5958
rect 9552 5956 9608 5958
rect 7762 1114 7818 1116
rect 7842 1114 7898 1116
rect 7922 1114 7978 1116
rect 8002 1114 8058 1116
rect 7762 1062 7808 1114
rect 7808 1062 7818 1114
rect 7842 1062 7872 1114
rect 7872 1062 7884 1114
rect 7884 1062 7898 1114
rect 7922 1062 7936 1114
rect 7936 1062 7948 1114
rect 7948 1062 7978 1114
rect 8002 1062 8012 1114
rect 8012 1062 8058 1114
rect 7762 1060 7818 1062
rect 7842 1060 7898 1062
rect 7922 1060 7978 1062
rect 8002 1060 8058 1062
rect 9312 4922 9368 4924
rect 9392 4922 9448 4924
rect 9472 4922 9528 4924
rect 9552 4922 9608 4924
rect 9312 4870 9358 4922
rect 9358 4870 9368 4922
rect 9392 4870 9422 4922
rect 9422 4870 9434 4922
rect 9434 4870 9448 4922
rect 9472 4870 9486 4922
rect 9486 4870 9498 4922
rect 9498 4870 9528 4922
rect 9552 4870 9562 4922
rect 9562 4870 9608 4922
rect 9312 4868 9368 4870
rect 9392 4868 9448 4870
rect 9472 4868 9528 4870
rect 9552 4868 9608 4870
rect 9312 3834 9368 3836
rect 9392 3834 9448 3836
rect 9472 3834 9528 3836
rect 9552 3834 9608 3836
rect 9312 3782 9358 3834
rect 9358 3782 9368 3834
rect 9392 3782 9422 3834
rect 9422 3782 9434 3834
rect 9434 3782 9448 3834
rect 9472 3782 9486 3834
rect 9486 3782 9498 3834
rect 9498 3782 9528 3834
rect 9552 3782 9562 3834
rect 9562 3782 9608 3834
rect 9312 3780 9368 3782
rect 9392 3780 9448 3782
rect 9472 3780 9528 3782
rect 9552 3780 9608 3782
rect 12412 10362 12468 10364
rect 12492 10362 12548 10364
rect 12572 10362 12628 10364
rect 12652 10362 12708 10364
rect 12412 10310 12458 10362
rect 12458 10310 12468 10362
rect 12492 10310 12522 10362
rect 12522 10310 12534 10362
rect 12534 10310 12548 10362
rect 12572 10310 12586 10362
rect 12586 10310 12598 10362
rect 12598 10310 12628 10362
rect 12652 10310 12662 10362
rect 12662 10310 12708 10362
rect 12412 10308 12468 10310
rect 12492 10308 12548 10310
rect 12572 10308 12628 10310
rect 12652 10308 12708 10310
rect 12412 9274 12468 9276
rect 12492 9274 12548 9276
rect 12572 9274 12628 9276
rect 12652 9274 12708 9276
rect 12412 9222 12458 9274
rect 12458 9222 12468 9274
rect 12492 9222 12522 9274
rect 12522 9222 12534 9274
rect 12534 9222 12548 9274
rect 12572 9222 12586 9274
rect 12586 9222 12598 9274
rect 12598 9222 12628 9274
rect 12652 9222 12662 9274
rect 12662 9222 12708 9274
rect 12412 9220 12468 9222
rect 12492 9220 12548 9222
rect 12572 9220 12628 9222
rect 12652 9220 12708 9222
rect 12412 8186 12468 8188
rect 12492 8186 12548 8188
rect 12572 8186 12628 8188
rect 12652 8186 12708 8188
rect 12412 8134 12458 8186
rect 12458 8134 12468 8186
rect 12492 8134 12522 8186
rect 12522 8134 12534 8186
rect 12534 8134 12548 8186
rect 12572 8134 12586 8186
rect 12586 8134 12598 8186
rect 12598 8134 12628 8186
rect 12652 8134 12662 8186
rect 12662 8134 12708 8186
rect 12412 8132 12468 8134
rect 12492 8132 12548 8134
rect 12572 8132 12628 8134
rect 12652 8132 12708 8134
rect 10862 6554 10918 6556
rect 10942 6554 10998 6556
rect 11022 6554 11078 6556
rect 11102 6554 11158 6556
rect 10862 6502 10908 6554
rect 10908 6502 10918 6554
rect 10942 6502 10972 6554
rect 10972 6502 10984 6554
rect 10984 6502 10998 6554
rect 11022 6502 11036 6554
rect 11036 6502 11048 6554
rect 11048 6502 11078 6554
rect 11102 6502 11112 6554
rect 11112 6502 11158 6554
rect 10862 6500 10918 6502
rect 10942 6500 10998 6502
rect 11022 6500 11078 6502
rect 11102 6500 11158 6502
rect 12412 7098 12468 7100
rect 12492 7098 12548 7100
rect 12572 7098 12628 7100
rect 12652 7098 12708 7100
rect 12412 7046 12458 7098
rect 12458 7046 12468 7098
rect 12492 7046 12522 7098
rect 12522 7046 12534 7098
rect 12534 7046 12548 7098
rect 12572 7046 12586 7098
rect 12586 7046 12598 7098
rect 12598 7046 12628 7098
rect 12652 7046 12662 7098
rect 12662 7046 12708 7098
rect 12412 7044 12468 7046
rect 12492 7044 12548 7046
rect 12572 7044 12628 7046
rect 12652 7044 12708 7046
rect 12412 6010 12468 6012
rect 12492 6010 12548 6012
rect 12572 6010 12628 6012
rect 12652 6010 12708 6012
rect 12412 5958 12458 6010
rect 12458 5958 12468 6010
rect 12492 5958 12522 6010
rect 12522 5958 12534 6010
rect 12534 5958 12548 6010
rect 12572 5958 12586 6010
rect 12586 5958 12598 6010
rect 12598 5958 12628 6010
rect 12652 5958 12662 6010
rect 12662 5958 12708 6010
rect 12412 5956 12468 5958
rect 12492 5956 12548 5958
rect 12572 5956 12628 5958
rect 12652 5956 12708 5958
rect 10862 5466 10918 5468
rect 10942 5466 10998 5468
rect 11022 5466 11078 5468
rect 11102 5466 11158 5468
rect 10862 5414 10908 5466
rect 10908 5414 10918 5466
rect 10942 5414 10972 5466
rect 10972 5414 10984 5466
rect 10984 5414 10998 5466
rect 11022 5414 11036 5466
rect 11036 5414 11048 5466
rect 11048 5414 11078 5466
rect 11102 5414 11112 5466
rect 11112 5414 11158 5466
rect 10862 5412 10918 5414
rect 10942 5412 10998 5414
rect 11022 5412 11078 5414
rect 11102 5412 11158 5414
rect 13962 11994 14018 11996
rect 14042 11994 14098 11996
rect 14122 11994 14178 11996
rect 14202 11994 14258 11996
rect 13962 11942 14008 11994
rect 14008 11942 14018 11994
rect 14042 11942 14072 11994
rect 14072 11942 14084 11994
rect 14084 11942 14098 11994
rect 14122 11942 14136 11994
rect 14136 11942 14148 11994
rect 14148 11942 14178 11994
rect 14202 11942 14212 11994
rect 14212 11942 14258 11994
rect 13962 11940 14018 11942
rect 14042 11940 14098 11942
rect 14122 11940 14178 11942
rect 14202 11940 14258 11942
rect 13962 10906 14018 10908
rect 14042 10906 14098 10908
rect 14122 10906 14178 10908
rect 14202 10906 14258 10908
rect 13962 10854 14008 10906
rect 14008 10854 14018 10906
rect 14042 10854 14072 10906
rect 14072 10854 14084 10906
rect 14084 10854 14098 10906
rect 14122 10854 14136 10906
rect 14136 10854 14148 10906
rect 14148 10854 14178 10906
rect 14202 10854 14212 10906
rect 14212 10854 14258 10906
rect 13962 10852 14018 10854
rect 14042 10852 14098 10854
rect 14122 10852 14178 10854
rect 14202 10852 14258 10854
rect 13962 9818 14018 9820
rect 14042 9818 14098 9820
rect 14122 9818 14178 9820
rect 14202 9818 14258 9820
rect 13962 9766 14008 9818
rect 14008 9766 14018 9818
rect 14042 9766 14072 9818
rect 14072 9766 14084 9818
rect 14084 9766 14098 9818
rect 14122 9766 14136 9818
rect 14136 9766 14148 9818
rect 14148 9766 14178 9818
rect 14202 9766 14212 9818
rect 14212 9766 14258 9818
rect 13962 9764 14018 9766
rect 14042 9764 14098 9766
rect 14122 9764 14178 9766
rect 14202 9764 14258 9766
rect 13962 8730 14018 8732
rect 14042 8730 14098 8732
rect 14122 8730 14178 8732
rect 14202 8730 14258 8732
rect 13962 8678 14008 8730
rect 14008 8678 14018 8730
rect 14042 8678 14072 8730
rect 14072 8678 14084 8730
rect 14084 8678 14098 8730
rect 14122 8678 14136 8730
rect 14136 8678 14148 8730
rect 14148 8678 14178 8730
rect 14202 8678 14212 8730
rect 14212 8678 14258 8730
rect 13962 8676 14018 8678
rect 14042 8676 14098 8678
rect 14122 8676 14178 8678
rect 14202 8676 14258 8678
rect 13962 7642 14018 7644
rect 14042 7642 14098 7644
rect 14122 7642 14178 7644
rect 14202 7642 14258 7644
rect 13962 7590 14008 7642
rect 14008 7590 14018 7642
rect 14042 7590 14072 7642
rect 14072 7590 14084 7642
rect 14084 7590 14098 7642
rect 14122 7590 14136 7642
rect 14136 7590 14148 7642
rect 14148 7590 14178 7642
rect 14202 7590 14212 7642
rect 14212 7590 14258 7642
rect 13962 7588 14018 7590
rect 14042 7588 14098 7590
rect 14122 7588 14178 7590
rect 14202 7588 14258 7590
rect 13962 6554 14018 6556
rect 14042 6554 14098 6556
rect 14122 6554 14178 6556
rect 14202 6554 14258 6556
rect 13962 6502 14008 6554
rect 14008 6502 14018 6554
rect 14042 6502 14072 6554
rect 14072 6502 14084 6554
rect 14084 6502 14098 6554
rect 14122 6502 14136 6554
rect 14136 6502 14148 6554
rect 14148 6502 14178 6554
rect 14202 6502 14212 6554
rect 14212 6502 14258 6554
rect 13962 6500 14018 6502
rect 14042 6500 14098 6502
rect 14122 6500 14178 6502
rect 14202 6500 14258 6502
rect 10862 4378 10918 4380
rect 10942 4378 10998 4380
rect 11022 4378 11078 4380
rect 11102 4378 11158 4380
rect 10862 4326 10908 4378
rect 10908 4326 10918 4378
rect 10942 4326 10972 4378
rect 10972 4326 10984 4378
rect 10984 4326 10998 4378
rect 11022 4326 11036 4378
rect 11036 4326 11048 4378
rect 11048 4326 11078 4378
rect 11102 4326 11112 4378
rect 11112 4326 11158 4378
rect 10862 4324 10918 4326
rect 10942 4324 10998 4326
rect 11022 4324 11078 4326
rect 11102 4324 11158 4326
rect 10862 3290 10918 3292
rect 10942 3290 10998 3292
rect 11022 3290 11078 3292
rect 11102 3290 11158 3292
rect 10862 3238 10908 3290
rect 10908 3238 10918 3290
rect 10942 3238 10972 3290
rect 10972 3238 10984 3290
rect 10984 3238 10998 3290
rect 11022 3238 11036 3290
rect 11036 3238 11048 3290
rect 11048 3238 11078 3290
rect 11102 3238 11112 3290
rect 11112 3238 11158 3290
rect 10862 3236 10918 3238
rect 10942 3236 10998 3238
rect 11022 3236 11078 3238
rect 11102 3236 11158 3238
rect 9312 2746 9368 2748
rect 9392 2746 9448 2748
rect 9472 2746 9528 2748
rect 9552 2746 9608 2748
rect 9312 2694 9358 2746
rect 9358 2694 9368 2746
rect 9392 2694 9422 2746
rect 9422 2694 9434 2746
rect 9434 2694 9448 2746
rect 9472 2694 9486 2746
rect 9486 2694 9498 2746
rect 9498 2694 9528 2746
rect 9552 2694 9562 2746
rect 9562 2694 9608 2746
rect 9312 2692 9368 2694
rect 9392 2692 9448 2694
rect 9472 2692 9528 2694
rect 9552 2692 9608 2694
rect 10862 2202 10918 2204
rect 10942 2202 10998 2204
rect 11022 2202 11078 2204
rect 11102 2202 11158 2204
rect 10862 2150 10908 2202
rect 10908 2150 10918 2202
rect 10942 2150 10972 2202
rect 10972 2150 10984 2202
rect 10984 2150 10998 2202
rect 11022 2150 11036 2202
rect 11036 2150 11048 2202
rect 11048 2150 11078 2202
rect 11102 2150 11112 2202
rect 11112 2150 11158 2202
rect 10862 2148 10918 2150
rect 10942 2148 10998 2150
rect 11022 2148 11078 2150
rect 11102 2148 11158 2150
rect 9312 1658 9368 1660
rect 9392 1658 9448 1660
rect 9472 1658 9528 1660
rect 9552 1658 9608 1660
rect 9312 1606 9358 1658
rect 9358 1606 9368 1658
rect 9392 1606 9422 1658
rect 9422 1606 9434 1658
rect 9434 1606 9448 1658
rect 9472 1606 9486 1658
rect 9486 1606 9498 1658
rect 9498 1606 9528 1658
rect 9552 1606 9562 1658
rect 9562 1606 9608 1658
rect 9312 1604 9368 1606
rect 9392 1604 9448 1606
rect 9472 1604 9528 1606
rect 9552 1604 9608 1606
rect 12412 4922 12468 4924
rect 12492 4922 12548 4924
rect 12572 4922 12628 4924
rect 12652 4922 12708 4924
rect 12412 4870 12458 4922
rect 12458 4870 12468 4922
rect 12492 4870 12522 4922
rect 12522 4870 12534 4922
rect 12534 4870 12548 4922
rect 12572 4870 12586 4922
rect 12586 4870 12598 4922
rect 12598 4870 12628 4922
rect 12652 4870 12662 4922
rect 12662 4870 12708 4922
rect 12412 4868 12468 4870
rect 12492 4868 12548 4870
rect 12572 4868 12628 4870
rect 12652 4868 12708 4870
rect 12412 3834 12468 3836
rect 12492 3834 12548 3836
rect 12572 3834 12628 3836
rect 12652 3834 12708 3836
rect 12412 3782 12458 3834
rect 12458 3782 12468 3834
rect 12492 3782 12522 3834
rect 12522 3782 12534 3834
rect 12534 3782 12548 3834
rect 12572 3782 12586 3834
rect 12586 3782 12598 3834
rect 12598 3782 12628 3834
rect 12652 3782 12662 3834
rect 12662 3782 12708 3834
rect 12412 3780 12468 3782
rect 12492 3780 12548 3782
rect 12572 3780 12628 3782
rect 12652 3780 12708 3782
rect 13962 5466 14018 5468
rect 14042 5466 14098 5468
rect 14122 5466 14178 5468
rect 14202 5466 14258 5468
rect 13962 5414 14008 5466
rect 14008 5414 14018 5466
rect 14042 5414 14072 5466
rect 14072 5414 14084 5466
rect 14084 5414 14098 5466
rect 14122 5414 14136 5466
rect 14136 5414 14148 5466
rect 14148 5414 14178 5466
rect 14202 5414 14212 5466
rect 14212 5414 14258 5466
rect 13962 5412 14018 5414
rect 14042 5412 14098 5414
rect 14122 5412 14178 5414
rect 14202 5412 14258 5414
rect 13962 4378 14018 4380
rect 14042 4378 14098 4380
rect 14122 4378 14178 4380
rect 14202 4378 14258 4380
rect 13962 4326 14008 4378
rect 14008 4326 14018 4378
rect 14042 4326 14072 4378
rect 14072 4326 14084 4378
rect 14084 4326 14098 4378
rect 14122 4326 14136 4378
rect 14136 4326 14148 4378
rect 14148 4326 14178 4378
rect 14202 4326 14212 4378
rect 14212 4326 14258 4378
rect 13962 4324 14018 4326
rect 14042 4324 14098 4326
rect 14122 4324 14178 4326
rect 14202 4324 14258 4326
rect 18418 18536 18474 18592
rect 17062 18522 17118 18524
rect 17142 18522 17198 18524
rect 17222 18522 17278 18524
rect 17302 18522 17358 18524
rect 17062 18470 17108 18522
rect 17108 18470 17118 18522
rect 17142 18470 17172 18522
rect 17172 18470 17184 18522
rect 17184 18470 17198 18522
rect 17222 18470 17236 18522
rect 17236 18470 17248 18522
rect 17248 18470 17278 18522
rect 17302 18470 17312 18522
rect 17312 18470 17358 18522
rect 17062 18468 17118 18470
rect 17142 18468 17198 18470
rect 17222 18468 17278 18470
rect 17302 18468 17358 18470
rect 15512 17978 15568 17980
rect 15592 17978 15648 17980
rect 15672 17978 15728 17980
rect 15752 17978 15808 17980
rect 15512 17926 15558 17978
rect 15558 17926 15568 17978
rect 15592 17926 15622 17978
rect 15622 17926 15634 17978
rect 15634 17926 15648 17978
rect 15672 17926 15686 17978
rect 15686 17926 15698 17978
rect 15698 17926 15728 17978
rect 15752 17926 15762 17978
rect 15762 17926 15808 17978
rect 15512 17924 15568 17926
rect 15592 17924 15648 17926
rect 15672 17924 15728 17926
rect 15752 17924 15808 17926
rect 15512 16890 15568 16892
rect 15592 16890 15648 16892
rect 15672 16890 15728 16892
rect 15752 16890 15808 16892
rect 15512 16838 15558 16890
rect 15558 16838 15568 16890
rect 15592 16838 15622 16890
rect 15622 16838 15634 16890
rect 15634 16838 15648 16890
rect 15672 16838 15686 16890
rect 15686 16838 15698 16890
rect 15698 16838 15728 16890
rect 15752 16838 15762 16890
rect 15762 16838 15808 16890
rect 15512 16836 15568 16838
rect 15592 16836 15648 16838
rect 15672 16836 15728 16838
rect 15752 16836 15808 16838
rect 15512 15802 15568 15804
rect 15592 15802 15648 15804
rect 15672 15802 15728 15804
rect 15752 15802 15808 15804
rect 15512 15750 15558 15802
rect 15558 15750 15568 15802
rect 15592 15750 15622 15802
rect 15622 15750 15634 15802
rect 15634 15750 15648 15802
rect 15672 15750 15686 15802
rect 15686 15750 15698 15802
rect 15698 15750 15728 15802
rect 15752 15750 15762 15802
rect 15762 15750 15808 15802
rect 15512 15748 15568 15750
rect 15592 15748 15648 15750
rect 15672 15748 15728 15750
rect 15752 15748 15808 15750
rect 15512 14714 15568 14716
rect 15592 14714 15648 14716
rect 15672 14714 15728 14716
rect 15752 14714 15808 14716
rect 15512 14662 15558 14714
rect 15558 14662 15568 14714
rect 15592 14662 15622 14714
rect 15622 14662 15634 14714
rect 15634 14662 15648 14714
rect 15672 14662 15686 14714
rect 15686 14662 15698 14714
rect 15698 14662 15728 14714
rect 15752 14662 15762 14714
rect 15762 14662 15808 14714
rect 15512 14660 15568 14662
rect 15592 14660 15648 14662
rect 15672 14660 15728 14662
rect 15752 14660 15808 14662
rect 17062 17434 17118 17436
rect 17142 17434 17198 17436
rect 17222 17434 17278 17436
rect 17302 17434 17358 17436
rect 17062 17382 17108 17434
rect 17108 17382 17118 17434
rect 17142 17382 17172 17434
rect 17172 17382 17184 17434
rect 17184 17382 17198 17434
rect 17222 17382 17236 17434
rect 17236 17382 17248 17434
rect 17248 17382 17278 17434
rect 17302 17382 17312 17434
rect 17312 17382 17358 17434
rect 17062 17380 17118 17382
rect 17142 17380 17198 17382
rect 17222 17380 17278 17382
rect 17302 17380 17358 17382
rect 17062 16346 17118 16348
rect 17142 16346 17198 16348
rect 17222 16346 17278 16348
rect 17302 16346 17358 16348
rect 17062 16294 17108 16346
rect 17108 16294 17118 16346
rect 17142 16294 17172 16346
rect 17172 16294 17184 16346
rect 17184 16294 17198 16346
rect 17222 16294 17236 16346
rect 17236 16294 17248 16346
rect 17248 16294 17278 16346
rect 17302 16294 17312 16346
rect 17312 16294 17358 16346
rect 17062 16292 17118 16294
rect 17142 16292 17198 16294
rect 17222 16292 17278 16294
rect 17302 16292 17358 16294
rect 15512 13626 15568 13628
rect 15592 13626 15648 13628
rect 15672 13626 15728 13628
rect 15752 13626 15808 13628
rect 15512 13574 15558 13626
rect 15558 13574 15568 13626
rect 15592 13574 15622 13626
rect 15622 13574 15634 13626
rect 15634 13574 15648 13626
rect 15672 13574 15686 13626
rect 15686 13574 15698 13626
rect 15698 13574 15728 13626
rect 15752 13574 15762 13626
rect 15762 13574 15808 13626
rect 15512 13572 15568 13574
rect 15592 13572 15648 13574
rect 15672 13572 15728 13574
rect 15752 13572 15808 13574
rect 17062 15258 17118 15260
rect 17142 15258 17198 15260
rect 17222 15258 17278 15260
rect 17302 15258 17358 15260
rect 17062 15206 17108 15258
rect 17108 15206 17118 15258
rect 17142 15206 17172 15258
rect 17172 15206 17184 15258
rect 17184 15206 17198 15258
rect 17222 15206 17236 15258
rect 17236 15206 17248 15258
rect 17248 15206 17278 15258
rect 17302 15206 17312 15258
rect 17312 15206 17358 15258
rect 17062 15204 17118 15206
rect 17142 15204 17198 15206
rect 17222 15204 17278 15206
rect 17302 15204 17358 15206
rect 17062 14170 17118 14172
rect 17142 14170 17198 14172
rect 17222 14170 17278 14172
rect 17302 14170 17358 14172
rect 17062 14118 17108 14170
rect 17108 14118 17118 14170
rect 17142 14118 17172 14170
rect 17172 14118 17184 14170
rect 17184 14118 17198 14170
rect 17222 14118 17236 14170
rect 17236 14118 17248 14170
rect 17248 14118 17278 14170
rect 17302 14118 17312 14170
rect 17312 14118 17358 14170
rect 17062 14116 17118 14118
rect 17142 14116 17198 14118
rect 17222 14116 17278 14118
rect 17302 14116 17358 14118
rect 15512 12538 15568 12540
rect 15592 12538 15648 12540
rect 15672 12538 15728 12540
rect 15752 12538 15808 12540
rect 15512 12486 15558 12538
rect 15558 12486 15568 12538
rect 15592 12486 15622 12538
rect 15622 12486 15634 12538
rect 15634 12486 15648 12538
rect 15672 12486 15686 12538
rect 15686 12486 15698 12538
rect 15698 12486 15728 12538
rect 15752 12486 15762 12538
rect 15762 12486 15808 12538
rect 15512 12484 15568 12486
rect 15592 12484 15648 12486
rect 15672 12484 15728 12486
rect 15752 12484 15808 12486
rect 15512 11450 15568 11452
rect 15592 11450 15648 11452
rect 15672 11450 15728 11452
rect 15752 11450 15808 11452
rect 15512 11398 15558 11450
rect 15558 11398 15568 11450
rect 15592 11398 15622 11450
rect 15622 11398 15634 11450
rect 15634 11398 15648 11450
rect 15672 11398 15686 11450
rect 15686 11398 15698 11450
rect 15698 11398 15728 11450
rect 15752 11398 15762 11450
rect 15762 11398 15808 11450
rect 15512 11396 15568 11398
rect 15592 11396 15648 11398
rect 15672 11396 15728 11398
rect 15752 11396 15808 11398
rect 15512 10362 15568 10364
rect 15592 10362 15648 10364
rect 15672 10362 15728 10364
rect 15752 10362 15808 10364
rect 15512 10310 15558 10362
rect 15558 10310 15568 10362
rect 15592 10310 15622 10362
rect 15622 10310 15634 10362
rect 15634 10310 15648 10362
rect 15672 10310 15686 10362
rect 15686 10310 15698 10362
rect 15698 10310 15728 10362
rect 15752 10310 15762 10362
rect 15762 10310 15808 10362
rect 15512 10308 15568 10310
rect 15592 10308 15648 10310
rect 15672 10308 15728 10310
rect 15752 10308 15808 10310
rect 15512 9274 15568 9276
rect 15592 9274 15648 9276
rect 15672 9274 15728 9276
rect 15752 9274 15808 9276
rect 15512 9222 15558 9274
rect 15558 9222 15568 9274
rect 15592 9222 15622 9274
rect 15622 9222 15634 9274
rect 15634 9222 15648 9274
rect 15672 9222 15686 9274
rect 15686 9222 15698 9274
rect 15698 9222 15728 9274
rect 15752 9222 15762 9274
rect 15762 9222 15808 9274
rect 15512 9220 15568 9222
rect 15592 9220 15648 9222
rect 15672 9220 15728 9222
rect 15752 9220 15808 9222
rect 15512 8186 15568 8188
rect 15592 8186 15648 8188
rect 15672 8186 15728 8188
rect 15752 8186 15808 8188
rect 15512 8134 15558 8186
rect 15558 8134 15568 8186
rect 15592 8134 15622 8186
rect 15622 8134 15634 8186
rect 15634 8134 15648 8186
rect 15672 8134 15686 8186
rect 15686 8134 15698 8186
rect 15698 8134 15728 8186
rect 15752 8134 15762 8186
rect 15762 8134 15808 8186
rect 15512 8132 15568 8134
rect 15592 8132 15648 8134
rect 15672 8132 15728 8134
rect 15752 8132 15808 8134
rect 15512 7098 15568 7100
rect 15592 7098 15648 7100
rect 15672 7098 15728 7100
rect 15752 7098 15808 7100
rect 15512 7046 15558 7098
rect 15558 7046 15568 7098
rect 15592 7046 15622 7098
rect 15622 7046 15634 7098
rect 15634 7046 15648 7098
rect 15672 7046 15686 7098
rect 15686 7046 15698 7098
rect 15698 7046 15728 7098
rect 15752 7046 15762 7098
rect 15762 7046 15808 7098
rect 15512 7044 15568 7046
rect 15592 7044 15648 7046
rect 15672 7044 15728 7046
rect 15752 7044 15808 7046
rect 15512 6010 15568 6012
rect 15592 6010 15648 6012
rect 15672 6010 15728 6012
rect 15752 6010 15808 6012
rect 15512 5958 15558 6010
rect 15558 5958 15568 6010
rect 15592 5958 15622 6010
rect 15622 5958 15634 6010
rect 15634 5958 15648 6010
rect 15672 5958 15686 6010
rect 15686 5958 15698 6010
rect 15698 5958 15728 6010
rect 15752 5958 15762 6010
rect 15762 5958 15808 6010
rect 15512 5956 15568 5958
rect 15592 5956 15648 5958
rect 15672 5956 15728 5958
rect 15752 5956 15808 5958
rect 13962 3290 14018 3292
rect 14042 3290 14098 3292
rect 14122 3290 14178 3292
rect 14202 3290 14258 3292
rect 13962 3238 14008 3290
rect 14008 3238 14018 3290
rect 14042 3238 14072 3290
rect 14072 3238 14084 3290
rect 14084 3238 14098 3290
rect 14122 3238 14136 3290
rect 14136 3238 14148 3290
rect 14148 3238 14178 3290
rect 14202 3238 14212 3290
rect 14212 3238 14258 3290
rect 13962 3236 14018 3238
rect 14042 3236 14098 3238
rect 14122 3236 14178 3238
rect 14202 3236 14258 3238
rect 12412 2746 12468 2748
rect 12492 2746 12548 2748
rect 12572 2746 12628 2748
rect 12652 2746 12708 2748
rect 12412 2694 12458 2746
rect 12458 2694 12468 2746
rect 12492 2694 12522 2746
rect 12522 2694 12534 2746
rect 12534 2694 12548 2746
rect 12572 2694 12586 2746
rect 12586 2694 12598 2746
rect 12598 2694 12628 2746
rect 12652 2694 12662 2746
rect 12662 2694 12708 2746
rect 12412 2692 12468 2694
rect 12492 2692 12548 2694
rect 12572 2692 12628 2694
rect 12652 2692 12708 2694
rect 12412 1658 12468 1660
rect 12492 1658 12548 1660
rect 12572 1658 12628 1660
rect 12652 1658 12708 1660
rect 12412 1606 12458 1658
rect 12458 1606 12468 1658
rect 12492 1606 12522 1658
rect 12522 1606 12534 1658
rect 12534 1606 12548 1658
rect 12572 1606 12586 1658
rect 12586 1606 12598 1658
rect 12598 1606 12628 1658
rect 12652 1606 12662 1658
rect 12662 1606 12708 1658
rect 12412 1604 12468 1606
rect 12492 1604 12548 1606
rect 12572 1604 12628 1606
rect 12652 1604 12708 1606
rect 17062 13082 17118 13084
rect 17142 13082 17198 13084
rect 17222 13082 17278 13084
rect 17302 13082 17358 13084
rect 17062 13030 17108 13082
rect 17108 13030 17118 13082
rect 17142 13030 17172 13082
rect 17172 13030 17184 13082
rect 17184 13030 17198 13082
rect 17222 13030 17236 13082
rect 17236 13030 17248 13082
rect 17248 13030 17278 13082
rect 17302 13030 17312 13082
rect 17312 13030 17358 13082
rect 17062 13028 17118 13030
rect 17142 13028 17198 13030
rect 17222 13028 17278 13030
rect 17302 13028 17358 13030
rect 17062 11994 17118 11996
rect 17142 11994 17198 11996
rect 17222 11994 17278 11996
rect 17302 11994 17358 11996
rect 17062 11942 17108 11994
rect 17108 11942 17118 11994
rect 17142 11942 17172 11994
rect 17172 11942 17184 11994
rect 17184 11942 17198 11994
rect 17222 11942 17236 11994
rect 17236 11942 17248 11994
rect 17248 11942 17278 11994
rect 17302 11942 17312 11994
rect 17312 11942 17358 11994
rect 17062 11940 17118 11942
rect 17142 11940 17198 11942
rect 17222 11940 17278 11942
rect 17302 11940 17358 11942
rect 18418 16088 18474 16144
rect 17062 10906 17118 10908
rect 17142 10906 17198 10908
rect 17222 10906 17278 10908
rect 17302 10906 17358 10908
rect 17062 10854 17108 10906
rect 17108 10854 17118 10906
rect 17142 10854 17172 10906
rect 17172 10854 17184 10906
rect 17184 10854 17198 10906
rect 17222 10854 17236 10906
rect 17236 10854 17248 10906
rect 17248 10854 17278 10906
rect 17302 10854 17312 10906
rect 17312 10854 17358 10906
rect 17062 10852 17118 10854
rect 17142 10852 17198 10854
rect 17222 10852 17278 10854
rect 17302 10852 17358 10854
rect 17062 9818 17118 9820
rect 17142 9818 17198 9820
rect 17222 9818 17278 9820
rect 17302 9818 17358 9820
rect 17062 9766 17108 9818
rect 17108 9766 17118 9818
rect 17142 9766 17172 9818
rect 17172 9766 17184 9818
rect 17184 9766 17198 9818
rect 17222 9766 17236 9818
rect 17236 9766 17248 9818
rect 17248 9766 17278 9818
rect 17302 9766 17312 9818
rect 17312 9766 17358 9818
rect 17062 9764 17118 9766
rect 17142 9764 17198 9766
rect 17222 9764 17278 9766
rect 17302 9764 17358 9766
rect 17062 8730 17118 8732
rect 17142 8730 17198 8732
rect 17222 8730 17278 8732
rect 17302 8730 17358 8732
rect 17062 8678 17108 8730
rect 17108 8678 17118 8730
rect 17142 8678 17172 8730
rect 17172 8678 17184 8730
rect 17184 8678 17198 8730
rect 17222 8678 17236 8730
rect 17236 8678 17248 8730
rect 17248 8678 17278 8730
rect 17302 8678 17312 8730
rect 17312 8678 17358 8730
rect 17062 8676 17118 8678
rect 17142 8676 17198 8678
rect 17222 8676 17278 8678
rect 17302 8676 17358 8678
rect 17062 7642 17118 7644
rect 17142 7642 17198 7644
rect 17222 7642 17278 7644
rect 17302 7642 17358 7644
rect 17062 7590 17108 7642
rect 17108 7590 17118 7642
rect 17142 7590 17172 7642
rect 17172 7590 17184 7642
rect 17184 7590 17198 7642
rect 17222 7590 17236 7642
rect 17236 7590 17248 7642
rect 17248 7590 17278 7642
rect 17302 7590 17312 7642
rect 17312 7590 17358 7642
rect 17062 7588 17118 7590
rect 17142 7588 17198 7590
rect 17222 7588 17278 7590
rect 17302 7588 17358 7590
rect 15512 4922 15568 4924
rect 15592 4922 15648 4924
rect 15672 4922 15728 4924
rect 15752 4922 15808 4924
rect 15512 4870 15558 4922
rect 15558 4870 15568 4922
rect 15592 4870 15622 4922
rect 15622 4870 15634 4922
rect 15634 4870 15648 4922
rect 15672 4870 15686 4922
rect 15686 4870 15698 4922
rect 15698 4870 15728 4922
rect 15752 4870 15762 4922
rect 15762 4870 15808 4922
rect 15512 4868 15568 4870
rect 15592 4868 15648 4870
rect 15672 4868 15728 4870
rect 15752 4868 15808 4870
rect 15512 3834 15568 3836
rect 15592 3834 15648 3836
rect 15672 3834 15728 3836
rect 15752 3834 15808 3836
rect 15512 3782 15558 3834
rect 15558 3782 15568 3834
rect 15592 3782 15622 3834
rect 15622 3782 15634 3834
rect 15634 3782 15648 3834
rect 15672 3782 15686 3834
rect 15686 3782 15698 3834
rect 15698 3782 15728 3834
rect 15752 3782 15762 3834
rect 15762 3782 15808 3834
rect 15512 3780 15568 3782
rect 15592 3780 15648 3782
rect 15672 3780 15728 3782
rect 15752 3780 15808 3782
rect 15512 2746 15568 2748
rect 15592 2746 15648 2748
rect 15672 2746 15728 2748
rect 15752 2746 15808 2748
rect 15512 2694 15558 2746
rect 15558 2694 15568 2746
rect 15592 2694 15622 2746
rect 15622 2694 15634 2746
rect 15634 2694 15648 2746
rect 15672 2694 15686 2746
rect 15686 2694 15698 2746
rect 15698 2694 15728 2746
rect 15752 2694 15762 2746
rect 15762 2694 15808 2746
rect 15512 2692 15568 2694
rect 15592 2692 15648 2694
rect 15672 2692 15728 2694
rect 15752 2692 15808 2694
rect 13962 2202 14018 2204
rect 14042 2202 14098 2204
rect 14122 2202 14178 2204
rect 14202 2202 14258 2204
rect 13962 2150 14008 2202
rect 14008 2150 14018 2202
rect 14042 2150 14072 2202
rect 14072 2150 14084 2202
rect 14084 2150 14098 2202
rect 14122 2150 14136 2202
rect 14136 2150 14148 2202
rect 14148 2150 14178 2202
rect 14202 2150 14212 2202
rect 14212 2150 14258 2202
rect 13962 2148 14018 2150
rect 14042 2148 14098 2150
rect 14122 2148 14178 2150
rect 14202 2148 14258 2150
rect 15512 1658 15568 1660
rect 15592 1658 15648 1660
rect 15672 1658 15728 1660
rect 15752 1658 15808 1660
rect 15512 1606 15558 1658
rect 15558 1606 15568 1658
rect 15592 1606 15622 1658
rect 15622 1606 15634 1658
rect 15634 1606 15648 1658
rect 15672 1606 15686 1658
rect 15686 1606 15698 1658
rect 15698 1606 15728 1658
rect 15752 1606 15762 1658
rect 15762 1606 15808 1658
rect 15512 1604 15568 1606
rect 15592 1604 15648 1606
rect 15672 1604 15728 1606
rect 15752 1604 15808 1606
rect 17062 6554 17118 6556
rect 17142 6554 17198 6556
rect 17222 6554 17278 6556
rect 17302 6554 17358 6556
rect 17062 6502 17108 6554
rect 17108 6502 17118 6554
rect 17142 6502 17172 6554
rect 17172 6502 17184 6554
rect 17184 6502 17198 6554
rect 17222 6502 17236 6554
rect 17236 6502 17248 6554
rect 17248 6502 17278 6554
rect 17302 6502 17312 6554
rect 17312 6502 17358 6554
rect 17062 6500 17118 6502
rect 17142 6500 17198 6502
rect 17222 6500 17278 6502
rect 17302 6500 17358 6502
rect 17062 5466 17118 5468
rect 17142 5466 17198 5468
rect 17222 5466 17278 5468
rect 17302 5466 17358 5468
rect 17062 5414 17108 5466
rect 17108 5414 17118 5466
rect 17142 5414 17172 5466
rect 17172 5414 17184 5466
rect 17184 5414 17198 5466
rect 17222 5414 17236 5466
rect 17236 5414 17248 5466
rect 17248 5414 17278 5466
rect 17302 5414 17312 5466
rect 17312 5414 17358 5466
rect 17062 5412 17118 5414
rect 17142 5412 17198 5414
rect 17222 5412 17278 5414
rect 17302 5412 17358 5414
rect 17062 4378 17118 4380
rect 17142 4378 17198 4380
rect 17222 4378 17278 4380
rect 17302 4378 17358 4380
rect 17062 4326 17108 4378
rect 17108 4326 17118 4378
rect 17142 4326 17172 4378
rect 17172 4326 17184 4378
rect 17184 4326 17198 4378
rect 17222 4326 17236 4378
rect 17236 4326 17248 4378
rect 17248 4326 17278 4378
rect 17302 4326 17312 4378
rect 17312 4326 17358 4378
rect 17062 4324 17118 4326
rect 17142 4324 17198 4326
rect 17222 4324 17278 4326
rect 17302 4324 17358 4326
rect 17062 3290 17118 3292
rect 17142 3290 17198 3292
rect 17222 3290 17278 3292
rect 17302 3290 17358 3292
rect 17062 3238 17108 3290
rect 17108 3238 17118 3290
rect 17142 3238 17172 3290
rect 17172 3238 17184 3290
rect 17184 3238 17198 3290
rect 17222 3238 17236 3290
rect 17236 3238 17248 3290
rect 17248 3238 17278 3290
rect 17302 3238 17312 3290
rect 17312 3238 17358 3290
rect 17062 3236 17118 3238
rect 17142 3236 17198 3238
rect 17222 3236 17278 3238
rect 17302 3236 17358 3238
rect 17062 2202 17118 2204
rect 17142 2202 17198 2204
rect 17222 2202 17278 2204
rect 17302 2202 17358 2204
rect 17062 2150 17108 2202
rect 17108 2150 17118 2202
rect 17142 2150 17172 2202
rect 17172 2150 17184 2202
rect 17184 2150 17198 2202
rect 17222 2150 17236 2202
rect 17236 2150 17248 2202
rect 17248 2150 17278 2202
rect 17302 2150 17312 2202
rect 17312 2150 17358 2202
rect 17062 2148 17118 2150
rect 17142 2148 17198 2150
rect 17222 2148 17278 2150
rect 17302 2148 17358 2150
rect 10862 1114 10918 1116
rect 10942 1114 10998 1116
rect 11022 1114 11078 1116
rect 11102 1114 11158 1116
rect 10862 1062 10908 1114
rect 10908 1062 10918 1114
rect 10942 1062 10972 1114
rect 10972 1062 10984 1114
rect 10984 1062 10998 1114
rect 11022 1062 11036 1114
rect 11036 1062 11048 1114
rect 11048 1062 11078 1114
rect 11102 1062 11112 1114
rect 11112 1062 11158 1114
rect 10862 1060 10918 1062
rect 10942 1060 10998 1062
rect 11022 1060 11078 1062
rect 11102 1060 11158 1062
rect 13962 1114 14018 1116
rect 14042 1114 14098 1116
rect 14122 1114 14178 1116
rect 14202 1114 14258 1116
rect 13962 1062 14008 1114
rect 14008 1062 14018 1114
rect 14042 1062 14072 1114
rect 14072 1062 14084 1114
rect 14084 1062 14098 1114
rect 14122 1062 14136 1114
rect 14136 1062 14148 1114
rect 14148 1062 14178 1114
rect 14202 1062 14212 1114
rect 14212 1062 14258 1114
rect 13962 1060 14018 1062
rect 14042 1060 14098 1062
rect 14122 1060 14178 1062
rect 14202 1060 14258 1062
rect 18612 17978 18668 17980
rect 18692 17978 18748 17980
rect 18772 17978 18828 17980
rect 18852 17978 18908 17980
rect 18612 17926 18658 17978
rect 18658 17926 18668 17978
rect 18692 17926 18722 17978
rect 18722 17926 18734 17978
rect 18734 17926 18748 17978
rect 18772 17926 18786 17978
rect 18786 17926 18798 17978
rect 18798 17926 18828 17978
rect 18852 17926 18862 17978
rect 18862 17926 18908 17978
rect 18612 17924 18668 17926
rect 18692 17924 18748 17926
rect 18772 17924 18828 17926
rect 18852 17924 18908 17926
rect 18612 16890 18668 16892
rect 18692 16890 18748 16892
rect 18772 16890 18828 16892
rect 18852 16890 18908 16892
rect 18612 16838 18658 16890
rect 18658 16838 18668 16890
rect 18692 16838 18722 16890
rect 18722 16838 18734 16890
rect 18734 16838 18748 16890
rect 18772 16838 18786 16890
rect 18786 16838 18798 16890
rect 18798 16838 18828 16890
rect 18852 16838 18862 16890
rect 18862 16838 18908 16890
rect 18612 16836 18668 16838
rect 18692 16836 18748 16838
rect 18772 16836 18828 16838
rect 18852 16836 18908 16838
rect 18612 15802 18668 15804
rect 18692 15802 18748 15804
rect 18772 15802 18828 15804
rect 18852 15802 18908 15804
rect 18612 15750 18658 15802
rect 18658 15750 18668 15802
rect 18692 15750 18722 15802
rect 18722 15750 18734 15802
rect 18734 15750 18748 15802
rect 18772 15750 18786 15802
rect 18786 15750 18798 15802
rect 18798 15750 18828 15802
rect 18852 15750 18862 15802
rect 18862 15750 18908 15802
rect 18612 15748 18668 15750
rect 18692 15748 18748 15750
rect 18772 15748 18828 15750
rect 18852 15748 18908 15750
rect 18612 14714 18668 14716
rect 18692 14714 18748 14716
rect 18772 14714 18828 14716
rect 18852 14714 18908 14716
rect 18612 14662 18658 14714
rect 18658 14662 18668 14714
rect 18692 14662 18722 14714
rect 18722 14662 18734 14714
rect 18734 14662 18748 14714
rect 18772 14662 18786 14714
rect 18786 14662 18798 14714
rect 18798 14662 18828 14714
rect 18852 14662 18862 14714
rect 18862 14662 18908 14714
rect 18612 14660 18668 14662
rect 18692 14660 18748 14662
rect 18772 14660 18828 14662
rect 18852 14660 18908 14662
rect 19062 13640 19118 13696
rect 18612 13626 18668 13628
rect 18692 13626 18748 13628
rect 18772 13626 18828 13628
rect 18852 13626 18908 13628
rect 18612 13574 18658 13626
rect 18658 13574 18668 13626
rect 18692 13574 18722 13626
rect 18722 13574 18734 13626
rect 18734 13574 18748 13626
rect 18772 13574 18786 13626
rect 18786 13574 18798 13626
rect 18798 13574 18828 13626
rect 18852 13574 18862 13626
rect 18862 13574 18908 13626
rect 18612 13572 18668 13574
rect 18692 13572 18748 13574
rect 18772 13572 18828 13574
rect 18852 13572 18908 13574
rect 18612 12538 18668 12540
rect 18692 12538 18748 12540
rect 18772 12538 18828 12540
rect 18852 12538 18908 12540
rect 18612 12486 18658 12538
rect 18658 12486 18668 12538
rect 18692 12486 18722 12538
rect 18722 12486 18734 12538
rect 18734 12486 18748 12538
rect 18772 12486 18786 12538
rect 18786 12486 18798 12538
rect 18798 12486 18828 12538
rect 18852 12486 18862 12538
rect 18862 12486 18908 12538
rect 18612 12484 18668 12486
rect 18692 12484 18748 12486
rect 18772 12484 18828 12486
rect 18852 12484 18908 12486
rect 18612 11450 18668 11452
rect 18692 11450 18748 11452
rect 18772 11450 18828 11452
rect 18852 11450 18908 11452
rect 18612 11398 18658 11450
rect 18658 11398 18668 11450
rect 18692 11398 18722 11450
rect 18722 11398 18734 11450
rect 18734 11398 18748 11450
rect 18772 11398 18786 11450
rect 18786 11398 18798 11450
rect 18798 11398 18828 11450
rect 18852 11398 18862 11450
rect 18862 11398 18908 11450
rect 18612 11396 18668 11398
rect 18692 11396 18748 11398
rect 18772 11396 18828 11398
rect 18852 11396 18908 11398
rect 18418 11212 18474 11248
rect 18418 11192 18420 11212
rect 18420 11192 18472 11212
rect 18472 11192 18474 11212
rect 18612 10362 18668 10364
rect 18692 10362 18748 10364
rect 18772 10362 18828 10364
rect 18852 10362 18908 10364
rect 18612 10310 18658 10362
rect 18658 10310 18668 10362
rect 18692 10310 18722 10362
rect 18722 10310 18734 10362
rect 18734 10310 18748 10362
rect 18772 10310 18786 10362
rect 18786 10310 18798 10362
rect 18798 10310 18828 10362
rect 18852 10310 18862 10362
rect 18862 10310 18908 10362
rect 18612 10308 18668 10310
rect 18692 10308 18748 10310
rect 18772 10308 18828 10310
rect 18852 10308 18908 10310
rect 18612 9274 18668 9276
rect 18692 9274 18748 9276
rect 18772 9274 18828 9276
rect 18852 9274 18908 9276
rect 18612 9222 18658 9274
rect 18658 9222 18668 9274
rect 18692 9222 18722 9274
rect 18722 9222 18734 9274
rect 18734 9222 18748 9274
rect 18772 9222 18786 9274
rect 18786 9222 18798 9274
rect 18798 9222 18828 9274
rect 18852 9222 18862 9274
rect 18862 9222 18908 9274
rect 18612 9220 18668 9222
rect 18692 9220 18748 9222
rect 18772 9220 18828 9222
rect 18852 9220 18908 9222
rect 18418 8744 18474 8800
rect 18612 8186 18668 8188
rect 18692 8186 18748 8188
rect 18772 8186 18828 8188
rect 18852 8186 18908 8188
rect 18612 8134 18658 8186
rect 18658 8134 18668 8186
rect 18692 8134 18722 8186
rect 18722 8134 18734 8186
rect 18734 8134 18748 8186
rect 18772 8134 18786 8186
rect 18786 8134 18798 8186
rect 18798 8134 18828 8186
rect 18852 8134 18862 8186
rect 18862 8134 18908 8186
rect 18612 8132 18668 8134
rect 18692 8132 18748 8134
rect 18772 8132 18828 8134
rect 18852 8132 18908 8134
rect 18612 7098 18668 7100
rect 18692 7098 18748 7100
rect 18772 7098 18828 7100
rect 18852 7098 18908 7100
rect 18612 7046 18658 7098
rect 18658 7046 18668 7098
rect 18692 7046 18722 7098
rect 18722 7046 18734 7098
rect 18734 7046 18748 7098
rect 18772 7046 18786 7098
rect 18786 7046 18798 7098
rect 18798 7046 18828 7098
rect 18852 7046 18862 7098
rect 18862 7046 18908 7098
rect 18612 7044 18668 7046
rect 18692 7044 18748 7046
rect 18772 7044 18828 7046
rect 18852 7044 18908 7046
rect 18418 6296 18474 6352
rect 18612 6010 18668 6012
rect 18692 6010 18748 6012
rect 18772 6010 18828 6012
rect 18852 6010 18908 6012
rect 18612 5958 18658 6010
rect 18658 5958 18668 6010
rect 18692 5958 18722 6010
rect 18722 5958 18734 6010
rect 18734 5958 18748 6010
rect 18772 5958 18786 6010
rect 18786 5958 18798 6010
rect 18798 5958 18828 6010
rect 18852 5958 18862 6010
rect 18862 5958 18908 6010
rect 18612 5956 18668 5958
rect 18692 5956 18748 5958
rect 18772 5956 18828 5958
rect 18852 5956 18908 5958
rect 18612 4922 18668 4924
rect 18692 4922 18748 4924
rect 18772 4922 18828 4924
rect 18852 4922 18908 4924
rect 18612 4870 18658 4922
rect 18658 4870 18668 4922
rect 18692 4870 18722 4922
rect 18722 4870 18734 4922
rect 18734 4870 18748 4922
rect 18772 4870 18786 4922
rect 18786 4870 18798 4922
rect 18798 4870 18828 4922
rect 18852 4870 18862 4922
rect 18862 4870 18908 4922
rect 18612 4868 18668 4870
rect 18692 4868 18748 4870
rect 18772 4868 18828 4870
rect 18852 4868 18908 4870
rect 19062 3848 19118 3904
rect 18612 3834 18668 3836
rect 18692 3834 18748 3836
rect 18772 3834 18828 3836
rect 18852 3834 18908 3836
rect 18612 3782 18658 3834
rect 18658 3782 18668 3834
rect 18692 3782 18722 3834
rect 18722 3782 18734 3834
rect 18734 3782 18748 3834
rect 18772 3782 18786 3834
rect 18786 3782 18798 3834
rect 18798 3782 18828 3834
rect 18852 3782 18862 3834
rect 18862 3782 18908 3834
rect 18612 3780 18668 3782
rect 18692 3780 18748 3782
rect 18772 3780 18828 3782
rect 18852 3780 18908 3782
rect 18612 2746 18668 2748
rect 18692 2746 18748 2748
rect 18772 2746 18828 2748
rect 18852 2746 18908 2748
rect 18612 2694 18658 2746
rect 18658 2694 18668 2746
rect 18692 2694 18722 2746
rect 18722 2694 18734 2746
rect 18734 2694 18748 2746
rect 18772 2694 18786 2746
rect 18786 2694 18798 2746
rect 18798 2694 18828 2746
rect 18852 2694 18862 2746
rect 18862 2694 18908 2746
rect 18612 2692 18668 2694
rect 18692 2692 18748 2694
rect 18772 2692 18828 2694
rect 18852 2692 18908 2694
rect 17062 1114 17118 1116
rect 17142 1114 17198 1116
rect 17222 1114 17278 1116
rect 17302 1114 17358 1116
rect 17062 1062 17108 1114
rect 17108 1062 17118 1114
rect 17142 1062 17172 1114
rect 17172 1062 17184 1114
rect 17184 1062 17198 1114
rect 17222 1062 17236 1114
rect 17236 1062 17248 1114
rect 17248 1062 17278 1114
rect 17302 1062 17312 1114
rect 17312 1062 17358 1114
rect 17062 1060 17118 1062
rect 17142 1060 17198 1062
rect 17222 1060 17278 1062
rect 17302 1060 17358 1062
rect 18612 1658 18668 1660
rect 18692 1658 18748 1660
rect 18772 1658 18828 1660
rect 18852 1658 18908 1660
rect 18612 1606 18658 1658
rect 18658 1606 18668 1658
rect 18692 1606 18722 1658
rect 18722 1606 18734 1658
rect 18734 1606 18748 1658
rect 18772 1606 18786 1658
rect 18786 1606 18798 1658
rect 18798 1606 18828 1658
rect 18852 1606 18862 1658
rect 18862 1606 18908 1658
rect 18612 1604 18668 1606
rect 18692 1604 18748 1606
rect 18772 1604 18828 1606
rect 18852 1604 18908 1606
rect 18418 1400 18474 1456
rect 3112 570 3168 572
rect 3192 570 3248 572
rect 3272 570 3328 572
rect 3352 570 3408 572
rect 3112 518 3158 570
rect 3158 518 3168 570
rect 3192 518 3222 570
rect 3222 518 3234 570
rect 3234 518 3248 570
rect 3272 518 3286 570
rect 3286 518 3298 570
rect 3298 518 3328 570
rect 3352 518 3362 570
rect 3362 518 3408 570
rect 3112 516 3168 518
rect 3192 516 3248 518
rect 3272 516 3328 518
rect 3352 516 3408 518
rect 6212 570 6268 572
rect 6292 570 6348 572
rect 6372 570 6428 572
rect 6452 570 6508 572
rect 6212 518 6258 570
rect 6258 518 6268 570
rect 6292 518 6322 570
rect 6322 518 6334 570
rect 6334 518 6348 570
rect 6372 518 6386 570
rect 6386 518 6398 570
rect 6398 518 6428 570
rect 6452 518 6462 570
rect 6462 518 6508 570
rect 6212 516 6268 518
rect 6292 516 6348 518
rect 6372 516 6428 518
rect 6452 516 6508 518
rect 9312 570 9368 572
rect 9392 570 9448 572
rect 9472 570 9528 572
rect 9552 570 9608 572
rect 9312 518 9358 570
rect 9358 518 9368 570
rect 9392 518 9422 570
rect 9422 518 9434 570
rect 9434 518 9448 570
rect 9472 518 9486 570
rect 9486 518 9498 570
rect 9498 518 9528 570
rect 9552 518 9562 570
rect 9562 518 9608 570
rect 9312 516 9368 518
rect 9392 516 9448 518
rect 9472 516 9528 518
rect 9552 516 9608 518
rect 12412 570 12468 572
rect 12492 570 12548 572
rect 12572 570 12628 572
rect 12652 570 12708 572
rect 12412 518 12458 570
rect 12458 518 12468 570
rect 12492 518 12522 570
rect 12522 518 12534 570
rect 12534 518 12548 570
rect 12572 518 12586 570
rect 12586 518 12598 570
rect 12598 518 12628 570
rect 12652 518 12662 570
rect 12662 518 12708 570
rect 12412 516 12468 518
rect 12492 516 12548 518
rect 12572 516 12628 518
rect 12652 516 12708 518
rect 15512 570 15568 572
rect 15592 570 15648 572
rect 15672 570 15728 572
rect 15752 570 15808 572
rect 15512 518 15558 570
rect 15558 518 15568 570
rect 15592 518 15622 570
rect 15622 518 15634 570
rect 15634 518 15648 570
rect 15672 518 15686 570
rect 15686 518 15698 570
rect 15698 518 15728 570
rect 15752 518 15762 570
rect 15762 518 15808 570
rect 15512 516 15568 518
rect 15592 516 15648 518
rect 15672 516 15728 518
rect 15752 516 15808 518
rect 18612 570 18668 572
rect 18692 570 18748 572
rect 18772 570 18828 572
rect 18852 570 18908 572
rect 18612 518 18658 570
rect 18658 518 18668 570
rect 18692 518 18722 570
rect 18722 518 18734 570
rect 18734 518 18748 570
rect 18772 518 18786 570
rect 18786 518 18798 570
rect 18798 518 18828 570
rect 18852 518 18862 570
rect 18862 518 18908 570
rect 18612 516 18668 518
rect 18692 516 18748 518
rect 18772 516 18828 518
rect 18852 516 18908 518
<< metal3 >>
rect 18413 18594 18479 18597
rect 19200 18594 20000 18624
rect 18413 18592 20000 18594
rect 18413 18536 18418 18592
rect 18474 18536 20000 18592
rect 18413 18534 20000 18536
rect 18413 18531 18479 18534
rect 1552 18528 1868 18529
rect 1552 18464 1558 18528
rect 1622 18464 1638 18528
rect 1702 18464 1718 18528
rect 1782 18464 1798 18528
rect 1862 18464 1868 18528
rect 1552 18463 1868 18464
rect 4652 18528 4968 18529
rect 4652 18464 4658 18528
rect 4722 18464 4738 18528
rect 4802 18464 4818 18528
rect 4882 18464 4898 18528
rect 4962 18464 4968 18528
rect 4652 18463 4968 18464
rect 7752 18528 8068 18529
rect 7752 18464 7758 18528
rect 7822 18464 7838 18528
rect 7902 18464 7918 18528
rect 7982 18464 7998 18528
rect 8062 18464 8068 18528
rect 7752 18463 8068 18464
rect 10852 18528 11168 18529
rect 10852 18464 10858 18528
rect 10922 18464 10938 18528
rect 11002 18464 11018 18528
rect 11082 18464 11098 18528
rect 11162 18464 11168 18528
rect 10852 18463 11168 18464
rect 13952 18528 14268 18529
rect 13952 18464 13958 18528
rect 14022 18464 14038 18528
rect 14102 18464 14118 18528
rect 14182 18464 14198 18528
rect 14262 18464 14268 18528
rect 13952 18463 14268 18464
rect 17052 18528 17368 18529
rect 17052 18464 17058 18528
rect 17122 18464 17138 18528
rect 17202 18464 17218 18528
rect 17282 18464 17298 18528
rect 17362 18464 17368 18528
rect 19200 18504 20000 18534
rect 17052 18463 17368 18464
rect 3102 17984 3418 17985
rect 3102 17920 3108 17984
rect 3172 17920 3188 17984
rect 3252 17920 3268 17984
rect 3332 17920 3348 17984
rect 3412 17920 3418 17984
rect 3102 17919 3418 17920
rect 6202 17984 6518 17985
rect 6202 17920 6208 17984
rect 6272 17920 6288 17984
rect 6352 17920 6368 17984
rect 6432 17920 6448 17984
rect 6512 17920 6518 17984
rect 6202 17919 6518 17920
rect 9302 17984 9618 17985
rect 9302 17920 9308 17984
rect 9372 17920 9388 17984
rect 9452 17920 9468 17984
rect 9532 17920 9548 17984
rect 9612 17920 9618 17984
rect 9302 17919 9618 17920
rect 12402 17984 12718 17985
rect 12402 17920 12408 17984
rect 12472 17920 12488 17984
rect 12552 17920 12568 17984
rect 12632 17920 12648 17984
rect 12712 17920 12718 17984
rect 12402 17919 12718 17920
rect 15502 17984 15818 17985
rect 15502 17920 15508 17984
rect 15572 17920 15588 17984
rect 15652 17920 15668 17984
rect 15732 17920 15748 17984
rect 15812 17920 15818 17984
rect 15502 17919 15818 17920
rect 18602 17984 18918 17985
rect 18602 17920 18608 17984
rect 18672 17920 18688 17984
rect 18752 17920 18768 17984
rect 18832 17920 18848 17984
rect 18912 17920 18918 17984
rect 18602 17919 18918 17920
rect 1552 17440 1868 17441
rect 1552 17376 1558 17440
rect 1622 17376 1638 17440
rect 1702 17376 1718 17440
rect 1782 17376 1798 17440
rect 1862 17376 1868 17440
rect 1552 17375 1868 17376
rect 4652 17440 4968 17441
rect 4652 17376 4658 17440
rect 4722 17376 4738 17440
rect 4802 17376 4818 17440
rect 4882 17376 4898 17440
rect 4962 17376 4968 17440
rect 4652 17375 4968 17376
rect 7752 17440 8068 17441
rect 7752 17376 7758 17440
rect 7822 17376 7838 17440
rect 7902 17376 7918 17440
rect 7982 17376 7998 17440
rect 8062 17376 8068 17440
rect 7752 17375 8068 17376
rect 10852 17440 11168 17441
rect 10852 17376 10858 17440
rect 10922 17376 10938 17440
rect 11002 17376 11018 17440
rect 11082 17376 11098 17440
rect 11162 17376 11168 17440
rect 10852 17375 11168 17376
rect 13952 17440 14268 17441
rect 13952 17376 13958 17440
rect 14022 17376 14038 17440
rect 14102 17376 14118 17440
rect 14182 17376 14198 17440
rect 14262 17376 14268 17440
rect 13952 17375 14268 17376
rect 17052 17440 17368 17441
rect 17052 17376 17058 17440
rect 17122 17376 17138 17440
rect 17202 17376 17218 17440
rect 17282 17376 17298 17440
rect 17362 17376 17368 17440
rect 17052 17375 17368 17376
rect 3102 16896 3418 16897
rect 3102 16832 3108 16896
rect 3172 16832 3188 16896
rect 3252 16832 3268 16896
rect 3332 16832 3348 16896
rect 3412 16832 3418 16896
rect 3102 16831 3418 16832
rect 6202 16896 6518 16897
rect 6202 16832 6208 16896
rect 6272 16832 6288 16896
rect 6352 16832 6368 16896
rect 6432 16832 6448 16896
rect 6512 16832 6518 16896
rect 6202 16831 6518 16832
rect 9302 16896 9618 16897
rect 9302 16832 9308 16896
rect 9372 16832 9388 16896
rect 9452 16832 9468 16896
rect 9532 16832 9548 16896
rect 9612 16832 9618 16896
rect 9302 16831 9618 16832
rect 12402 16896 12718 16897
rect 12402 16832 12408 16896
rect 12472 16832 12488 16896
rect 12552 16832 12568 16896
rect 12632 16832 12648 16896
rect 12712 16832 12718 16896
rect 12402 16831 12718 16832
rect 15502 16896 15818 16897
rect 15502 16832 15508 16896
rect 15572 16832 15588 16896
rect 15652 16832 15668 16896
rect 15732 16832 15748 16896
rect 15812 16832 15818 16896
rect 15502 16831 15818 16832
rect 18602 16896 18918 16897
rect 18602 16832 18608 16896
rect 18672 16832 18688 16896
rect 18752 16832 18768 16896
rect 18832 16832 18848 16896
rect 18912 16832 18918 16896
rect 18602 16831 18918 16832
rect 1552 16352 1868 16353
rect 1552 16288 1558 16352
rect 1622 16288 1638 16352
rect 1702 16288 1718 16352
rect 1782 16288 1798 16352
rect 1862 16288 1868 16352
rect 1552 16287 1868 16288
rect 4652 16352 4968 16353
rect 4652 16288 4658 16352
rect 4722 16288 4738 16352
rect 4802 16288 4818 16352
rect 4882 16288 4898 16352
rect 4962 16288 4968 16352
rect 4652 16287 4968 16288
rect 7752 16352 8068 16353
rect 7752 16288 7758 16352
rect 7822 16288 7838 16352
rect 7902 16288 7918 16352
rect 7982 16288 7998 16352
rect 8062 16288 8068 16352
rect 7752 16287 8068 16288
rect 10852 16352 11168 16353
rect 10852 16288 10858 16352
rect 10922 16288 10938 16352
rect 11002 16288 11018 16352
rect 11082 16288 11098 16352
rect 11162 16288 11168 16352
rect 10852 16287 11168 16288
rect 13952 16352 14268 16353
rect 13952 16288 13958 16352
rect 14022 16288 14038 16352
rect 14102 16288 14118 16352
rect 14182 16288 14198 16352
rect 14262 16288 14268 16352
rect 13952 16287 14268 16288
rect 17052 16352 17368 16353
rect 17052 16288 17058 16352
rect 17122 16288 17138 16352
rect 17202 16288 17218 16352
rect 17282 16288 17298 16352
rect 17362 16288 17368 16352
rect 17052 16287 17368 16288
rect 18413 16146 18479 16149
rect 19200 16146 20000 16176
rect 18413 16144 20000 16146
rect 18413 16088 18418 16144
rect 18474 16088 20000 16144
rect 18413 16086 20000 16088
rect 18413 16083 18479 16086
rect 19200 16056 20000 16086
rect 3102 15808 3418 15809
rect 3102 15744 3108 15808
rect 3172 15744 3188 15808
rect 3252 15744 3268 15808
rect 3332 15744 3348 15808
rect 3412 15744 3418 15808
rect 3102 15743 3418 15744
rect 6202 15808 6518 15809
rect 6202 15744 6208 15808
rect 6272 15744 6288 15808
rect 6352 15744 6368 15808
rect 6432 15744 6448 15808
rect 6512 15744 6518 15808
rect 6202 15743 6518 15744
rect 9302 15808 9618 15809
rect 9302 15744 9308 15808
rect 9372 15744 9388 15808
rect 9452 15744 9468 15808
rect 9532 15744 9548 15808
rect 9612 15744 9618 15808
rect 9302 15743 9618 15744
rect 12402 15808 12718 15809
rect 12402 15744 12408 15808
rect 12472 15744 12488 15808
rect 12552 15744 12568 15808
rect 12632 15744 12648 15808
rect 12712 15744 12718 15808
rect 12402 15743 12718 15744
rect 15502 15808 15818 15809
rect 15502 15744 15508 15808
rect 15572 15744 15588 15808
rect 15652 15744 15668 15808
rect 15732 15744 15748 15808
rect 15812 15744 15818 15808
rect 15502 15743 15818 15744
rect 18602 15808 18918 15809
rect 18602 15744 18608 15808
rect 18672 15744 18688 15808
rect 18752 15744 18768 15808
rect 18832 15744 18848 15808
rect 18912 15744 18918 15808
rect 18602 15743 18918 15744
rect 1552 15264 1868 15265
rect 1552 15200 1558 15264
rect 1622 15200 1638 15264
rect 1702 15200 1718 15264
rect 1782 15200 1798 15264
rect 1862 15200 1868 15264
rect 1552 15199 1868 15200
rect 4652 15264 4968 15265
rect 4652 15200 4658 15264
rect 4722 15200 4738 15264
rect 4802 15200 4818 15264
rect 4882 15200 4898 15264
rect 4962 15200 4968 15264
rect 4652 15199 4968 15200
rect 7752 15264 8068 15265
rect 7752 15200 7758 15264
rect 7822 15200 7838 15264
rect 7902 15200 7918 15264
rect 7982 15200 7998 15264
rect 8062 15200 8068 15264
rect 7752 15199 8068 15200
rect 10852 15264 11168 15265
rect 10852 15200 10858 15264
rect 10922 15200 10938 15264
rect 11002 15200 11018 15264
rect 11082 15200 11098 15264
rect 11162 15200 11168 15264
rect 10852 15199 11168 15200
rect 13952 15264 14268 15265
rect 13952 15200 13958 15264
rect 14022 15200 14038 15264
rect 14102 15200 14118 15264
rect 14182 15200 14198 15264
rect 14262 15200 14268 15264
rect 13952 15199 14268 15200
rect 17052 15264 17368 15265
rect 17052 15200 17058 15264
rect 17122 15200 17138 15264
rect 17202 15200 17218 15264
rect 17282 15200 17298 15264
rect 17362 15200 17368 15264
rect 17052 15199 17368 15200
rect 3102 14720 3418 14721
rect 3102 14656 3108 14720
rect 3172 14656 3188 14720
rect 3252 14656 3268 14720
rect 3332 14656 3348 14720
rect 3412 14656 3418 14720
rect 3102 14655 3418 14656
rect 6202 14720 6518 14721
rect 6202 14656 6208 14720
rect 6272 14656 6288 14720
rect 6352 14656 6368 14720
rect 6432 14656 6448 14720
rect 6512 14656 6518 14720
rect 6202 14655 6518 14656
rect 9302 14720 9618 14721
rect 9302 14656 9308 14720
rect 9372 14656 9388 14720
rect 9452 14656 9468 14720
rect 9532 14656 9548 14720
rect 9612 14656 9618 14720
rect 9302 14655 9618 14656
rect 12402 14720 12718 14721
rect 12402 14656 12408 14720
rect 12472 14656 12488 14720
rect 12552 14656 12568 14720
rect 12632 14656 12648 14720
rect 12712 14656 12718 14720
rect 12402 14655 12718 14656
rect 15502 14720 15818 14721
rect 15502 14656 15508 14720
rect 15572 14656 15588 14720
rect 15652 14656 15668 14720
rect 15732 14656 15748 14720
rect 15812 14656 15818 14720
rect 15502 14655 15818 14656
rect 18602 14720 18918 14721
rect 18602 14656 18608 14720
rect 18672 14656 18688 14720
rect 18752 14656 18768 14720
rect 18832 14656 18848 14720
rect 18912 14656 18918 14720
rect 18602 14655 18918 14656
rect 1552 14176 1868 14177
rect 1552 14112 1558 14176
rect 1622 14112 1638 14176
rect 1702 14112 1718 14176
rect 1782 14112 1798 14176
rect 1862 14112 1868 14176
rect 1552 14111 1868 14112
rect 4652 14176 4968 14177
rect 4652 14112 4658 14176
rect 4722 14112 4738 14176
rect 4802 14112 4818 14176
rect 4882 14112 4898 14176
rect 4962 14112 4968 14176
rect 4652 14111 4968 14112
rect 7752 14176 8068 14177
rect 7752 14112 7758 14176
rect 7822 14112 7838 14176
rect 7902 14112 7918 14176
rect 7982 14112 7998 14176
rect 8062 14112 8068 14176
rect 7752 14111 8068 14112
rect 10852 14176 11168 14177
rect 10852 14112 10858 14176
rect 10922 14112 10938 14176
rect 11002 14112 11018 14176
rect 11082 14112 11098 14176
rect 11162 14112 11168 14176
rect 10852 14111 11168 14112
rect 13952 14176 14268 14177
rect 13952 14112 13958 14176
rect 14022 14112 14038 14176
rect 14102 14112 14118 14176
rect 14182 14112 14198 14176
rect 14262 14112 14268 14176
rect 13952 14111 14268 14112
rect 17052 14176 17368 14177
rect 17052 14112 17058 14176
rect 17122 14112 17138 14176
rect 17202 14112 17218 14176
rect 17282 14112 17298 14176
rect 17362 14112 17368 14176
rect 17052 14111 17368 14112
rect 19057 13698 19123 13701
rect 19200 13698 20000 13728
rect 19057 13696 20000 13698
rect 19057 13640 19062 13696
rect 19118 13640 20000 13696
rect 19057 13638 20000 13640
rect 19057 13635 19123 13638
rect 3102 13632 3418 13633
rect 3102 13568 3108 13632
rect 3172 13568 3188 13632
rect 3252 13568 3268 13632
rect 3332 13568 3348 13632
rect 3412 13568 3418 13632
rect 3102 13567 3418 13568
rect 6202 13632 6518 13633
rect 6202 13568 6208 13632
rect 6272 13568 6288 13632
rect 6352 13568 6368 13632
rect 6432 13568 6448 13632
rect 6512 13568 6518 13632
rect 6202 13567 6518 13568
rect 9302 13632 9618 13633
rect 9302 13568 9308 13632
rect 9372 13568 9388 13632
rect 9452 13568 9468 13632
rect 9532 13568 9548 13632
rect 9612 13568 9618 13632
rect 9302 13567 9618 13568
rect 12402 13632 12718 13633
rect 12402 13568 12408 13632
rect 12472 13568 12488 13632
rect 12552 13568 12568 13632
rect 12632 13568 12648 13632
rect 12712 13568 12718 13632
rect 12402 13567 12718 13568
rect 15502 13632 15818 13633
rect 15502 13568 15508 13632
rect 15572 13568 15588 13632
rect 15652 13568 15668 13632
rect 15732 13568 15748 13632
rect 15812 13568 15818 13632
rect 15502 13567 15818 13568
rect 18602 13632 18918 13633
rect 18602 13568 18608 13632
rect 18672 13568 18688 13632
rect 18752 13568 18768 13632
rect 18832 13568 18848 13632
rect 18912 13568 18918 13632
rect 19200 13608 20000 13638
rect 18602 13567 18918 13568
rect 1552 13088 1868 13089
rect 1552 13024 1558 13088
rect 1622 13024 1638 13088
rect 1702 13024 1718 13088
rect 1782 13024 1798 13088
rect 1862 13024 1868 13088
rect 1552 13023 1868 13024
rect 4652 13088 4968 13089
rect 4652 13024 4658 13088
rect 4722 13024 4738 13088
rect 4802 13024 4818 13088
rect 4882 13024 4898 13088
rect 4962 13024 4968 13088
rect 4652 13023 4968 13024
rect 7752 13088 8068 13089
rect 7752 13024 7758 13088
rect 7822 13024 7838 13088
rect 7902 13024 7918 13088
rect 7982 13024 7998 13088
rect 8062 13024 8068 13088
rect 7752 13023 8068 13024
rect 10852 13088 11168 13089
rect 10852 13024 10858 13088
rect 10922 13024 10938 13088
rect 11002 13024 11018 13088
rect 11082 13024 11098 13088
rect 11162 13024 11168 13088
rect 10852 13023 11168 13024
rect 13952 13088 14268 13089
rect 13952 13024 13958 13088
rect 14022 13024 14038 13088
rect 14102 13024 14118 13088
rect 14182 13024 14198 13088
rect 14262 13024 14268 13088
rect 13952 13023 14268 13024
rect 17052 13088 17368 13089
rect 17052 13024 17058 13088
rect 17122 13024 17138 13088
rect 17202 13024 17218 13088
rect 17282 13024 17298 13088
rect 17362 13024 17368 13088
rect 17052 13023 17368 13024
rect 3102 12544 3418 12545
rect 3102 12480 3108 12544
rect 3172 12480 3188 12544
rect 3252 12480 3268 12544
rect 3332 12480 3348 12544
rect 3412 12480 3418 12544
rect 3102 12479 3418 12480
rect 6202 12544 6518 12545
rect 6202 12480 6208 12544
rect 6272 12480 6288 12544
rect 6352 12480 6368 12544
rect 6432 12480 6448 12544
rect 6512 12480 6518 12544
rect 6202 12479 6518 12480
rect 9302 12544 9618 12545
rect 9302 12480 9308 12544
rect 9372 12480 9388 12544
rect 9452 12480 9468 12544
rect 9532 12480 9548 12544
rect 9612 12480 9618 12544
rect 9302 12479 9618 12480
rect 12402 12544 12718 12545
rect 12402 12480 12408 12544
rect 12472 12480 12488 12544
rect 12552 12480 12568 12544
rect 12632 12480 12648 12544
rect 12712 12480 12718 12544
rect 12402 12479 12718 12480
rect 15502 12544 15818 12545
rect 15502 12480 15508 12544
rect 15572 12480 15588 12544
rect 15652 12480 15668 12544
rect 15732 12480 15748 12544
rect 15812 12480 15818 12544
rect 15502 12479 15818 12480
rect 18602 12544 18918 12545
rect 18602 12480 18608 12544
rect 18672 12480 18688 12544
rect 18752 12480 18768 12544
rect 18832 12480 18848 12544
rect 18912 12480 18918 12544
rect 18602 12479 18918 12480
rect 1552 12000 1868 12001
rect 1552 11936 1558 12000
rect 1622 11936 1638 12000
rect 1702 11936 1718 12000
rect 1782 11936 1798 12000
rect 1862 11936 1868 12000
rect 1552 11935 1868 11936
rect 4652 12000 4968 12001
rect 4652 11936 4658 12000
rect 4722 11936 4738 12000
rect 4802 11936 4818 12000
rect 4882 11936 4898 12000
rect 4962 11936 4968 12000
rect 4652 11935 4968 11936
rect 7752 12000 8068 12001
rect 7752 11936 7758 12000
rect 7822 11936 7838 12000
rect 7902 11936 7918 12000
rect 7982 11936 7998 12000
rect 8062 11936 8068 12000
rect 7752 11935 8068 11936
rect 10852 12000 11168 12001
rect 10852 11936 10858 12000
rect 10922 11936 10938 12000
rect 11002 11936 11018 12000
rect 11082 11936 11098 12000
rect 11162 11936 11168 12000
rect 10852 11935 11168 11936
rect 13952 12000 14268 12001
rect 13952 11936 13958 12000
rect 14022 11936 14038 12000
rect 14102 11936 14118 12000
rect 14182 11936 14198 12000
rect 14262 11936 14268 12000
rect 13952 11935 14268 11936
rect 17052 12000 17368 12001
rect 17052 11936 17058 12000
rect 17122 11936 17138 12000
rect 17202 11936 17218 12000
rect 17282 11936 17298 12000
rect 17362 11936 17368 12000
rect 17052 11935 17368 11936
rect 3102 11456 3418 11457
rect 3102 11392 3108 11456
rect 3172 11392 3188 11456
rect 3252 11392 3268 11456
rect 3332 11392 3348 11456
rect 3412 11392 3418 11456
rect 3102 11391 3418 11392
rect 6202 11456 6518 11457
rect 6202 11392 6208 11456
rect 6272 11392 6288 11456
rect 6352 11392 6368 11456
rect 6432 11392 6448 11456
rect 6512 11392 6518 11456
rect 6202 11391 6518 11392
rect 9302 11456 9618 11457
rect 9302 11392 9308 11456
rect 9372 11392 9388 11456
rect 9452 11392 9468 11456
rect 9532 11392 9548 11456
rect 9612 11392 9618 11456
rect 9302 11391 9618 11392
rect 12402 11456 12718 11457
rect 12402 11392 12408 11456
rect 12472 11392 12488 11456
rect 12552 11392 12568 11456
rect 12632 11392 12648 11456
rect 12712 11392 12718 11456
rect 12402 11391 12718 11392
rect 15502 11456 15818 11457
rect 15502 11392 15508 11456
rect 15572 11392 15588 11456
rect 15652 11392 15668 11456
rect 15732 11392 15748 11456
rect 15812 11392 15818 11456
rect 15502 11391 15818 11392
rect 18602 11456 18918 11457
rect 18602 11392 18608 11456
rect 18672 11392 18688 11456
rect 18752 11392 18768 11456
rect 18832 11392 18848 11456
rect 18912 11392 18918 11456
rect 18602 11391 18918 11392
rect 18413 11250 18479 11253
rect 19200 11250 20000 11280
rect 18413 11248 20000 11250
rect 18413 11192 18418 11248
rect 18474 11192 20000 11248
rect 18413 11190 20000 11192
rect 18413 11187 18479 11190
rect 19200 11160 20000 11190
rect 1552 10912 1868 10913
rect 1552 10848 1558 10912
rect 1622 10848 1638 10912
rect 1702 10848 1718 10912
rect 1782 10848 1798 10912
rect 1862 10848 1868 10912
rect 1552 10847 1868 10848
rect 4652 10912 4968 10913
rect 4652 10848 4658 10912
rect 4722 10848 4738 10912
rect 4802 10848 4818 10912
rect 4882 10848 4898 10912
rect 4962 10848 4968 10912
rect 4652 10847 4968 10848
rect 7752 10912 8068 10913
rect 7752 10848 7758 10912
rect 7822 10848 7838 10912
rect 7902 10848 7918 10912
rect 7982 10848 7998 10912
rect 8062 10848 8068 10912
rect 7752 10847 8068 10848
rect 10852 10912 11168 10913
rect 10852 10848 10858 10912
rect 10922 10848 10938 10912
rect 11002 10848 11018 10912
rect 11082 10848 11098 10912
rect 11162 10848 11168 10912
rect 10852 10847 11168 10848
rect 13952 10912 14268 10913
rect 13952 10848 13958 10912
rect 14022 10848 14038 10912
rect 14102 10848 14118 10912
rect 14182 10848 14198 10912
rect 14262 10848 14268 10912
rect 13952 10847 14268 10848
rect 17052 10912 17368 10913
rect 17052 10848 17058 10912
rect 17122 10848 17138 10912
rect 17202 10848 17218 10912
rect 17282 10848 17298 10912
rect 17362 10848 17368 10912
rect 17052 10847 17368 10848
rect 3102 10368 3418 10369
rect 3102 10304 3108 10368
rect 3172 10304 3188 10368
rect 3252 10304 3268 10368
rect 3332 10304 3348 10368
rect 3412 10304 3418 10368
rect 3102 10303 3418 10304
rect 6202 10368 6518 10369
rect 6202 10304 6208 10368
rect 6272 10304 6288 10368
rect 6352 10304 6368 10368
rect 6432 10304 6448 10368
rect 6512 10304 6518 10368
rect 6202 10303 6518 10304
rect 9302 10368 9618 10369
rect 9302 10304 9308 10368
rect 9372 10304 9388 10368
rect 9452 10304 9468 10368
rect 9532 10304 9548 10368
rect 9612 10304 9618 10368
rect 9302 10303 9618 10304
rect 12402 10368 12718 10369
rect 12402 10304 12408 10368
rect 12472 10304 12488 10368
rect 12552 10304 12568 10368
rect 12632 10304 12648 10368
rect 12712 10304 12718 10368
rect 12402 10303 12718 10304
rect 15502 10368 15818 10369
rect 15502 10304 15508 10368
rect 15572 10304 15588 10368
rect 15652 10304 15668 10368
rect 15732 10304 15748 10368
rect 15812 10304 15818 10368
rect 15502 10303 15818 10304
rect 18602 10368 18918 10369
rect 18602 10304 18608 10368
rect 18672 10304 18688 10368
rect 18752 10304 18768 10368
rect 18832 10304 18848 10368
rect 18912 10304 18918 10368
rect 18602 10303 18918 10304
rect 1552 9824 1868 9825
rect 1552 9760 1558 9824
rect 1622 9760 1638 9824
rect 1702 9760 1718 9824
rect 1782 9760 1798 9824
rect 1862 9760 1868 9824
rect 1552 9759 1868 9760
rect 4652 9824 4968 9825
rect 4652 9760 4658 9824
rect 4722 9760 4738 9824
rect 4802 9760 4818 9824
rect 4882 9760 4898 9824
rect 4962 9760 4968 9824
rect 4652 9759 4968 9760
rect 7752 9824 8068 9825
rect 7752 9760 7758 9824
rect 7822 9760 7838 9824
rect 7902 9760 7918 9824
rect 7982 9760 7998 9824
rect 8062 9760 8068 9824
rect 7752 9759 8068 9760
rect 10852 9824 11168 9825
rect 10852 9760 10858 9824
rect 10922 9760 10938 9824
rect 11002 9760 11018 9824
rect 11082 9760 11098 9824
rect 11162 9760 11168 9824
rect 10852 9759 11168 9760
rect 13952 9824 14268 9825
rect 13952 9760 13958 9824
rect 14022 9760 14038 9824
rect 14102 9760 14118 9824
rect 14182 9760 14198 9824
rect 14262 9760 14268 9824
rect 13952 9759 14268 9760
rect 17052 9824 17368 9825
rect 17052 9760 17058 9824
rect 17122 9760 17138 9824
rect 17202 9760 17218 9824
rect 17282 9760 17298 9824
rect 17362 9760 17368 9824
rect 17052 9759 17368 9760
rect 3102 9280 3418 9281
rect 3102 9216 3108 9280
rect 3172 9216 3188 9280
rect 3252 9216 3268 9280
rect 3332 9216 3348 9280
rect 3412 9216 3418 9280
rect 3102 9215 3418 9216
rect 6202 9280 6518 9281
rect 6202 9216 6208 9280
rect 6272 9216 6288 9280
rect 6352 9216 6368 9280
rect 6432 9216 6448 9280
rect 6512 9216 6518 9280
rect 6202 9215 6518 9216
rect 9302 9280 9618 9281
rect 9302 9216 9308 9280
rect 9372 9216 9388 9280
rect 9452 9216 9468 9280
rect 9532 9216 9548 9280
rect 9612 9216 9618 9280
rect 9302 9215 9618 9216
rect 12402 9280 12718 9281
rect 12402 9216 12408 9280
rect 12472 9216 12488 9280
rect 12552 9216 12568 9280
rect 12632 9216 12648 9280
rect 12712 9216 12718 9280
rect 12402 9215 12718 9216
rect 15502 9280 15818 9281
rect 15502 9216 15508 9280
rect 15572 9216 15588 9280
rect 15652 9216 15668 9280
rect 15732 9216 15748 9280
rect 15812 9216 15818 9280
rect 15502 9215 15818 9216
rect 18602 9280 18918 9281
rect 18602 9216 18608 9280
rect 18672 9216 18688 9280
rect 18752 9216 18768 9280
rect 18832 9216 18848 9280
rect 18912 9216 18918 9280
rect 18602 9215 18918 9216
rect 18413 8802 18479 8805
rect 19200 8802 20000 8832
rect 18413 8800 20000 8802
rect 18413 8744 18418 8800
rect 18474 8744 20000 8800
rect 18413 8742 20000 8744
rect 18413 8739 18479 8742
rect 1552 8736 1868 8737
rect 1552 8672 1558 8736
rect 1622 8672 1638 8736
rect 1702 8672 1718 8736
rect 1782 8672 1798 8736
rect 1862 8672 1868 8736
rect 1552 8671 1868 8672
rect 4652 8736 4968 8737
rect 4652 8672 4658 8736
rect 4722 8672 4738 8736
rect 4802 8672 4818 8736
rect 4882 8672 4898 8736
rect 4962 8672 4968 8736
rect 4652 8671 4968 8672
rect 7752 8736 8068 8737
rect 7752 8672 7758 8736
rect 7822 8672 7838 8736
rect 7902 8672 7918 8736
rect 7982 8672 7998 8736
rect 8062 8672 8068 8736
rect 7752 8671 8068 8672
rect 10852 8736 11168 8737
rect 10852 8672 10858 8736
rect 10922 8672 10938 8736
rect 11002 8672 11018 8736
rect 11082 8672 11098 8736
rect 11162 8672 11168 8736
rect 10852 8671 11168 8672
rect 13952 8736 14268 8737
rect 13952 8672 13958 8736
rect 14022 8672 14038 8736
rect 14102 8672 14118 8736
rect 14182 8672 14198 8736
rect 14262 8672 14268 8736
rect 13952 8671 14268 8672
rect 17052 8736 17368 8737
rect 17052 8672 17058 8736
rect 17122 8672 17138 8736
rect 17202 8672 17218 8736
rect 17282 8672 17298 8736
rect 17362 8672 17368 8736
rect 19200 8712 20000 8742
rect 17052 8671 17368 8672
rect 3102 8192 3418 8193
rect 3102 8128 3108 8192
rect 3172 8128 3188 8192
rect 3252 8128 3268 8192
rect 3332 8128 3348 8192
rect 3412 8128 3418 8192
rect 3102 8127 3418 8128
rect 6202 8192 6518 8193
rect 6202 8128 6208 8192
rect 6272 8128 6288 8192
rect 6352 8128 6368 8192
rect 6432 8128 6448 8192
rect 6512 8128 6518 8192
rect 6202 8127 6518 8128
rect 9302 8192 9618 8193
rect 9302 8128 9308 8192
rect 9372 8128 9388 8192
rect 9452 8128 9468 8192
rect 9532 8128 9548 8192
rect 9612 8128 9618 8192
rect 9302 8127 9618 8128
rect 12402 8192 12718 8193
rect 12402 8128 12408 8192
rect 12472 8128 12488 8192
rect 12552 8128 12568 8192
rect 12632 8128 12648 8192
rect 12712 8128 12718 8192
rect 12402 8127 12718 8128
rect 15502 8192 15818 8193
rect 15502 8128 15508 8192
rect 15572 8128 15588 8192
rect 15652 8128 15668 8192
rect 15732 8128 15748 8192
rect 15812 8128 15818 8192
rect 15502 8127 15818 8128
rect 18602 8192 18918 8193
rect 18602 8128 18608 8192
rect 18672 8128 18688 8192
rect 18752 8128 18768 8192
rect 18832 8128 18848 8192
rect 18912 8128 18918 8192
rect 18602 8127 18918 8128
rect 1552 7648 1868 7649
rect 1552 7584 1558 7648
rect 1622 7584 1638 7648
rect 1702 7584 1718 7648
rect 1782 7584 1798 7648
rect 1862 7584 1868 7648
rect 1552 7583 1868 7584
rect 4652 7648 4968 7649
rect 4652 7584 4658 7648
rect 4722 7584 4738 7648
rect 4802 7584 4818 7648
rect 4882 7584 4898 7648
rect 4962 7584 4968 7648
rect 4652 7583 4968 7584
rect 7752 7648 8068 7649
rect 7752 7584 7758 7648
rect 7822 7584 7838 7648
rect 7902 7584 7918 7648
rect 7982 7584 7998 7648
rect 8062 7584 8068 7648
rect 7752 7583 8068 7584
rect 10852 7648 11168 7649
rect 10852 7584 10858 7648
rect 10922 7584 10938 7648
rect 11002 7584 11018 7648
rect 11082 7584 11098 7648
rect 11162 7584 11168 7648
rect 10852 7583 11168 7584
rect 13952 7648 14268 7649
rect 13952 7584 13958 7648
rect 14022 7584 14038 7648
rect 14102 7584 14118 7648
rect 14182 7584 14198 7648
rect 14262 7584 14268 7648
rect 13952 7583 14268 7584
rect 17052 7648 17368 7649
rect 17052 7584 17058 7648
rect 17122 7584 17138 7648
rect 17202 7584 17218 7648
rect 17282 7584 17298 7648
rect 17362 7584 17368 7648
rect 17052 7583 17368 7584
rect 3102 7104 3418 7105
rect 3102 7040 3108 7104
rect 3172 7040 3188 7104
rect 3252 7040 3268 7104
rect 3332 7040 3348 7104
rect 3412 7040 3418 7104
rect 3102 7039 3418 7040
rect 6202 7104 6518 7105
rect 6202 7040 6208 7104
rect 6272 7040 6288 7104
rect 6352 7040 6368 7104
rect 6432 7040 6448 7104
rect 6512 7040 6518 7104
rect 6202 7039 6518 7040
rect 9302 7104 9618 7105
rect 9302 7040 9308 7104
rect 9372 7040 9388 7104
rect 9452 7040 9468 7104
rect 9532 7040 9548 7104
rect 9612 7040 9618 7104
rect 9302 7039 9618 7040
rect 12402 7104 12718 7105
rect 12402 7040 12408 7104
rect 12472 7040 12488 7104
rect 12552 7040 12568 7104
rect 12632 7040 12648 7104
rect 12712 7040 12718 7104
rect 12402 7039 12718 7040
rect 15502 7104 15818 7105
rect 15502 7040 15508 7104
rect 15572 7040 15588 7104
rect 15652 7040 15668 7104
rect 15732 7040 15748 7104
rect 15812 7040 15818 7104
rect 15502 7039 15818 7040
rect 18602 7104 18918 7105
rect 18602 7040 18608 7104
rect 18672 7040 18688 7104
rect 18752 7040 18768 7104
rect 18832 7040 18848 7104
rect 18912 7040 18918 7104
rect 18602 7039 18918 7040
rect 1552 6560 1868 6561
rect 1552 6496 1558 6560
rect 1622 6496 1638 6560
rect 1702 6496 1718 6560
rect 1782 6496 1798 6560
rect 1862 6496 1868 6560
rect 1552 6495 1868 6496
rect 4652 6560 4968 6561
rect 4652 6496 4658 6560
rect 4722 6496 4738 6560
rect 4802 6496 4818 6560
rect 4882 6496 4898 6560
rect 4962 6496 4968 6560
rect 4652 6495 4968 6496
rect 7752 6560 8068 6561
rect 7752 6496 7758 6560
rect 7822 6496 7838 6560
rect 7902 6496 7918 6560
rect 7982 6496 7998 6560
rect 8062 6496 8068 6560
rect 7752 6495 8068 6496
rect 10852 6560 11168 6561
rect 10852 6496 10858 6560
rect 10922 6496 10938 6560
rect 11002 6496 11018 6560
rect 11082 6496 11098 6560
rect 11162 6496 11168 6560
rect 10852 6495 11168 6496
rect 13952 6560 14268 6561
rect 13952 6496 13958 6560
rect 14022 6496 14038 6560
rect 14102 6496 14118 6560
rect 14182 6496 14198 6560
rect 14262 6496 14268 6560
rect 13952 6495 14268 6496
rect 17052 6560 17368 6561
rect 17052 6496 17058 6560
rect 17122 6496 17138 6560
rect 17202 6496 17218 6560
rect 17282 6496 17298 6560
rect 17362 6496 17368 6560
rect 17052 6495 17368 6496
rect 18413 6354 18479 6357
rect 19200 6354 20000 6384
rect 18413 6352 20000 6354
rect 18413 6296 18418 6352
rect 18474 6296 20000 6352
rect 18413 6294 20000 6296
rect 18413 6291 18479 6294
rect 19200 6264 20000 6294
rect 3102 6016 3418 6017
rect 3102 5952 3108 6016
rect 3172 5952 3188 6016
rect 3252 5952 3268 6016
rect 3332 5952 3348 6016
rect 3412 5952 3418 6016
rect 3102 5951 3418 5952
rect 6202 6016 6518 6017
rect 6202 5952 6208 6016
rect 6272 5952 6288 6016
rect 6352 5952 6368 6016
rect 6432 5952 6448 6016
rect 6512 5952 6518 6016
rect 6202 5951 6518 5952
rect 9302 6016 9618 6017
rect 9302 5952 9308 6016
rect 9372 5952 9388 6016
rect 9452 5952 9468 6016
rect 9532 5952 9548 6016
rect 9612 5952 9618 6016
rect 9302 5951 9618 5952
rect 12402 6016 12718 6017
rect 12402 5952 12408 6016
rect 12472 5952 12488 6016
rect 12552 5952 12568 6016
rect 12632 5952 12648 6016
rect 12712 5952 12718 6016
rect 12402 5951 12718 5952
rect 15502 6016 15818 6017
rect 15502 5952 15508 6016
rect 15572 5952 15588 6016
rect 15652 5952 15668 6016
rect 15732 5952 15748 6016
rect 15812 5952 15818 6016
rect 15502 5951 15818 5952
rect 18602 6016 18918 6017
rect 18602 5952 18608 6016
rect 18672 5952 18688 6016
rect 18752 5952 18768 6016
rect 18832 5952 18848 6016
rect 18912 5952 18918 6016
rect 18602 5951 18918 5952
rect 1552 5472 1868 5473
rect 1552 5408 1558 5472
rect 1622 5408 1638 5472
rect 1702 5408 1718 5472
rect 1782 5408 1798 5472
rect 1862 5408 1868 5472
rect 1552 5407 1868 5408
rect 4652 5472 4968 5473
rect 4652 5408 4658 5472
rect 4722 5408 4738 5472
rect 4802 5408 4818 5472
rect 4882 5408 4898 5472
rect 4962 5408 4968 5472
rect 4652 5407 4968 5408
rect 7752 5472 8068 5473
rect 7752 5408 7758 5472
rect 7822 5408 7838 5472
rect 7902 5408 7918 5472
rect 7982 5408 7998 5472
rect 8062 5408 8068 5472
rect 7752 5407 8068 5408
rect 10852 5472 11168 5473
rect 10852 5408 10858 5472
rect 10922 5408 10938 5472
rect 11002 5408 11018 5472
rect 11082 5408 11098 5472
rect 11162 5408 11168 5472
rect 10852 5407 11168 5408
rect 13952 5472 14268 5473
rect 13952 5408 13958 5472
rect 14022 5408 14038 5472
rect 14102 5408 14118 5472
rect 14182 5408 14198 5472
rect 14262 5408 14268 5472
rect 13952 5407 14268 5408
rect 17052 5472 17368 5473
rect 17052 5408 17058 5472
rect 17122 5408 17138 5472
rect 17202 5408 17218 5472
rect 17282 5408 17298 5472
rect 17362 5408 17368 5472
rect 17052 5407 17368 5408
rect 3102 4928 3418 4929
rect 3102 4864 3108 4928
rect 3172 4864 3188 4928
rect 3252 4864 3268 4928
rect 3332 4864 3348 4928
rect 3412 4864 3418 4928
rect 3102 4863 3418 4864
rect 6202 4928 6518 4929
rect 6202 4864 6208 4928
rect 6272 4864 6288 4928
rect 6352 4864 6368 4928
rect 6432 4864 6448 4928
rect 6512 4864 6518 4928
rect 6202 4863 6518 4864
rect 9302 4928 9618 4929
rect 9302 4864 9308 4928
rect 9372 4864 9388 4928
rect 9452 4864 9468 4928
rect 9532 4864 9548 4928
rect 9612 4864 9618 4928
rect 9302 4863 9618 4864
rect 12402 4928 12718 4929
rect 12402 4864 12408 4928
rect 12472 4864 12488 4928
rect 12552 4864 12568 4928
rect 12632 4864 12648 4928
rect 12712 4864 12718 4928
rect 12402 4863 12718 4864
rect 15502 4928 15818 4929
rect 15502 4864 15508 4928
rect 15572 4864 15588 4928
rect 15652 4864 15668 4928
rect 15732 4864 15748 4928
rect 15812 4864 15818 4928
rect 15502 4863 15818 4864
rect 18602 4928 18918 4929
rect 18602 4864 18608 4928
rect 18672 4864 18688 4928
rect 18752 4864 18768 4928
rect 18832 4864 18848 4928
rect 18912 4864 18918 4928
rect 18602 4863 18918 4864
rect 1552 4384 1868 4385
rect 1552 4320 1558 4384
rect 1622 4320 1638 4384
rect 1702 4320 1718 4384
rect 1782 4320 1798 4384
rect 1862 4320 1868 4384
rect 1552 4319 1868 4320
rect 4652 4384 4968 4385
rect 4652 4320 4658 4384
rect 4722 4320 4738 4384
rect 4802 4320 4818 4384
rect 4882 4320 4898 4384
rect 4962 4320 4968 4384
rect 4652 4319 4968 4320
rect 7752 4384 8068 4385
rect 7752 4320 7758 4384
rect 7822 4320 7838 4384
rect 7902 4320 7918 4384
rect 7982 4320 7998 4384
rect 8062 4320 8068 4384
rect 7752 4319 8068 4320
rect 10852 4384 11168 4385
rect 10852 4320 10858 4384
rect 10922 4320 10938 4384
rect 11002 4320 11018 4384
rect 11082 4320 11098 4384
rect 11162 4320 11168 4384
rect 10852 4319 11168 4320
rect 13952 4384 14268 4385
rect 13952 4320 13958 4384
rect 14022 4320 14038 4384
rect 14102 4320 14118 4384
rect 14182 4320 14198 4384
rect 14262 4320 14268 4384
rect 13952 4319 14268 4320
rect 17052 4384 17368 4385
rect 17052 4320 17058 4384
rect 17122 4320 17138 4384
rect 17202 4320 17218 4384
rect 17282 4320 17298 4384
rect 17362 4320 17368 4384
rect 17052 4319 17368 4320
rect 19057 3906 19123 3909
rect 19200 3906 20000 3936
rect 19057 3904 20000 3906
rect 19057 3848 19062 3904
rect 19118 3848 20000 3904
rect 19057 3846 20000 3848
rect 19057 3843 19123 3846
rect 3102 3840 3418 3841
rect 3102 3776 3108 3840
rect 3172 3776 3188 3840
rect 3252 3776 3268 3840
rect 3332 3776 3348 3840
rect 3412 3776 3418 3840
rect 3102 3775 3418 3776
rect 6202 3840 6518 3841
rect 6202 3776 6208 3840
rect 6272 3776 6288 3840
rect 6352 3776 6368 3840
rect 6432 3776 6448 3840
rect 6512 3776 6518 3840
rect 6202 3775 6518 3776
rect 9302 3840 9618 3841
rect 9302 3776 9308 3840
rect 9372 3776 9388 3840
rect 9452 3776 9468 3840
rect 9532 3776 9548 3840
rect 9612 3776 9618 3840
rect 9302 3775 9618 3776
rect 12402 3840 12718 3841
rect 12402 3776 12408 3840
rect 12472 3776 12488 3840
rect 12552 3776 12568 3840
rect 12632 3776 12648 3840
rect 12712 3776 12718 3840
rect 12402 3775 12718 3776
rect 15502 3840 15818 3841
rect 15502 3776 15508 3840
rect 15572 3776 15588 3840
rect 15652 3776 15668 3840
rect 15732 3776 15748 3840
rect 15812 3776 15818 3840
rect 15502 3775 15818 3776
rect 18602 3840 18918 3841
rect 18602 3776 18608 3840
rect 18672 3776 18688 3840
rect 18752 3776 18768 3840
rect 18832 3776 18848 3840
rect 18912 3776 18918 3840
rect 19200 3816 20000 3846
rect 18602 3775 18918 3776
rect 1552 3296 1868 3297
rect 1552 3232 1558 3296
rect 1622 3232 1638 3296
rect 1702 3232 1718 3296
rect 1782 3232 1798 3296
rect 1862 3232 1868 3296
rect 1552 3231 1868 3232
rect 4652 3296 4968 3297
rect 4652 3232 4658 3296
rect 4722 3232 4738 3296
rect 4802 3232 4818 3296
rect 4882 3232 4898 3296
rect 4962 3232 4968 3296
rect 4652 3231 4968 3232
rect 7752 3296 8068 3297
rect 7752 3232 7758 3296
rect 7822 3232 7838 3296
rect 7902 3232 7918 3296
rect 7982 3232 7998 3296
rect 8062 3232 8068 3296
rect 7752 3231 8068 3232
rect 10852 3296 11168 3297
rect 10852 3232 10858 3296
rect 10922 3232 10938 3296
rect 11002 3232 11018 3296
rect 11082 3232 11098 3296
rect 11162 3232 11168 3296
rect 10852 3231 11168 3232
rect 13952 3296 14268 3297
rect 13952 3232 13958 3296
rect 14022 3232 14038 3296
rect 14102 3232 14118 3296
rect 14182 3232 14198 3296
rect 14262 3232 14268 3296
rect 13952 3231 14268 3232
rect 17052 3296 17368 3297
rect 17052 3232 17058 3296
rect 17122 3232 17138 3296
rect 17202 3232 17218 3296
rect 17282 3232 17298 3296
rect 17362 3232 17368 3296
rect 17052 3231 17368 3232
rect 3102 2752 3418 2753
rect 3102 2688 3108 2752
rect 3172 2688 3188 2752
rect 3252 2688 3268 2752
rect 3332 2688 3348 2752
rect 3412 2688 3418 2752
rect 3102 2687 3418 2688
rect 6202 2752 6518 2753
rect 6202 2688 6208 2752
rect 6272 2688 6288 2752
rect 6352 2688 6368 2752
rect 6432 2688 6448 2752
rect 6512 2688 6518 2752
rect 6202 2687 6518 2688
rect 9302 2752 9618 2753
rect 9302 2688 9308 2752
rect 9372 2688 9388 2752
rect 9452 2688 9468 2752
rect 9532 2688 9548 2752
rect 9612 2688 9618 2752
rect 9302 2687 9618 2688
rect 12402 2752 12718 2753
rect 12402 2688 12408 2752
rect 12472 2688 12488 2752
rect 12552 2688 12568 2752
rect 12632 2688 12648 2752
rect 12712 2688 12718 2752
rect 12402 2687 12718 2688
rect 15502 2752 15818 2753
rect 15502 2688 15508 2752
rect 15572 2688 15588 2752
rect 15652 2688 15668 2752
rect 15732 2688 15748 2752
rect 15812 2688 15818 2752
rect 15502 2687 15818 2688
rect 18602 2752 18918 2753
rect 18602 2688 18608 2752
rect 18672 2688 18688 2752
rect 18752 2688 18768 2752
rect 18832 2688 18848 2752
rect 18912 2688 18918 2752
rect 18602 2687 18918 2688
rect 1552 2208 1868 2209
rect 1552 2144 1558 2208
rect 1622 2144 1638 2208
rect 1702 2144 1718 2208
rect 1782 2144 1798 2208
rect 1862 2144 1868 2208
rect 1552 2143 1868 2144
rect 4652 2208 4968 2209
rect 4652 2144 4658 2208
rect 4722 2144 4738 2208
rect 4802 2144 4818 2208
rect 4882 2144 4898 2208
rect 4962 2144 4968 2208
rect 4652 2143 4968 2144
rect 7752 2208 8068 2209
rect 7752 2144 7758 2208
rect 7822 2144 7838 2208
rect 7902 2144 7918 2208
rect 7982 2144 7998 2208
rect 8062 2144 8068 2208
rect 7752 2143 8068 2144
rect 10852 2208 11168 2209
rect 10852 2144 10858 2208
rect 10922 2144 10938 2208
rect 11002 2144 11018 2208
rect 11082 2144 11098 2208
rect 11162 2144 11168 2208
rect 10852 2143 11168 2144
rect 13952 2208 14268 2209
rect 13952 2144 13958 2208
rect 14022 2144 14038 2208
rect 14102 2144 14118 2208
rect 14182 2144 14198 2208
rect 14262 2144 14268 2208
rect 13952 2143 14268 2144
rect 17052 2208 17368 2209
rect 17052 2144 17058 2208
rect 17122 2144 17138 2208
rect 17202 2144 17218 2208
rect 17282 2144 17298 2208
rect 17362 2144 17368 2208
rect 17052 2143 17368 2144
rect 3102 1664 3418 1665
rect 3102 1600 3108 1664
rect 3172 1600 3188 1664
rect 3252 1600 3268 1664
rect 3332 1600 3348 1664
rect 3412 1600 3418 1664
rect 3102 1599 3418 1600
rect 6202 1664 6518 1665
rect 6202 1600 6208 1664
rect 6272 1600 6288 1664
rect 6352 1600 6368 1664
rect 6432 1600 6448 1664
rect 6512 1600 6518 1664
rect 6202 1599 6518 1600
rect 9302 1664 9618 1665
rect 9302 1600 9308 1664
rect 9372 1600 9388 1664
rect 9452 1600 9468 1664
rect 9532 1600 9548 1664
rect 9612 1600 9618 1664
rect 9302 1599 9618 1600
rect 12402 1664 12718 1665
rect 12402 1600 12408 1664
rect 12472 1600 12488 1664
rect 12552 1600 12568 1664
rect 12632 1600 12648 1664
rect 12712 1600 12718 1664
rect 12402 1599 12718 1600
rect 15502 1664 15818 1665
rect 15502 1600 15508 1664
rect 15572 1600 15588 1664
rect 15652 1600 15668 1664
rect 15732 1600 15748 1664
rect 15812 1600 15818 1664
rect 15502 1599 15818 1600
rect 18602 1664 18918 1665
rect 18602 1600 18608 1664
rect 18672 1600 18688 1664
rect 18752 1600 18768 1664
rect 18832 1600 18848 1664
rect 18912 1600 18918 1664
rect 18602 1599 18918 1600
rect 18413 1458 18479 1461
rect 19200 1458 20000 1488
rect 18413 1456 20000 1458
rect 18413 1400 18418 1456
rect 18474 1400 20000 1456
rect 18413 1398 20000 1400
rect 18413 1395 18479 1398
rect 19200 1368 20000 1398
rect 1552 1120 1868 1121
rect 1552 1056 1558 1120
rect 1622 1056 1638 1120
rect 1702 1056 1718 1120
rect 1782 1056 1798 1120
rect 1862 1056 1868 1120
rect 1552 1055 1868 1056
rect 4652 1120 4968 1121
rect 4652 1056 4658 1120
rect 4722 1056 4738 1120
rect 4802 1056 4818 1120
rect 4882 1056 4898 1120
rect 4962 1056 4968 1120
rect 4652 1055 4968 1056
rect 7752 1120 8068 1121
rect 7752 1056 7758 1120
rect 7822 1056 7838 1120
rect 7902 1056 7918 1120
rect 7982 1056 7998 1120
rect 8062 1056 8068 1120
rect 7752 1055 8068 1056
rect 10852 1120 11168 1121
rect 10852 1056 10858 1120
rect 10922 1056 10938 1120
rect 11002 1056 11018 1120
rect 11082 1056 11098 1120
rect 11162 1056 11168 1120
rect 10852 1055 11168 1056
rect 13952 1120 14268 1121
rect 13952 1056 13958 1120
rect 14022 1056 14038 1120
rect 14102 1056 14118 1120
rect 14182 1056 14198 1120
rect 14262 1056 14268 1120
rect 13952 1055 14268 1056
rect 17052 1120 17368 1121
rect 17052 1056 17058 1120
rect 17122 1056 17138 1120
rect 17202 1056 17218 1120
rect 17282 1056 17298 1120
rect 17362 1056 17368 1120
rect 17052 1055 17368 1056
rect 3102 576 3418 577
rect 3102 512 3108 576
rect 3172 512 3188 576
rect 3252 512 3268 576
rect 3332 512 3348 576
rect 3412 512 3418 576
rect 3102 511 3418 512
rect 6202 576 6518 577
rect 6202 512 6208 576
rect 6272 512 6288 576
rect 6352 512 6368 576
rect 6432 512 6448 576
rect 6512 512 6518 576
rect 6202 511 6518 512
rect 9302 576 9618 577
rect 9302 512 9308 576
rect 9372 512 9388 576
rect 9452 512 9468 576
rect 9532 512 9548 576
rect 9612 512 9618 576
rect 9302 511 9618 512
rect 12402 576 12718 577
rect 12402 512 12408 576
rect 12472 512 12488 576
rect 12552 512 12568 576
rect 12632 512 12648 576
rect 12712 512 12718 576
rect 12402 511 12718 512
rect 15502 576 15818 577
rect 15502 512 15508 576
rect 15572 512 15588 576
rect 15652 512 15668 576
rect 15732 512 15748 576
rect 15812 512 15818 576
rect 15502 511 15818 512
rect 18602 576 18918 577
rect 18602 512 18608 576
rect 18672 512 18688 576
rect 18752 512 18768 576
rect 18832 512 18848 576
rect 18912 512 18918 576
rect 18602 511 18918 512
<< via3 >>
rect 1558 18524 1622 18528
rect 1558 18468 1562 18524
rect 1562 18468 1618 18524
rect 1618 18468 1622 18524
rect 1558 18464 1622 18468
rect 1638 18524 1702 18528
rect 1638 18468 1642 18524
rect 1642 18468 1698 18524
rect 1698 18468 1702 18524
rect 1638 18464 1702 18468
rect 1718 18524 1782 18528
rect 1718 18468 1722 18524
rect 1722 18468 1778 18524
rect 1778 18468 1782 18524
rect 1718 18464 1782 18468
rect 1798 18524 1862 18528
rect 1798 18468 1802 18524
rect 1802 18468 1858 18524
rect 1858 18468 1862 18524
rect 1798 18464 1862 18468
rect 4658 18524 4722 18528
rect 4658 18468 4662 18524
rect 4662 18468 4718 18524
rect 4718 18468 4722 18524
rect 4658 18464 4722 18468
rect 4738 18524 4802 18528
rect 4738 18468 4742 18524
rect 4742 18468 4798 18524
rect 4798 18468 4802 18524
rect 4738 18464 4802 18468
rect 4818 18524 4882 18528
rect 4818 18468 4822 18524
rect 4822 18468 4878 18524
rect 4878 18468 4882 18524
rect 4818 18464 4882 18468
rect 4898 18524 4962 18528
rect 4898 18468 4902 18524
rect 4902 18468 4958 18524
rect 4958 18468 4962 18524
rect 4898 18464 4962 18468
rect 7758 18524 7822 18528
rect 7758 18468 7762 18524
rect 7762 18468 7818 18524
rect 7818 18468 7822 18524
rect 7758 18464 7822 18468
rect 7838 18524 7902 18528
rect 7838 18468 7842 18524
rect 7842 18468 7898 18524
rect 7898 18468 7902 18524
rect 7838 18464 7902 18468
rect 7918 18524 7982 18528
rect 7918 18468 7922 18524
rect 7922 18468 7978 18524
rect 7978 18468 7982 18524
rect 7918 18464 7982 18468
rect 7998 18524 8062 18528
rect 7998 18468 8002 18524
rect 8002 18468 8058 18524
rect 8058 18468 8062 18524
rect 7998 18464 8062 18468
rect 10858 18524 10922 18528
rect 10858 18468 10862 18524
rect 10862 18468 10918 18524
rect 10918 18468 10922 18524
rect 10858 18464 10922 18468
rect 10938 18524 11002 18528
rect 10938 18468 10942 18524
rect 10942 18468 10998 18524
rect 10998 18468 11002 18524
rect 10938 18464 11002 18468
rect 11018 18524 11082 18528
rect 11018 18468 11022 18524
rect 11022 18468 11078 18524
rect 11078 18468 11082 18524
rect 11018 18464 11082 18468
rect 11098 18524 11162 18528
rect 11098 18468 11102 18524
rect 11102 18468 11158 18524
rect 11158 18468 11162 18524
rect 11098 18464 11162 18468
rect 13958 18524 14022 18528
rect 13958 18468 13962 18524
rect 13962 18468 14018 18524
rect 14018 18468 14022 18524
rect 13958 18464 14022 18468
rect 14038 18524 14102 18528
rect 14038 18468 14042 18524
rect 14042 18468 14098 18524
rect 14098 18468 14102 18524
rect 14038 18464 14102 18468
rect 14118 18524 14182 18528
rect 14118 18468 14122 18524
rect 14122 18468 14178 18524
rect 14178 18468 14182 18524
rect 14118 18464 14182 18468
rect 14198 18524 14262 18528
rect 14198 18468 14202 18524
rect 14202 18468 14258 18524
rect 14258 18468 14262 18524
rect 14198 18464 14262 18468
rect 17058 18524 17122 18528
rect 17058 18468 17062 18524
rect 17062 18468 17118 18524
rect 17118 18468 17122 18524
rect 17058 18464 17122 18468
rect 17138 18524 17202 18528
rect 17138 18468 17142 18524
rect 17142 18468 17198 18524
rect 17198 18468 17202 18524
rect 17138 18464 17202 18468
rect 17218 18524 17282 18528
rect 17218 18468 17222 18524
rect 17222 18468 17278 18524
rect 17278 18468 17282 18524
rect 17218 18464 17282 18468
rect 17298 18524 17362 18528
rect 17298 18468 17302 18524
rect 17302 18468 17358 18524
rect 17358 18468 17362 18524
rect 17298 18464 17362 18468
rect 3108 17980 3172 17984
rect 3108 17924 3112 17980
rect 3112 17924 3168 17980
rect 3168 17924 3172 17980
rect 3108 17920 3172 17924
rect 3188 17980 3252 17984
rect 3188 17924 3192 17980
rect 3192 17924 3248 17980
rect 3248 17924 3252 17980
rect 3188 17920 3252 17924
rect 3268 17980 3332 17984
rect 3268 17924 3272 17980
rect 3272 17924 3328 17980
rect 3328 17924 3332 17980
rect 3268 17920 3332 17924
rect 3348 17980 3412 17984
rect 3348 17924 3352 17980
rect 3352 17924 3408 17980
rect 3408 17924 3412 17980
rect 3348 17920 3412 17924
rect 6208 17980 6272 17984
rect 6208 17924 6212 17980
rect 6212 17924 6268 17980
rect 6268 17924 6272 17980
rect 6208 17920 6272 17924
rect 6288 17980 6352 17984
rect 6288 17924 6292 17980
rect 6292 17924 6348 17980
rect 6348 17924 6352 17980
rect 6288 17920 6352 17924
rect 6368 17980 6432 17984
rect 6368 17924 6372 17980
rect 6372 17924 6428 17980
rect 6428 17924 6432 17980
rect 6368 17920 6432 17924
rect 6448 17980 6512 17984
rect 6448 17924 6452 17980
rect 6452 17924 6508 17980
rect 6508 17924 6512 17980
rect 6448 17920 6512 17924
rect 9308 17980 9372 17984
rect 9308 17924 9312 17980
rect 9312 17924 9368 17980
rect 9368 17924 9372 17980
rect 9308 17920 9372 17924
rect 9388 17980 9452 17984
rect 9388 17924 9392 17980
rect 9392 17924 9448 17980
rect 9448 17924 9452 17980
rect 9388 17920 9452 17924
rect 9468 17980 9532 17984
rect 9468 17924 9472 17980
rect 9472 17924 9528 17980
rect 9528 17924 9532 17980
rect 9468 17920 9532 17924
rect 9548 17980 9612 17984
rect 9548 17924 9552 17980
rect 9552 17924 9608 17980
rect 9608 17924 9612 17980
rect 9548 17920 9612 17924
rect 12408 17980 12472 17984
rect 12408 17924 12412 17980
rect 12412 17924 12468 17980
rect 12468 17924 12472 17980
rect 12408 17920 12472 17924
rect 12488 17980 12552 17984
rect 12488 17924 12492 17980
rect 12492 17924 12548 17980
rect 12548 17924 12552 17980
rect 12488 17920 12552 17924
rect 12568 17980 12632 17984
rect 12568 17924 12572 17980
rect 12572 17924 12628 17980
rect 12628 17924 12632 17980
rect 12568 17920 12632 17924
rect 12648 17980 12712 17984
rect 12648 17924 12652 17980
rect 12652 17924 12708 17980
rect 12708 17924 12712 17980
rect 12648 17920 12712 17924
rect 15508 17980 15572 17984
rect 15508 17924 15512 17980
rect 15512 17924 15568 17980
rect 15568 17924 15572 17980
rect 15508 17920 15572 17924
rect 15588 17980 15652 17984
rect 15588 17924 15592 17980
rect 15592 17924 15648 17980
rect 15648 17924 15652 17980
rect 15588 17920 15652 17924
rect 15668 17980 15732 17984
rect 15668 17924 15672 17980
rect 15672 17924 15728 17980
rect 15728 17924 15732 17980
rect 15668 17920 15732 17924
rect 15748 17980 15812 17984
rect 15748 17924 15752 17980
rect 15752 17924 15808 17980
rect 15808 17924 15812 17980
rect 15748 17920 15812 17924
rect 18608 17980 18672 17984
rect 18608 17924 18612 17980
rect 18612 17924 18668 17980
rect 18668 17924 18672 17980
rect 18608 17920 18672 17924
rect 18688 17980 18752 17984
rect 18688 17924 18692 17980
rect 18692 17924 18748 17980
rect 18748 17924 18752 17980
rect 18688 17920 18752 17924
rect 18768 17980 18832 17984
rect 18768 17924 18772 17980
rect 18772 17924 18828 17980
rect 18828 17924 18832 17980
rect 18768 17920 18832 17924
rect 18848 17980 18912 17984
rect 18848 17924 18852 17980
rect 18852 17924 18908 17980
rect 18908 17924 18912 17980
rect 18848 17920 18912 17924
rect 1558 17436 1622 17440
rect 1558 17380 1562 17436
rect 1562 17380 1618 17436
rect 1618 17380 1622 17436
rect 1558 17376 1622 17380
rect 1638 17436 1702 17440
rect 1638 17380 1642 17436
rect 1642 17380 1698 17436
rect 1698 17380 1702 17436
rect 1638 17376 1702 17380
rect 1718 17436 1782 17440
rect 1718 17380 1722 17436
rect 1722 17380 1778 17436
rect 1778 17380 1782 17436
rect 1718 17376 1782 17380
rect 1798 17436 1862 17440
rect 1798 17380 1802 17436
rect 1802 17380 1858 17436
rect 1858 17380 1862 17436
rect 1798 17376 1862 17380
rect 4658 17436 4722 17440
rect 4658 17380 4662 17436
rect 4662 17380 4718 17436
rect 4718 17380 4722 17436
rect 4658 17376 4722 17380
rect 4738 17436 4802 17440
rect 4738 17380 4742 17436
rect 4742 17380 4798 17436
rect 4798 17380 4802 17436
rect 4738 17376 4802 17380
rect 4818 17436 4882 17440
rect 4818 17380 4822 17436
rect 4822 17380 4878 17436
rect 4878 17380 4882 17436
rect 4818 17376 4882 17380
rect 4898 17436 4962 17440
rect 4898 17380 4902 17436
rect 4902 17380 4958 17436
rect 4958 17380 4962 17436
rect 4898 17376 4962 17380
rect 7758 17436 7822 17440
rect 7758 17380 7762 17436
rect 7762 17380 7818 17436
rect 7818 17380 7822 17436
rect 7758 17376 7822 17380
rect 7838 17436 7902 17440
rect 7838 17380 7842 17436
rect 7842 17380 7898 17436
rect 7898 17380 7902 17436
rect 7838 17376 7902 17380
rect 7918 17436 7982 17440
rect 7918 17380 7922 17436
rect 7922 17380 7978 17436
rect 7978 17380 7982 17436
rect 7918 17376 7982 17380
rect 7998 17436 8062 17440
rect 7998 17380 8002 17436
rect 8002 17380 8058 17436
rect 8058 17380 8062 17436
rect 7998 17376 8062 17380
rect 10858 17436 10922 17440
rect 10858 17380 10862 17436
rect 10862 17380 10918 17436
rect 10918 17380 10922 17436
rect 10858 17376 10922 17380
rect 10938 17436 11002 17440
rect 10938 17380 10942 17436
rect 10942 17380 10998 17436
rect 10998 17380 11002 17436
rect 10938 17376 11002 17380
rect 11018 17436 11082 17440
rect 11018 17380 11022 17436
rect 11022 17380 11078 17436
rect 11078 17380 11082 17436
rect 11018 17376 11082 17380
rect 11098 17436 11162 17440
rect 11098 17380 11102 17436
rect 11102 17380 11158 17436
rect 11158 17380 11162 17436
rect 11098 17376 11162 17380
rect 13958 17436 14022 17440
rect 13958 17380 13962 17436
rect 13962 17380 14018 17436
rect 14018 17380 14022 17436
rect 13958 17376 14022 17380
rect 14038 17436 14102 17440
rect 14038 17380 14042 17436
rect 14042 17380 14098 17436
rect 14098 17380 14102 17436
rect 14038 17376 14102 17380
rect 14118 17436 14182 17440
rect 14118 17380 14122 17436
rect 14122 17380 14178 17436
rect 14178 17380 14182 17436
rect 14118 17376 14182 17380
rect 14198 17436 14262 17440
rect 14198 17380 14202 17436
rect 14202 17380 14258 17436
rect 14258 17380 14262 17436
rect 14198 17376 14262 17380
rect 17058 17436 17122 17440
rect 17058 17380 17062 17436
rect 17062 17380 17118 17436
rect 17118 17380 17122 17436
rect 17058 17376 17122 17380
rect 17138 17436 17202 17440
rect 17138 17380 17142 17436
rect 17142 17380 17198 17436
rect 17198 17380 17202 17436
rect 17138 17376 17202 17380
rect 17218 17436 17282 17440
rect 17218 17380 17222 17436
rect 17222 17380 17278 17436
rect 17278 17380 17282 17436
rect 17218 17376 17282 17380
rect 17298 17436 17362 17440
rect 17298 17380 17302 17436
rect 17302 17380 17358 17436
rect 17358 17380 17362 17436
rect 17298 17376 17362 17380
rect 3108 16892 3172 16896
rect 3108 16836 3112 16892
rect 3112 16836 3168 16892
rect 3168 16836 3172 16892
rect 3108 16832 3172 16836
rect 3188 16892 3252 16896
rect 3188 16836 3192 16892
rect 3192 16836 3248 16892
rect 3248 16836 3252 16892
rect 3188 16832 3252 16836
rect 3268 16892 3332 16896
rect 3268 16836 3272 16892
rect 3272 16836 3328 16892
rect 3328 16836 3332 16892
rect 3268 16832 3332 16836
rect 3348 16892 3412 16896
rect 3348 16836 3352 16892
rect 3352 16836 3408 16892
rect 3408 16836 3412 16892
rect 3348 16832 3412 16836
rect 6208 16892 6272 16896
rect 6208 16836 6212 16892
rect 6212 16836 6268 16892
rect 6268 16836 6272 16892
rect 6208 16832 6272 16836
rect 6288 16892 6352 16896
rect 6288 16836 6292 16892
rect 6292 16836 6348 16892
rect 6348 16836 6352 16892
rect 6288 16832 6352 16836
rect 6368 16892 6432 16896
rect 6368 16836 6372 16892
rect 6372 16836 6428 16892
rect 6428 16836 6432 16892
rect 6368 16832 6432 16836
rect 6448 16892 6512 16896
rect 6448 16836 6452 16892
rect 6452 16836 6508 16892
rect 6508 16836 6512 16892
rect 6448 16832 6512 16836
rect 9308 16892 9372 16896
rect 9308 16836 9312 16892
rect 9312 16836 9368 16892
rect 9368 16836 9372 16892
rect 9308 16832 9372 16836
rect 9388 16892 9452 16896
rect 9388 16836 9392 16892
rect 9392 16836 9448 16892
rect 9448 16836 9452 16892
rect 9388 16832 9452 16836
rect 9468 16892 9532 16896
rect 9468 16836 9472 16892
rect 9472 16836 9528 16892
rect 9528 16836 9532 16892
rect 9468 16832 9532 16836
rect 9548 16892 9612 16896
rect 9548 16836 9552 16892
rect 9552 16836 9608 16892
rect 9608 16836 9612 16892
rect 9548 16832 9612 16836
rect 12408 16892 12472 16896
rect 12408 16836 12412 16892
rect 12412 16836 12468 16892
rect 12468 16836 12472 16892
rect 12408 16832 12472 16836
rect 12488 16892 12552 16896
rect 12488 16836 12492 16892
rect 12492 16836 12548 16892
rect 12548 16836 12552 16892
rect 12488 16832 12552 16836
rect 12568 16892 12632 16896
rect 12568 16836 12572 16892
rect 12572 16836 12628 16892
rect 12628 16836 12632 16892
rect 12568 16832 12632 16836
rect 12648 16892 12712 16896
rect 12648 16836 12652 16892
rect 12652 16836 12708 16892
rect 12708 16836 12712 16892
rect 12648 16832 12712 16836
rect 15508 16892 15572 16896
rect 15508 16836 15512 16892
rect 15512 16836 15568 16892
rect 15568 16836 15572 16892
rect 15508 16832 15572 16836
rect 15588 16892 15652 16896
rect 15588 16836 15592 16892
rect 15592 16836 15648 16892
rect 15648 16836 15652 16892
rect 15588 16832 15652 16836
rect 15668 16892 15732 16896
rect 15668 16836 15672 16892
rect 15672 16836 15728 16892
rect 15728 16836 15732 16892
rect 15668 16832 15732 16836
rect 15748 16892 15812 16896
rect 15748 16836 15752 16892
rect 15752 16836 15808 16892
rect 15808 16836 15812 16892
rect 15748 16832 15812 16836
rect 18608 16892 18672 16896
rect 18608 16836 18612 16892
rect 18612 16836 18668 16892
rect 18668 16836 18672 16892
rect 18608 16832 18672 16836
rect 18688 16892 18752 16896
rect 18688 16836 18692 16892
rect 18692 16836 18748 16892
rect 18748 16836 18752 16892
rect 18688 16832 18752 16836
rect 18768 16892 18832 16896
rect 18768 16836 18772 16892
rect 18772 16836 18828 16892
rect 18828 16836 18832 16892
rect 18768 16832 18832 16836
rect 18848 16892 18912 16896
rect 18848 16836 18852 16892
rect 18852 16836 18908 16892
rect 18908 16836 18912 16892
rect 18848 16832 18912 16836
rect 1558 16348 1622 16352
rect 1558 16292 1562 16348
rect 1562 16292 1618 16348
rect 1618 16292 1622 16348
rect 1558 16288 1622 16292
rect 1638 16348 1702 16352
rect 1638 16292 1642 16348
rect 1642 16292 1698 16348
rect 1698 16292 1702 16348
rect 1638 16288 1702 16292
rect 1718 16348 1782 16352
rect 1718 16292 1722 16348
rect 1722 16292 1778 16348
rect 1778 16292 1782 16348
rect 1718 16288 1782 16292
rect 1798 16348 1862 16352
rect 1798 16292 1802 16348
rect 1802 16292 1858 16348
rect 1858 16292 1862 16348
rect 1798 16288 1862 16292
rect 4658 16348 4722 16352
rect 4658 16292 4662 16348
rect 4662 16292 4718 16348
rect 4718 16292 4722 16348
rect 4658 16288 4722 16292
rect 4738 16348 4802 16352
rect 4738 16292 4742 16348
rect 4742 16292 4798 16348
rect 4798 16292 4802 16348
rect 4738 16288 4802 16292
rect 4818 16348 4882 16352
rect 4818 16292 4822 16348
rect 4822 16292 4878 16348
rect 4878 16292 4882 16348
rect 4818 16288 4882 16292
rect 4898 16348 4962 16352
rect 4898 16292 4902 16348
rect 4902 16292 4958 16348
rect 4958 16292 4962 16348
rect 4898 16288 4962 16292
rect 7758 16348 7822 16352
rect 7758 16292 7762 16348
rect 7762 16292 7818 16348
rect 7818 16292 7822 16348
rect 7758 16288 7822 16292
rect 7838 16348 7902 16352
rect 7838 16292 7842 16348
rect 7842 16292 7898 16348
rect 7898 16292 7902 16348
rect 7838 16288 7902 16292
rect 7918 16348 7982 16352
rect 7918 16292 7922 16348
rect 7922 16292 7978 16348
rect 7978 16292 7982 16348
rect 7918 16288 7982 16292
rect 7998 16348 8062 16352
rect 7998 16292 8002 16348
rect 8002 16292 8058 16348
rect 8058 16292 8062 16348
rect 7998 16288 8062 16292
rect 10858 16348 10922 16352
rect 10858 16292 10862 16348
rect 10862 16292 10918 16348
rect 10918 16292 10922 16348
rect 10858 16288 10922 16292
rect 10938 16348 11002 16352
rect 10938 16292 10942 16348
rect 10942 16292 10998 16348
rect 10998 16292 11002 16348
rect 10938 16288 11002 16292
rect 11018 16348 11082 16352
rect 11018 16292 11022 16348
rect 11022 16292 11078 16348
rect 11078 16292 11082 16348
rect 11018 16288 11082 16292
rect 11098 16348 11162 16352
rect 11098 16292 11102 16348
rect 11102 16292 11158 16348
rect 11158 16292 11162 16348
rect 11098 16288 11162 16292
rect 13958 16348 14022 16352
rect 13958 16292 13962 16348
rect 13962 16292 14018 16348
rect 14018 16292 14022 16348
rect 13958 16288 14022 16292
rect 14038 16348 14102 16352
rect 14038 16292 14042 16348
rect 14042 16292 14098 16348
rect 14098 16292 14102 16348
rect 14038 16288 14102 16292
rect 14118 16348 14182 16352
rect 14118 16292 14122 16348
rect 14122 16292 14178 16348
rect 14178 16292 14182 16348
rect 14118 16288 14182 16292
rect 14198 16348 14262 16352
rect 14198 16292 14202 16348
rect 14202 16292 14258 16348
rect 14258 16292 14262 16348
rect 14198 16288 14262 16292
rect 17058 16348 17122 16352
rect 17058 16292 17062 16348
rect 17062 16292 17118 16348
rect 17118 16292 17122 16348
rect 17058 16288 17122 16292
rect 17138 16348 17202 16352
rect 17138 16292 17142 16348
rect 17142 16292 17198 16348
rect 17198 16292 17202 16348
rect 17138 16288 17202 16292
rect 17218 16348 17282 16352
rect 17218 16292 17222 16348
rect 17222 16292 17278 16348
rect 17278 16292 17282 16348
rect 17218 16288 17282 16292
rect 17298 16348 17362 16352
rect 17298 16292 17302 16348
rect 17302 16292 17358 16348
rect 17358 16292 17362 16348
rect 17298 16288 17362 16292
rect 3108 15804 3172 15808
rect 3108 15748 3112 15804
rect 3112 15748 3168 15804
rect 3168 15748 3172 15804
rect 3108 15744 3172 15748
rect 3188 15804 3252 15808
rect 3188 15748 3192 15804
rect 3192 15748 3248 15804
rect 3248 15748 3252 15804
rect 3188 15744 3252 15748
rect 3268 15804 3332 15808
rect 3268 15748 3272 15804
rect 3272 15748 3328 15804
rect 3328 15748 3332 15804
rect 3268 15744 3332 15748
rect 3348 15804 3412 15808
rect 3348 15748 3352 15804
rect 3352 15748 3408 15804
rect 3408 15748 3412 15804
rect 3348 15744 3412 15748
rect 6208 15804 6272 15808
rect 6208 15748 6212 15804
rect 6212 15748 6268 15804
rect 6268 15748 6272 15804
rect 6208 15744 6272 15748
rect 6288 15804 6352 15808
rect 6288 15748 6292 15804
rect 6292 15748 6348 15804
rect 6348 15748 6352 15804
rect 6288 15744 6352 15748
rect 6368 15804 6432 15808
rect 6368 15748 6372 15804
rect 6372 15748 6428 15804
rect 6428 15748 6432 15804
rect 6368 15744 6432 15748
rect 6448 15804 6512 15808
rect 6448 15748 6452 15804
rect 6452 15748 6508 15804
rect 6508 15748 6512 15804
rect 6448 15744 6512 15748
rect 9308 15804 9372 15808
rect 9308 15748 9312 15804
rect 9312 15748 9368 15804
rect 9368 15748 9372 15804
rect 9308 15744 9372 15748
rect 9388 15804 9452 15808
rect 9388 15748 9392 15804
rect 9392 15748 9448 15804
rect 9448 15748 9452 15804
rect 9388 15744 9452 15748
rect 9468 15804 9532 15808
rect 9468 15748 9472 15804
rect 9472 15748 9528 15804
rect 9528 15748 9532 15804
rect 9468 15744 9532 15748
rect 9548 15804 9612 15808
rect 9548 15748 9552 15804
rect 9552 15748 9608 15804
rect 9608 15748 9612 15804
rect 9548 15744 9612 15748
rect 12408 15804 12472 15808
rect 12408 15748 12412 15804
rect 12412 15748 12468 15804
rect 12468 15748 12472 15804
rect 12408 15744 12472 15748
rect 12488 15804 12552 15808
rect 12488 15748 12492 15804
rect 12492 15748 12548 15804
rect 12548 15748 12552 15804
rect 12488 15744 12552 15748
rect 12568 15804 12632 15808
rect 12568 15748 12572 15804
rect 12572 15748 12628 15804
rect 12628 15748 12632 15804
rect 12568 15744 12632 15748
rect 12648 15804 12712 15808
rect 12648 15748 12652 15804
rect 12652 15748 12708 15804
rect 12708 15748 12712 15804
rect 12648 15744 12712 15748
rect 15508 15804 15572 15808
rect 15508 15748 15512 15804
rect 15512 15748 15568 15804
rect 15568 15748 15572 15804
rect 15508 15744 15572 15748
rect 15588 15804 15652 15808
rect 15588 15748 15592 15804
rect 15592 15748 15648 15804
rect 15648 15748 15652 15804
rect 15588 15744 15652 15748
rect 15668 15804 15732 15808
rect 15668 15748 15672 15804
rect 15672 15748 15728 15804
rect 15728 15748 15732 15804
rect 15668 15744 15732 15748
rect 15748 15804 15812 15808
rect 15748 15748 15752 15804
rect 15752 15748 15808 15804
rect 15808 15748 15812 15804
rect 15748 15744 15812 15748
rect 18608 15804 18672 15808
rect 18608 15748 18612 15804
rect 18612 15748 18668 15804
rect 18668 15748 18672 15804
rect 18608 15744 18672 15748
rect 18688 15804 18752 15808
rect 18688 15748 18692 15804
rect 18692 15748 18748 15804
rect 18748 15748 18752 15804
rect 18688 15744 18752 15748
rect 18768 15804 18832 15808
rect 18768 15748 18772 15804
rect 18772 15748 18828 15804
rect 18828 15748 18832 15804
rect 18768 15744 18832 15748
rect 18848 15804 18912 15808
rect 18848 15748 18852 15804
rect 18852 15748 18908 15804
rect 18908 15748 18912 15804
rect 18848 15744 18912 15748
rect 1558 15260 1622 15264
rect 1558 15204 1562 15260
rect 1562 15204 1618 15260
rect 1618 15204 1622 15260
rect 1558 15200 1622 15204
rect 1638 15260 1702 15264
rect 1638 15204 1642 15260
rect 1642 15204 1698 15260
rect 1698 15204 1702 15260
rect 1638 15200 1702 15204
rect 1718 15260 1782 15264
rect 1718 15204 1722 15260
rect 1722 15204 1778 15260
rect 1778 15204 1782 15260
rect 1718 15200 1782 15204
rect 1798 15260 1862 15264
rect 1798 15204 1802 15260
rect 1802 15204 1858 15260
rect 1858 15204 1862 15260
rect 1798 15200 1862 15204
rect 4658 15260 4722 15264
rect 4658 15204 4662 15260
rect 4662 15204 4718 15260
rect 4718 15204 4722 15260
rect 4658 15200 4722 15204
rect 4738 15260 4802 15264
rect 4738 15204 4742 15260
rect 4742 15204 4798 15260
rect 4798 15204 4802 15260
rect 4738 15200 4802 15204
rect 4818 15260 4882 15264
rect 4818 15204 4822 15260
rect 4822 15204 4878 15260
rect 4878 15204 4882 15260
rect 4818 15200 4882 15204
rect 4898 15260 4962 15264
rect 4898 15204 4902 15260
rect 4902 15204 4958 15260
rect 4958 15204 4962 15260
rect 4898 15200 4962 15204
rect 7758 15260 7822 15264
rect 7758 15204 7762 15260
rect 7762 15204 7818 15260
rect 7818 15204 7822 15260
rect 7758 15200 7822 15204
rect 7838 15260 7902 15264
rect 7838 15204 7842 15260
rect 7842 15204 7898 15260
rect 7898 15204 7902 15260
rect 7838 15200 7902 15204
rect 7918 15260 7982 15264
rect 7918 15204 7922 15260
rect 7922 15204 7978 15260
rect 7978 15204 7982 15260
rect 7918 15200 7982 15204
rect 7998 15260 8062 15264
rect 7998 15204 8002 15260
rect 8002 15204 8058 15260
rect 8058 15204 8062 15260
rect 7998 15200 8062 15204
rect 10858 15260 10922 15264
rect 10858 15204 10862 15260
rect 10862 15204 10918 15260
rect 10918 15204 10922 15260
rect 10858 15200 10922 15204
rect 10938 15260 11002 15264
rect 10938 15204 10942 15260
rect 10942 15204 10998 15260
rect 10998 15204 11002 15260
rect 10938 15200 11002 15204
rect 11018 15260 11082 15264
rect 11018 15204 11022 15260
rect 11022 15204 11078 15260
rect 11078 15204 11082 15260
rect 11018 15200 11082 15204
rect 11098 15260 11162 15264
rect 11098 15204 11102 15260
rect 11102 15204 11158 15260
rect 11158 15204 11162 15260
rect 11098 15200 11162 15204
rect 13958 15260 14022 15264
rect 13958 15204 13962 15260
rect 13962 15204 14018 15260
rect 14018 15204 14022 15260
rect 13958 15200 14022 15204
rect 14038 15260 14102 15264
rect 14038 15204 14042 15260
rect 14042 15204 14098 15260
rect 14098 15204 14102 15260
rect 14038 15200 14102 15204
rect 14118 15260 14182 15264
rect 14118 15204 14122 15260
rect 14122 15204 14178 15260
rect 14178 15204 14182 15260
rect 14118 15200 14182 15204
rect 14198 15260 14262 15264
rect 14198 15204 14202 15260
rect 14202 15204 14258 15260
rect 14258 15204 14262 15260
rect 14198 15200 14262 15204
rect 17058 15260 17122 15264
rect 17058 15204 17062 15260
rect 17062 15204 17118 15260
rect 17118 15204 17122 15260
rect 17058 15200 17122 15204
rect 17138 15260 17202 15264
rect 17138 15204 17142 15260
rect 17142 15204 17198 15260
rect 17198 15204 17202 15260
rect 17138 15200 17202 15204
rect 17218 15260 17282 15264
rect 17218 15204 17222 15260
rect 17222 15204 17278 15260
rect 17278 15204 17282 15260
rect 17218 15200 17282 15204
rect 17298 15260 17362 15264
rect 17298 15204 17302 15260
rect 17302 15204 17358 15260
rect 17358 15204 17362 15260
rect 17298 15200 17362 15204
rect 3108 14716 3172 14720
rect 3108 14660 3112 14716
rect 3112 14660 3168 14716
rect 3168 14660 3172 14716
rect 3108 14656 3172 14660
rect 3188 14716 3252 14720
rect 3188 14660 3192 14716
rect 3192 14660 3248 14716
rect 3248 14660 3252 14716
rect 3188 14656 3252 14660
rect 3268 14716 3332 14720
rect 3268 14660 3272 14716
rect 3272 14660 3328 14716
rect 3328 14660 3332 14716
rect 3268 14656 3332 14660
rect 3348 14716 3412 14720
rect 3348 14660 3352 14716
rect 3352 14660 3408 14716
rect 3408 14660 3412 14716
rect 3348 14656 3412 14660
rect 6208 14716 6272 14720
rect 6208 14660 6212 14716
rect 6212 14660 6268 14716
rect 6268 14660 6272 14716
rect 6208 14656 6272 14660
rect 6288 14716 6352 14720
rect 6288 14660 6292 14716
rect 6292 14660 6348 14716
rect 6348 14660 6352 14716
rect 6288 14656 6352 14660
rect 6368 14716 6432 14720
rect 6368 14660 6372 14716
rect 6372 14660 6428 14716
rect 6428 14660 6432 14716
rect 6368 14656 6432 14660
rect 6448 14716 6512 14720
rect 6448 14660 6452 14716
rect 6452 14660 6508 14716
rect 6508 14660 6512 14716
rect 6448 14656 6512 14660
rect 9308 14716 9372 14720
rect 9308 14660 9312 14716
rect 9312 14660 9368 14716
rect 9368 14660 9372 14716
rect 9308 14656 9372 14660
rect 9388 14716 9452 14720
rect 9388 14660 9392 14716
rect 9392 14660 9448 14716
rect 9448 14660 9452 14716
rect 9388 14656 9452 14660
rect 9468 14716 9532 14720
rect 9468 14660 9472 14716
rect 9472 14660 9528 14716
rect 9528 14660 9532 14716
rect 9468 14656 9532 14660
rect 9548 14716 9612 14720
rect 9548 14660 9552 14716
rect 9552 14660 9608 14716
rect 9608 14660 9612 14716
rect 9548 14656 9612 14660
rect 12408 14716 12472 14720
rect 12408 14660 12412 14716
rect 12412 14660 12468 14716
rect 12468 14660 12472 14716
rect 12408 14656 12472 14660
rect 12488 14716 12552 14720
rect 12488 14660 12492 14716
rect 12492 14660 12548 14716
rect 12548 14660 12552 14716
rect 12488 14656 12552 14660
rect 12568 14716 12632 14720
rect 12568 14660 12572 14716
rect 12572 14660 12628 14716
rect 12628 14660 12632 14716
rect 12568 14656 12632 14660
rect 12648 14716 12712 14720
rect 12648 14660 12652 14716
rect 12652 14660 12708 14716
rect 12708 14660 12712 14716
rect 12648 14656 12712 14660
rect 15508 14716 15572 14720
rect 15508 14660 15512 14716
rect 15512 14660 15568 14716
rect 15568 14660 15572 14716
rect 15508 14656 15572 14660
rect 15588 14716 15652 14720
rect 15588 14660 15592 14716
rect 15592 14660 15648 14716
rect 15648 14660 15652 14716
rect 15588 14656 15652 14660
rect 15668 14716 15732 14720
rect 15668 14660 15672 14716
rect 15672 14660 15728 14716
rect 15728 14660 15732 14716
rect 15668 14656 15732 14660
rect 15748 14716 15812 14720
rect 15748 14660 15752 14716
rect 15752 14660 15808 14716
rect 15808 14660 15812 14716
rect 15748 14656 15812 14660
rect 18608 14716 18672 14720
rect 18608 14660 18612 14716
rect 18612 14660 18668 14716
rect 18668 14660 18672 14716
rect 18608 14656 18672 14660
rect 18688 14716 18752 14720
rect 18688 14660 18692 14716
rect 18692 14660 18748 14716
rect 18748 14660 18752 14716
rect 18688 14656 18752 14660
rect 18768 14716 18832 14720
rect 18768 14660 18772 14716
rect 18772 14660 18828 14716
rect 18828 14660 18832 14716
rect 18768 14656 18832 14660
rect 18848 14716 18912 14720
rect 18848 14660 18852 14716
rect 18852 14660 18908 14716
rect 18908 14660 18912 14716
rect 18848 14656 18912 14660
rect 1558 14172 1622 14176
rect 1558 14116 1562 14172
rect 1562 14116 1618 14172
rect 1618 14116 1622 14172
rect 1558 14112 1622 14116
rect 1638 14172 1702 14176
rect 1638 14116 1642 14172
rect 1642 14116 1698 14172
rect 1698 14116 1702 14172
rect 1638 14112 1702 14116
rect 1718 14172 1782 14176
rect 1718 14116 1722 14172
rect 1722 14116 1778 14172
rect 1778 14116 1782 14172
rect 1718 14112 1782 14116
rect 1798 14172 1862 14176
rect 1798 14116 1802 14172
rect 1802 14116 1858 14172
rect 1858 14116 1862 14172
rect 1798 14112 1862 14116
rect 4658 14172 4722 14176
rect 4658 14116 4662 14172
rect 4662 14116 4718 14172
rect 4718 14116 4722 14172
rect 4658 14112 4722 14116
rect 4738 14172 4802 14176
rect 4738 14116 4742 14172
rect 4742 14116 4798 14172
rect 4798 14116 4802 14172
rect 4738 14112 4802 14116
rect 4818 14172 4882 14176
rect 4818 14116 4822 14172
rect 4822 14116 4878 14172
rect 4878 14116 4882 14172
rect 4818 14112 4882 14116
rect 4898 14172 4962 14176
rect 4898 14116 4902 14172
rect 4902 14116 4958 14172
rect 4958 14116 4962 14172
rect 4898 14112 4962 14116
rect 7758 14172 7822 14176
rect 7758 14116 7762 14172
rect 7762 14116 7818 14172
rect 7818 14116 7822 14172
rect 7758 14112 7822 14116
rect 7838 14172 7902 14176
rect 7838 14116 7842 14172
rect 7842 14116 7898 14172
rect 7898 14116 7902 14172
rect 7838 14112 7902 14116
rect 7918 14172 7982 14176
rect 7918 14116 7922 14172
rect 7922 14116 7978 14172
rect 7978 14116 7982 14172
rect 7918 14112 7982 14116
rect 7998 14172 8062 14176
rect 7998 14116 8002 14172
rect 8002 14116 8058 14172
rect 8058 14116 8062 14172
rect 7998 14112 8062 14116
rect 10858 14172 10922 14176
rect 10858 14116 10862 14172
rect 10862 14116 10918 14172
rect 10918 14116 10922 14172
rect 10858 14112 10922 14116
rect 10938 14172 11002 14176
rect 10938 14116 10942 14172
rect 10942 14116 10998 14172
rect 10998 14116 11002 14172
rect 10938 14112 11002 14116
rect 11018 14172 11082 14176
rect 11018 14116 11022 14172
rect 11022 14116 11078 14172
rect 11078 14116 11082 14172
rect 11018 14112 11082 14116
rect 11098 14172 11162 14176
rect 11098 14116 11102 14172
rect 11102 14116 11158 14172
rect 11158 14116 11162 14172
rect 11098 14112 11162 14116
rect 13958 14172 14022 14176
rect 13958 14116 13962 14172
rect 13962 14116 14018 14172
rect 14018 14116 14022 14172
rect 13958 14112 14022 14116
rect 14038 14172 14102 14176
rect 14038 14116 14042 14172
rect 14042 14116 14098 14172
rect 14098 14116 14102 14172
rect 14038 14112 14102 14116
rect 14118 14172 14182 14176
rect 14118 14116 14122 14172
rect 14122 14116 14178 14172
rect 14178 14116 14182 14172
rect 14118 14112 14182 14116
rect 14198 14172 14262 14176
rect 14198 14116 14202 14172
rect 14202 14116 14258 14172
rect 14258 14116 14262 14172
rect 14198 14112 14262 14116
rect 17058 14172 17122 14176
rect 17058 14116 17062 14172
rect 17062 14116 17118 14172
rect 17118 14116 17122 14172
rect 17058 14112 17122 14116
rect 17138 14172 17202 14176
rect 17138 14116 17142 14172
rect 17142 14116 17198 14172
rect 17198 14116 17202 14172
rect 17138 14112 17202 14116
rect 17218 14172 17282 14176
rect 17218 14116 17222 14172
rect 17222 14116 17278 14172
rect 17278 14116 17282 14172
rect 17218 14112 17282 14116
rect 17298 14172 17362 14176
rect 17298 14116 17302 14172
rect 17302 14116 17358 14172
rect 17358 14116 17362 14172
rect 17298 14112 17362 14116
rect 3108 13628 3172 13632
rect 3108 13572 3112 13628
rect 3112 13572 3168 13628
rect 3168 13572 3172 13628
rect 3108 13568 3172 13572
rect 3188 13628 3252 13632
rect 3188 13572 3192 13628
rect 3192 13572 3248 13628
rect 3248 13572 3252 13628
rect 3188 13568 3252 13572
rect 3268 13628 3332 13632
rect 3268 13572 3272 13628
rect 3272 13572 3328 13628
rect 3328 13572 3332 13628
rect 3268 13568 3332 13572
rect 3348 13628 3412 13632
rect 3348 13572 3352 13628
rect 3352 13572 3408 13628
rect 3408 13572 3412 13628
rect 3348 13568 3412 13572
rect 6208 13628 6272 13632
rect 6208 13572 6212 13628
rect 6212 13572 6268 13628
rect 6268 13572 6272 13628
rect 6208 13568 6272 13572
rect 6288 13628 6352 13632
rect 6288 13572 6292 13628
rect 6292 13572 6348 13628
rect 6348 13572 6352 13628
rect 6288 13568 6352 13572
rect 6368 13628 6432 13632
rect 6368 13572 6372 13628
rect 6372 13572 6428 13628
rect 6428 13572 6432 13628
rect 6368 13568 6432 13572
rect 6448 13628 6512 13632
rect 6448 13572 6452 13628
rect 6452 13572 6508 13628
rect 6508 13572 6512 13628
rect 6448 13568 6512 13572
rect 9308 13628 9372 13632
rect 9308 13572 9312 13628
rect 9312 13572 9368 13628
rect 9368 13572 9372 13628
rect 9308 13568 9372 13572
rect 9388 13628 9452 13632
rect 9388 13572 9392 13628
rect 9392 13572 9448 13628
rect 9448 13572 9452 13628
rect 9388 13568 9452 13572
rect 9468 13628 9532 13632
rect 9468 13572 9472 13628
rect 9472 13572 9528 13628
rect 9528 13572 9532 13628
rect 9468 13568 9532 13572
rect 9548 13628 9612 13632
rect 9548 13572 9552 13628
rect 9552 13572 9608 13628
rect 9608 13572 9612 13628
rect 9548 13568 9612 13572
rect 12408 13628 12472 13632
rect 12408 13572 12412 13628
rect 12412 13572 12468 13628
rect 12468 13572 12472 13628
rect 12408 13568 12472 13572
rect 12488 13628 12552 13632
rect 12488 13572 12492 13628
rect 12492 13572 12548 13628
rect 12548 13572 12552 13628
rect 12488 13568 12552 13572
rect 12568 13628 12632 13632
rect 12568 13572 12572 13628
rect 12572 13572 12628 13628
rect 12628 13572 12632 13628
rect 12568 13568 12632 13572
rect 12648 13628 12712 13632
rect 12648 13572 12652 13628
rect 12652 13572 12708 13628
rect 12708 13572 12712 13628
rect 12648 13568 12712 13572
rect 15508 13628 15572 13632
rect 15508 13572 15512 13628
rect 15512 13572 15568 13628
rect 15568 13572 15572 13628
rect 15508 13568 15572 13572
rect 15588 13628 15652 13632
rect 15588 13572 15592 13628
rect 15592 13572 15648 13628
rect 15648 13572 15652 13628
rect 15588 13568 15652 13572
rect 15668 13628 15732 13632
rect 15668 13572 15672 13628
rect 15672 13572 15728 13628
rect 15728 13572 15732 13628
rect 15668 13568 15732 13572
rect 15748 13628 15812 13632
rect 15748 13572 15752 13628
rect 15752 13572 15808 13628
rect 15808 13572 15812 13628
rect 15748 13568 15812 13572
rect 18608 13628 18672 13632
rect 18608 13572 18612 13628
rect 18612 13572 18668 13628
rect 18668 13572 18672 13628
rect 18608 13568 18672 13572
rect 18688 13628 18752 13632
rect 18688 13572 18692 13628
rect 18692 13572 18748 13628
rect 18748 13572 18752 13628
rect 18688 13568 18752 13572
rect 18768 13628 18832 13632
rect 18768 13572 18772 13628
rect 18772 13572 18828 13628
rect 18828 13572 18832 13628
rect 18768 13568 18832 13572
rect 18848 13628 18912 13632
rect 18848 13572 18852 13628
rect 18852 13572 18908 13628
rect 18908 13572 18912 13628
rect 18848 13568 18912 13572
rect 1558 13084 1622 13088
rect 1558 13028 1562 13084
rect 1562 13028 1618 13084
rect 1618 13028 1622 13084
rect 1558 13024 1622 13028
rect 1638 13084 1702 13088
rect 1638 13028 1642 13084
rect 1642 13028 1698 13084
rect 1698 13028 1702 13084
rect 1638 13024 1702 13028
rect 1718 13084 1782 13088
rect 1718 13028 1722 13084
rect 1722 13028 1778 13084
rect 1778 13028 1782 13084
rect 1718 13024 1782 13028
rect 1798 13084 1862 13088
rect 1798 13028 1802 13084
rect 1802 13028 1858 13084
rect 1858 13028 1862 13084
rect 1798 13024 1862 13028
rect 4658 13084 4722 13088
rect 4658 13028 4662 13084
rect 4662 13028 4718 13084
rect 4718 13028 4722 13084
rect 4658 13024 4722 13028
rect 4738 13084 4802 13088
rect 4738 13028 4742 13084
rect 4742 13028 4798 13084
rect 4798 13028 4802 13084
rect 4738 13024 4802 13028
rect 4818 13084 4882 13088
rect 4818 13028 4822 13084
rect 4822 13028 4878 13084
rect 4878 13028 4882 13084
rect 4818 13024 4882 13028
rect 4898 13084 4962 13088
rect 4898 13028 4902 13084
rect 4902 13028 4958 13084
rect 4958 13028 4962 13084
rect 4898 13024 4962 13028
rect 7758 13084 7822 13088
rect 7758 13028 7762 13084
rect 7762 13028 7818 13084
rect 7818 13028 7822 13084
rect 7758 13024 7822 13028
rect 7838 13084 7902 13088
rect 7838 13028 7842 13084
rect 7842 13028 7898 13084
rect 7898 13028 7902 13084
rect 7838 13024 7902 13028
rect 7918 13084 7982 13088
rect 7918 13028 7922 13084
rect 7922 13028 7978 13084
rect 7978 13028 7982 13084
rect 7918 13024 7982 13028
rect 7998 13084 8062 13088
rect 7998 13028 8002 13084
rect 8002 13028 8058 13084
rect 8058 13028 8062 13084
rect 7998 13024 8062 13028
rect 10858 13084 10922 13088
rect 10858 13028 10862 13084
rect 10862 13028 10918 13084
rect 10918 13028 10922 13084
rect 10858 13024 10922 13028
rect 10938 13084 11002 13088
rect 10938 13028 10942 13084
rect 10942 13028 10998 13084
rect 10998 13028 11002 13084
rect 10938 13024 11002 13028
rect 11018 13084 11082 13088
rect 11018 13028 11022 13084
rect 11022 13028 11078 13084
rect 11078 13028 11082 13084
rect 11018 13024 11082 13028
rect 11098 13084 11162 13088
rect 11098 13028 11102 13084
rect 11102 13028 11158 13084
rect 11158 13028 11162 13084
rect 11098 13024 11162 13028
rect 13958 13084 14022 13088
rect 13958 13028 13962 13084
rect 13962 13028 14018 13084
rect 14018 13028 14022 13084
rect 13958 13024 14022 13028
rect 14038 13084 14102 13088
rect 14038 13028 14042 13084
rect 14042 13028 14098 13084
rect 14098 13028 14102 13084
rect 14038 13024 14102 13028
rect 14118 13084 14182 13088
rect 14118 13028 14122 13084
rect 14122 13028 14178 13084
rect 14178 13028 14182 13084
rect 14118 13024 14182 13028
rect 14198 13084 14262 13088
rect 14198 13028 14202 13084
rect 14202 13028 14258 13084
rect 14258 13028 14262 13084
rect 14198 13024 14262 13028
rect 17058 13084 17122 13088
rect 17058 13028 17062 13084
rect 17062 13028 17118 13084
rect 17118 13028 17122 13084
rect 17058 13024 17122 13028
rect 17138 13084 17202 13088
rect 17138 13028 17142 13084
rect 17142 13028 17198 13084
rect 17198 13028 17202 13084
rect 17138 13024 17202 13028
rect 17218 13084 17282 13088
rect 17218 13028 17222 13084
rect 17222 13028 17278 13084
rect 17278 13028 17282 13084
rect 17218 13024 17282 13028
rect 17298 13084 17362 13088
rect 17298 13028 17302 13084
rect 17302 13028 17358 13084
rect 17358 13028 17362 13084
rect 17298 13024 17362 13028
rect 3108 12540 3172 12544
rect 3108 12484 3112 12540
rect 3112 12484 3168 12540
rect 3168 12484 3172 12540
rect 3108 12480 3172 12484
rect 3188 12540 3252 12544
rect 3188 12484 3192 12540
rect 3192 12484 3248 12540
rect 3248 12484 3252 12540
rect 3188 12480 3252 12484
rect 3268 12540 3332 12544
rect 3268 12484 3272 12540
rect 3272 12484 3328 12540
rect 3328 12484 3332 12540
rect 3268 12480 3332 12484
rect 3348 12540 3412 12544
rect 3348 12484 3352 12540
rect 3352 12484 3408 12540
rect 3408 12484 3412 12540
rect 3348 12480 3412 12484
rect 6208 12540 6272 12544
rect 6208 12484 6212 12540
rect 6212 12484 6268 12540
rect 6268 12484 6272 12540
rect 6208 12480 6272 12484
rect 6288 12540 6352 12544
rect 6288 12484 6292 12540
rect 6292 12484 6348 12540
rect 6348 12484 6352 12540
rect 6288 12480 6352 12484
rect 6368 12540 6432 12544
rect 6368 12484 6372 12540
rect 6372 12484 6428 12540
rect 6428 12484 6432 12540
rect 6368 12480 6432 12484
rect 6448 12540 6512 12544
rect 6448 12484 6452 12540
rect 6452 12484 6508 12540
rect 6508 12484 6512 12540
rect 6448 12480 6512 12484
rect 9308 12540 9372 12544
rect 9308 12484 9312 12540
rect 9312 12484 9368 12540
rect 9368 12484 9372 12540
rect 9308 12480 9372 12484
rect 9388 12540 9452 12544
rect 9388 12484 9392 12540
rect 9392 12484 9448 12540
rect 9448 12484 9452 12540
rect 9388 12480 9452 12484
rect 9468 12540 9532 12544
rect 9468 12484 9472 12540
rect 9472 12484 9528 12540
rect 9528 12484 9532 12540
rect 9468 12480 9532 12484
rect 9548 12540 9612 12544
rect 9548 12484 9552 12540
rect 9552 12484 9608 12540
rect 9608 12484 9612 12540
rect 9548 12480 9612 12484
rect 12408 12540 12472 12544
rect 12408 12484 12412 12540
rect 12412 12484 12468 12540
rect 12468 12484 12472 12540
rect 12408 12480 12472 12484
rect 12488 12540 12552 12544
rect 12488 12484 12492 12540
rect 12492 12484 12548 12540
rect 12548 12484 12552 12540
rect 12488 12480 12552 12484
rect 12568 12540 12632 12544
rect 12568 12484 12572 12540
rect 12572 12484 12628 12540
rect 12628 12484 12632 12540
rect 12568 12480 12632 12484
rect 12648 12540 12712 12544
rect 12648 12484 12652 12540
rect 12652 12484 12708 12540
rect 12708 12484 12712 12540
rect 12648 12480 12712 12484
rect 15508 12540 15572 12544
rect 15508 12484 15512 12540
rect 15512 12484 15568 12540
rect 15568 12484 15572 12540
rect 15508 12480 15572 12484
rect 15588 12540 15652 12544
rect 15588 12484 15592 12540
rect 15592 12484 15648 12540
rect 15648 12484 15652 12540
rect 15588 12480 15652 12484
rect 15668 12540 15732 12544
rect 15668 12484 15672 12540
rect 15672 12484 15728 12540
rect 15728 12484 15732 12540
rect 15668 12480 15732 12484
rect 15748 12540 15812 12544
rect 15748 12484 15752 12540
rect 15752 12484 15808 12540
rect 15808 12484 15812 12540
rect 15748 12480 15812 12484
rect 18608 12540 18672 12544
rect 18608 12484 18612 12540
rect 18612 12484 18668 12540
rect 18668 12484 18672 12540
rect 18608 12480 18672 12484
rect 18688 12540 18752 12544
rect 18688 12484 18692 12540
rect 18692 12484 18748 12540
rect 18748 12484 18752 12540
rect 18688 12480 18752 12484
rect 18768 12540 18832 12544
rect 18768 12484 18772 12540
rect 18772 12484 18828 12540
rect 18828 12484 18832 12540
rect 18768 12480 18832 12484
rect 18848 12540 18912 12544
rect 18848 12484 18852 12540
rect 18852 12484 18908 12540
rect 18908 12484 18912 12540
rect 18848 12480 18912 12484
rect 1558 11996 1622 12000
rect 1558 11940 1562 11996
rect 1562 11940 1618 11996
rect 1618 11940 1622 11996
rect 1558 11936 1622 11940
rect 1638 11996 1702 12000
rect 1638 11940 1642 11996
rect 1642 11940 1698 11996
rect 1698 11940 1702 11996
rect 1638 11936 1702 11940
rect 1718 11996 1782 12000
rect 1718 11940 1722 11996
rect 1722 11940 1778 11996
rect 1778 11940 1782 11996
rect 1718 11936 1782 11940
rect 1798 11996 1862 12000
rect 1798 11940 1802 11996
rect 1802 11940 1858 11996
rect 1858 11940 1862 11996
rect 1798 11936 1862 11940
rect 4658 11996 4722 12000
rect 4658 11940 4662 11996
rect 4662 11940 4718 11996
rect 4718 11940 4722 11996
rect 4658 11936 4722 11940
rect 4738 11996 4802 12000
rect 4738 11940 4742 11996
rect 4742 11940 4798 11996
rect 4798 11940 4802 11996
rect 4738 11936 4802 11940
rect 4818 11996 4882 12000
rect 4818 11940 4822 11996
rect 4822 11940 4878 11996
rect 4878 11940 4882 11996
rect 4818 11936 4882 11940
rect 4898 11996 4962 12000
rect 4898 11940 4902 11996
rect 4902 11940 4958 11996
rect 4958 11940 4962 11996
rect 4898 11936 4962 11940
rect 7758 11996 7822 12000
rect 7758 11940 7762 11996
rect 7762 11940 7818 11996
rect 7818 11940 7822 11996
rect 7758 11936 7822 11940
rect 7838 11996 7902 12000
rect 7838 11940 7842 11996
rect 7842 11940 7898 11996
rect 7898 11940 7902 11996
rect 7838 11936 7902 11940
rect 7918 11996 7982 12000
rect 7918 11940 7922 11996
rect 7922 11940 7978 11996
rect 7978 11940 7982 11996
rect 7918 11936 7982 11940
rect 7998 11996 8062 12000
rect 7998 11940 8002 11996
rect 8002 11940 8058 11996
rect 8058 11940 8062 11996
rect 7998 11936 8062 11940
rect 10858 11996 10922 12000
rect 10858 11940 10862 11996
rect 10862 11940 10918 11996
rect 10918 11940 10922 11996
rect 10858 11936 10922 11940
rect 10938 11996 11002 12000
rect 10938 11940 10942 11996
rect 10942 11940 10998 11996
rect 10998 11940 11002 11996
rect 10938 11936 11002 11940
rect 11018 11996 11082 12000
rect 11018 11940 11022 11996
rect 11022 11940 11078 11996
rect 11078 11940 11082 11996
rect 11018 11936 11082 11940
rect 11098 11996 11162 12000
rect 11098 11940 11102 11996
rect 11102 11940 11158 11996
rect 11158 11940 11162 11996
rect 11098 11936 11162 11940
rect 13958 11996 14022 12000
rect 13958 11940 13962 11996
rect 13962 11940 14018 11996
rect 14018 11940 14022 11996
rect 13958 11936 14022 11940
rect 14038 11996 14102 12000
rect 14038 11940 14042 11996
rect 14042 11940 14098 11996
rect 14098 11940 14102 11996
rect 14038 11936 14102 11940
rect 14118 11996 14182 12000
rect 14118 11940 14122 11996
rect 14122 11940 14178 11996
rect 14178 11940 14182 11996
rect 14118 11936 14182 11940
rect 14198 11996 14262 12000
rect 14198 11940 14202 11996
rect 14202 11940 14258 11996
rect 14258 11940 14262 11996
rect 14198 11936 14262 11940
rect 17058 11996 17122 12000
rect 17058 11940 17062 11996
rect 17062 11940 17118 11996
rect 17118 11940 17122 11996
rect 17058 11936 17122 11940
rect 17138 11996 17202 12000
rect 17138 11940 17142 11996
rect 17142 11940 17198 11996
rect 17198 11940 17202 11996
rect 17138 11936 17202 11940
rect 17218 11996 17282 12000
rect 17218 11940 17222 11996
rect 17222 11940 17278 11996
rect 17278 11940 17282 11996
rect 17218 11936 17282 11940
rect 17298 11996 17362 12000
rect 17298 11940 17302 11996
rect 17302 11940 17358 11996
rect 17358 11940 17362 11996
rect 17298 11936 17362 11940
rect 3108 11452 3172 11456
rect 3108 11396 3112 11452
rect 3112 11396 3168 11452
rect 3168 11396 3172 11452
rect 3108 11392 3172 11396
rect 3188 11452 3252 11456
rect 3188 11396 3192 11452
rect 3192 11396 3248 11452
rect 3248 11396 3252 11452
rect 3188 11392 3252 11396
rect 3268 11452 3332 11456
rect 3268 11396 3272 11452
rect 3272 11396 3328 11452
rect 3328 11396 3332 11452
rect 3268 11392 3332 11396
rect 3348 11452 3412 11456
rect 3348 11396 3352 11452
rect 3352 11396 3408 11452
rect 3408 11396 3412 11452
rect 3348 11392 3412 11396
rect 6208 11452 6272 11456
rect 6208 11396 6212 11452
rect 6212 11396 6268 11452
rect 6268 11396 6272 11452
rect 6208 11392 6272 11396
rect 6288 11452 6352 11456
rect 6288 11396 6292 11452
rect 6292 11396 6348 11452
rect 6348 11396 6352 11452
rect 6288 11392 6352 11396
rect 6368 11452 6432 11456
rect 6368 11396 6372 11452
rect 6372 11396 6428 11452
rect 6428 11396 6432 11452
rect 6368 11392 6432 11396
rect 6448 11452 6512 11456
rect 6448 11396 6452 11452
rect 6452 11396 6508 11452
rect 6508 11396 6512 11452
rect 6448 11392 6512 11396
rect 9308 11452 9372 11456
rect 9308 11396 9312 11452
rect 9312 11396 9368 11452
rect 9368 11396 9372 11452
rect 9308 11392 9372 11396
rect 9388 11452 9452 11456
rect 9388 11396 9392 11452
rect 9392 11396 9448 11452
rect 9448 11396 9452 11452
rect 9388 11392 9452 11396
rect 9468 11452 9532 11456
rect 9468 11396 9472 11452
rect 9472 11396 9528 11452
rect 9528 11396 9532 11452
rect 9468 11392 9532 11396
rect 9548 11452 9612 11456
rect 9548 11396 9552 11452
rect 9552 11396 9608 11452
rect 9608 11396 9612 11452
rect 9548 11392 9612 11396
rect 12408 11452 12472 11456
rect 12408 11396 12412 11452
rect 12412 11396 12468 11452
rect 12468 11396 12472 11452
rect 12408 11392 12472 11396
rect 12488 11452 12552 11456
rect 12488 11396 12492 11452
rect 12492 11396 12548 11452
rect 12548 11396 12552 11452
rect 12488 11392 12552 11396
rect 12568 11452 12632 11456
rect 12568 11396 12572 11452
rect 12572 11396 12628 11452
rect 12628 11396 12632 11452
rect 12568 11392 12632 11396
rect 12648 11452 12712 11456
rect 12648 11396 12652 11452
rect 12652 11396 12708 11452
rect 12708 11396 12712 11452
rect 12648 11392 12712 11396
rect 15508 11452 15572 11456
rect 15508 11396 15512 11452
rect 15512 11396 15568 11452
rect 15568 11396 15572 11452
rect 15508 11392 15572 11396
rect 15588 11452 15652 11456
rect 15588 11396 15592 11452
rect 15592 11396 15648 11452
rect 15648 11396 15652 11452
rect 15588 11392 15652 11396
rect 15668 11452 15732 11456
rect 15668 11396 15672 11452
rect 15672 11396 15728 11452
rect 15728 11396 15732 11452
rect 15668 11392 15732 11396
rect 15748 11452 15812 11456
rect 15748 11396 15752 11452
rect 15752 11396 15808 11452
rect 15808 11396 15812 11452
rect 15748 11392 15812 11396
rect 18608 11452 18672 11456
rect 18608 11396 18612 11452
rect 18612 11396 18668 11452
rect 18668 11396 18672 11452
rect 18608 11392 18672 11396
rect 18688 11452 18752 11456
rect 18688 11396 18692 11452
rect 18692 11396 18748 11452
rect 18748 11396 18752 11452
rect 18688 11392 18752 11396
rect 18768 11452 18832 11456
rect 18768 11396 18772 11452
rect 18772 11396 18828 11452
rect 18828 11396 18832 11452
rect 18768 11392 18832 11396
rect 18848 11452 18912 11456
rect 18848 11396 18852 11452
rect 18852 11396 18908 11452
rect 18908 11396 18912 11452
rect 18848 11392 18912 11396
rect 1558 10908 1622 10912
rect 1558 10852 1562 10908
rect 1562 10852 1618 10908
rect 1618 10852 1622 10908
rect 1558 10848 1622 10852
rect 1638 10908 1702 10912
rect 1638 10852 1642 10908
rect 1642 10852 1698 10908
rect 1698 10852 1702 10908
rect 1638 10848 1702 10852
rect 1718 10908 1782 10912
rect 1718 10852 1722 10908
rect 1722 10852 1778 10908
rect 1778 10852 1782 10908
rect 1718 10848 1782 10852
rect 1798 10908 1862 10912
rect 1798 10852 1802 10908
rect 1802 10852 1858 10908
rect 1858 10852 1862 10908
rect 1798 10848 1862 10852
rect 4658 10908 4722 10912
rect 4658 10852 4662 10908
rect 4662 10852 4718 10908
rect 4718 10852 4722 10908
rect 4658 10848 4722 10852
rect 4738 10908 4802 10912
rect 4738 10852 4742 10908
rect 4742 10852 4798 10908
rect 4798 10852 4802 10908
rect 4738 10848 4802 10852
rect 4818 10908 4882 10912
rect 4818 10852 4822 10908
rect 4822 10852 4878 10908
rect 4878 10852 4882 10908
rect 4818 10848 4882 10852
rect 4898 10908 4962 10912
rect 4898 10852 4902 10908
rect 4902 10852 4958 10908
rect 4958 10852 4962 10908
rect 4898 10848 4962 10852
rect 7758 10908 7822 10912
rect 7758 10852 7762 10908
rect 7762 10852 7818 10908
rect 7818 10852 7822 10908
rect 7758 10848 7822 10852
rect 7838 10908 7902 10912
rect 7838 10852 7842 10908
rect 7842 10852 7898 10908
rect 7898 10852 7902 10908
rect 7838 10848 7902 10852
rect 7918 10908 7982 10912
rect 7918 10852 7922 10908
rect 7922 10852 7978 10908
rect 7978 10852 7982 10908
rect 7918 10848 7982 10852
rect 7998 10908 8062 10912
rect 7998 10852 8002 10908
rect 8002 10852 8058 10908
rect 8058 10852 8062 10908
rect 7998 10848 8062 10852
rect 10858 10908 10922 10912
rect 10858 10852 10862 10908
rect 10862 10852 10918 10908
rect 10918 10852 10922 10908
rect 10858 10848 10922 10852
rect 10938 10908 11002 10912
rect 10938 10852 10942 10908
rect 10942 10852 10998 10908
rect 10998 10852 11002 10908
rect 10938 10848 11002 10852
rect 11018 10908 11082 10912
rect 11018 10852 11022 10908
rect 11022 10852 11078 10908
rect 11078 10852 11082 10908
rect 11018 10848 11082 10852
rect 11098 10908 11162 10912
rect 11098 10852 11102 10908
rect 11102 10852 11158 10908
rect 11158 10852 11162 10908
rect 11098 10848 11162 10852
rect 13958 10908 14022 10912
rect 13958 10852 13962 10908
rect 13962 10852 14018 10908
rect 14018 10852 14022 10908
rect 13958 10848 14022 10852
rect 14038 10908 14102 10912
rect 14038 10852 14042 10908
rect 14042 10852 14098 10908
rect 14098 10852 14102 10908
rect 14038 10848 14102 10852
rect 14118 10908 14182 10912
rect 14118 10852 14122 10908
rect 14122 10852 14178 10908
rect 14178 10852 14182 10908
rect 14118 10848 14182 10852
rect 14198 10908 14262 10912
rect 14198 10852 14202 10908
rect 14202 10852 14258 10908
rect 14258 10852 14262 10908
rect 14198 10848 14262 10852
rect 17058 10908 17122 10912
rect 17058 10852 17062 10908
rect 17062 10852 17118 10908
rect 17118 10852 17122 10908
rect 17058 10848 17122 10852
rect 17138 10908 17202 10912
rect 17138 10852 17142 10908
rect 17142 10852 17198 10908
rect 17198 10852 17202 10908
rect 17138 10848 17202 10852
rect 17218 10908 17282 10912
rect 17218 10852 17222 10908
rect 17222 10852 17278 10908
rect 17278 10852 17282 10908
rect 17218 10848 17282 10852
rect 17298 10908 17362 10912
rect 17298 10852 17302 10908
rect 17302 10852 17358 10908
rect 17358 10852 17362 10908
rect 17298 10848 17362 10852
rect 3108 10364 3172 10368
rect 3108 10308 3112 10364
rect 3112 10308 3168 10364
rect 3168 10308 3172 10364
rect 3108 10304 3172 10308
rect 3188 10364 3252 10368
rect 3188 10308 3192 10364
rect 3192 10308 3248 10364
rect 3248 10308 3252 10364
rect 3188 10304 3252 10308
rect 3268 10364 3332 10368
rect 3268 10308 3272 10364
rect 3272 10308 3328 10364
rect 3328 10308 3332 10364
rect 3268 10304 3332 10308
rect 3348 10364 3412 10368
rect 3348 10308 3352 10364
rect 3352 10308 3408 10364
rect 3408 10308 3412 10364
rect 3348 10304 3412 10308
rect 6208 10364 6272 10368
rect 6208 10308 6212 10364
rect 6212 10308 6268 10364
rect 6268 10308 6272 10364
rect 6208 10304 6272 10308
rect 6288 10364 6352 10368
rect 6288 10308 6292 10364
rect 6292 10308 6348 10364
rect 6348 10308 6352 10364
rect 6288 10304 6352 10308
rect 6368 10364 6432 10368
rect 6368 10308 6372 10364
rect 6372 10308 6428 10364
rect 6428 10308 6432 10364
rect 6368 10304 6432 10308
rect 6448 10364 6512 10368
rect 6448 10308 6452 10364
rect 6452 10308 6508 10364
rect 6508 10308 6512 10364
rect 6448 10304 6512 10308
rect 9308 10364 9372 10368
rect 9308 10308 9312 10364
rect 9312 10308 9368 10364
rect 9368 10308 9372 10364
rect 9308 10304 9372 10308
rect 9388 10364 9452 10368
rect 9388 10308 9392 10364
rect 9392 10308 9448 10364
rect 9448 10308 9452 10364
rect 9388 10304 9452 10308
rect 9468 10364 9532 10368
rect 9468 10308 9472 10364
rect 9472 10308 9528 10364
rect 9528 10308 9532 10364
rect 9468 10304 9532 10308
rect 9548 10364 9612 10368
rect 9548 10308 9552 10364
rect 9552 10308 9608 10364
rect 9608 10308 9612 10364
rect 9548 10304 9612 10308
rect 12408 10364 12472 10368
rect 12408 10308 12412 10364
rect 12412 10308 12468 10364
rect 12468 10308 12472 10364
rect 12408 10304 12472 10308
rect 12488 10364 12552 10368
rect 12488 10308 12492 10364
rect 12492 10308 12548 10364
rect 12548 10308 12552 10364
rect 12488 10304 12552 10308
rect 12568 10364 12632 10368
rect 12568 10308 12572 10364
rect 12572 10308 12628 10364
rect 12628 10308 12632 10364
rect 12568 10304 12632 10308
rect 12648 10364 12712 10368
rect 12648 10308 12652 10364
rect 12652 10308 12708 10364
rect 12708 10308 12712 10364
rect 12648 10304 12712 10308
rect 15508 10364 15572 10368
rect 15508 10308 15512 10364
rect 15512 10308 15568 10364
rect 15568 10308 15572 10364
rect 15508 10304 15572 10308
rect 15588 10364 15652 10368
rect 15588 10308 15592 10364
rect 15592 10308 15648 10364
rect 15648 10308 15652 10364
rect 15588 10304 15652 10308
rect 15668 10364 15732 10368
rect 15668 10308 15672 10364
rect 15672 10308 15728 10364
rect 15728 10308 15732 10364
rect 15668 10304 15732 10308
rect 15748 10364 15812 10368
rect 15748 10308 15752 10364
rect 15752 10308 15808 10364
rect 15808 10308 15812 10364
rect 15748 10304 15812 10308
rect 18608 10364 18672 10368
rect 18608 10308 18612 10364
rect 18612 10308 18668 10364
rect 18668 10308 18672 10364
rect 18608 10304 18672 10308
rect 18688 10364 18752 10368
rect 18688 10308 18692 10364
rect 18692 10308 18748 10364
rect 18748 10308 18752 10364
rect 18688 10304 18752 10308
rect 18768 10364 18832 10368
rect 18768 10308 18772 10364
rect 18772 10308 18828 10364
rect 18828 10308 18832 10364
rect 18768 10304 18832 10308
rect 18848 10364 18912 10368
rect 18848 10308 18852 10364
rect 18852 10308 18908 10364
rect 18908 10308 18912 10364
rect 18848 10304 18912 10308
rect 1558 9820 1622 9824
rect 1558 9764 1562 9820
rect 1562 9764 1618 9820
rect 1618 9764 1622 9820
rect 1558 9760 1622 9764
rect 1638 9820 1702 9824
rect 1638 9764 1642 9820
rect 1642 9764 1698 9820
rect 1698 9764 1702 9820
rect 1638 9760 1702 9764
rect 1718 9820 1782 9824
rect 1718 9764 1722 9820
rect 1722 9764 1778 9820
rect 1778 9764 1782 9820
rect 1718 9760 1782 9764
rect 1798 9820 1862 9824
rect 1798 9764 1802 9820
rect 1802 9764 1858 9820
rect 1858 9764 1862 9820
rect 1798 9760 1862 9764
rect 4658 9820 4722 9824
rect 4658 9764 4662 9820
rect 4662 9764 4718 9820
rect 4718 9764 4722 9820
rect 4658 9760 4722 9764
rect 4738 9820 4802 9824
rect 4738 9764 4742 9820
rect 4742 9764 4798 9820
rect 4798 9764 4802 9820
rect 4738 9760 4802 9764
rect 4818 9820 4882 9824
rect 4818 9764 4822 9820
rect 4822 9764 4878 9820
rect 4878 9764 4882 9820
rect 4818 9760 4882 9764
rect 4898 9820 4962 9824
rect 4898 9764 4902 9820
rect 4902 9764 4958 9820
rect 4958 9764 4962 9820
rect 4898 9760 4962 9764
rect 7758 9820 7822 9824
rect 7758 9764 7762 9820
rect 7762 9764 7818 9820
rect 7818 9764 7822 9820
rect 7758 9760 7822 9764
rect 7838 9820 7902 9824
rect 7838 9764 7842 9820
rect 7842 9764 7898 9820
rect 7898 9764 7902 9820
rect 7838 9760 7902 9764
rect 7918 9820 7982 9824
rect 7918 9764 7922 9820
rect 7922 9764 7978 9820
rect 7978 9764 7982 9820
rect 7918 9760 7982 9764
rect 7998 9820 8062 9824
rect 7998 9764 8002 9820
rect 8002 9764 8058 9820
rect 8058 9764 8062 9820
rect 7998 9760 8062 9764
rect 10858 9820 10922 9824
rect 10858 9764 10862 9820
rect 10862 9764 10918 9820
rect 10918 9764 10922 9820
rect 10858 9760 10922 9764
rect 10938 9820 11002 9824
rect 10938 9764 10942 9820
rect 10942 9764 10998 9820
rect 10998 9764 11002 9820
rect 10938 9760 11002 9764
rect 11018 9820 11082 9824
rect 11018 9764 11022 9820
rect 11022 9764 11078 9820
rect 11078 9764 11082 9820
rect 11018 9760 11082 9764
rect 11098 9820 11162 9824
rect 11098 9764 11102 9820
rect 11102 9764 11158 9820
rect 11158 9764 11162 9820
rect 11098 9760 11162 9764
rect 13958 9820 14022 9824
rect 13958 9764 13962 9820
rect 13962 9764 14018 9820
rect 14018 9764 14022 9820
rect 13958 9760 14022 9764
rect 14038 9820 14102 9824
rect 14038 9764 14042 9820
rect 14042 9764 14098 9820
rect 14098 9764 14102 9820
rect 14038 9760 14102 9764
rect 14118 9820 14182 9824
rect 14118 9764 14122 9820
rect 14122 9764 14178 9820
rect 14178 9764 14182 9820
rect 14118 9760 14182 9764
rect 14198 9820 14262 9824
rect 14198 9764 14202 9820
rect 14202 9764 14258 9820
rect 14258 9764 14262 9820
rect 14198 9760 14262 9764
rect 17058 9820 17122 9824
rect 17058 9764 17062 9820
rect 17062 9764 17118 9820
rect 17118 9764 17122 9820
rect 17058 9760 17122 9764
rect 17138 9820 17202 9824
rect 17138 9764 17142 9820
rect 17142 9764 17198 9820
rect 17198 9764 17202 9820
rect 17138 9760 17202 9764
rect 17218 9820 17282 9824
rect 17218 9764 17222 9820
rect 17222 9764 17278 9820
rect 17278 9764 17282 9820
rect 17218 9760 17282 9764
rect 17298 9820 17362 9824
rect 17298 9764 17302 9820
rect 17302 9764 17358 9820
rect 17358 9764 17362 9820
rect 17298 9760 17362 9764
rect 3108 9276 3172 9280
rect 3108 9220 3112 9276
rect 3112 9220 3168 9276
rect 3168 9220 3172 9276
rect 3108 9216 3172 9220
rect 3188 9276 3252 9280
rect 3188 9220 3192 9276
rect 3192 9220 3248 9276
rect 3248 9220 3252 9276
rect 3188 9216 3252 9220
rect 3268 9276 3332 9280
rect 3268 9220 3272 9276
rect 3272 9220 3328 9276
rect 3328 9220 3332 9276
rect 3268 9216 3332 9220
rect 3348 9276 3412 9280
rect 3348 9220 3352 9276
rect 3352 9220 3408 9276
rect 3408 9220 3412 9276
rect 3348 9216 3412 9220
rect 6208 9276 6272 9280
rect 6208 9220 6212 9276
rect 6212 9220 6268 9276
rect 6268 9220 6272 9276
rect 6208 9216 6272 9220
rect 6288 9276 6352 9280
rect 6288 9220 6292 9276
rect 6292 9220 6348 9276
rect 6348 9220 6352 9276
rect 6288 9216 6352 9220
rect 6368 9276 6432 9280
rect 6368 9220 6372 9276
rect 6372 9220 6428 9276
rect 6428 9220 6432 9276
rect 6368 9216 6432 9220
rect 6448 9276 6512 9280
rect 6448 9220 6452 9276
rect 6452 9220 6508 9276
rect 6508 9220 6512 9276
rect 6448 9216 6512 9220
rect 9308 9276 9372 9280
rect 9308 9220 9312 9276
rect 9312 9220 9368 9276
rect 9368 9220 9372 9276
rect 9308 9216 9372 9220
rect 9388 9276 9452 9280
rect 9388 9220 9392 9276
rect 9392 9220 9448 9276
rect 9448 9220 9452 9276
rect 9388 9216 9452 9220
rect 9468 9276 9532 9280
rect 9468 9220 9472 9276
rect 9472 9220 9528 9276
rect 9528 9220 9532 9276
rect 9468 9216 9532 9220
rect 9548 9276 9612 9280
rect 9548 9220 9552 9276
rect 9552 9220 9608 9276
rect 9608 9220 9612 9276
rect 9548 9216 9612 9220
rect 12408 9276 12472 9280
rect 12408 9220 12412 9276
rect 12412 9220 12468 9276
rect 12468 9220 12472 9276
rect 12408 9216 12472 9220
rect 12488 9276 12552 9280
rect 12488 9220 12492 9276
rect 12492 9220 12548 9276
rect 12548 9220 12552 9276
rect 12488 9216 12552 9220
rect 12568 9276 12632 9280
rect 12568 9220 12572 9276
rect 12572 9220 12628 9276
rect 12628 9220 12632 9276
rect 12568 9216 12632 9220
rect 12648 9276 12712 9280
rect 12648 9220 12652 9276
rect 12652 9220 12708 9276
rect 12708 9220 12712 9276
rect 12648 9216 12712 9220
rect 15508 9276 15572 9280
rect 15508 9220 15512 9276
rect 15512 9220 15568 9276
rect 15568 9220 15572 9276
rect 15508 9216 15572 9220
rect 15588 9276 15652 9280
rect 15588 9220 15592 9276
rect 15592 9220 15648 9276
rect 15648 9220 15652 9276
rect 15588 9216 15652 9220
rect 15668 9276 15732 9280
rect 15668 9220 15672 9276
rect 15672 9220 15728 9276
rect 15728 9220 15732 9276
rect 15668 9216 15732 9220
rect 15748 9276 15812 9280
rect 15748 9220 15752 9276
rect 15752 9220 15808 9276
rect 15808 9220 15812 9276
rect 15748 9216 15812 9220
rect 18608 9276 18672 9280
rect 18608 9220 18612 9276
rect 18612 9220 18668 9276
rect 18668 9220 18672 9276
rect 18608 9216 18672 9220
rect 18688 9276 18752 9280
rect 18688 9220 18692 9276
rect 18692 9220 18748 9276
rect 18748 9220 18752 9276
rect 18688 9216 18752 9220
rect 18768 9276 18832 9280
rect 18768 9220 18772 9276
rect 18772 9220 18828 9276
rect 18828 9220 18832 9276
rect 18768 9216 18832 9220
rect 18848 9276 18912 9280
rect 18848 9220 18852 9276
rect 18852 9220 18908 9276
rect 18908 9220 18912 9276
rect 18848 9216 18912 9220
rect 1558 8732 1622 8736
rect 1558 8676 1562 8732
rect 1562 8676 1618 8732
rect 1618 8676 1622 8732
rect 1558 8672 1622 8676
rect 1638 8732 1702 8736
rect 1638 8676 1642 8732
rect 1642 8676 1698 8732
rect 1698 8676 1702 8732
rect 1638 8672 1702 8676
rect 1718 8732 1782 8736
rect 1718 8676 1722 8732
rect 1722 8676 1778 8732
rect 1778 8676 1782 8732
rect 1718 8672 1782 8676
rect 1798 8732 1862 8736
rect 1798 8676 1802 8732
rect 1802 8676 1858 8732
rect 1858 8676 1862 8732
rect 1798 8672 1862 8676
rect 4658 8732 4722 8736
rect 4658 8676 4662 8732
rect 4662 8676 4718 8732
rect 4718 8676 4722 8732
rect 4658 8672 4722 8676
rect 4738 8732 4802 8736
rect 4738 8676 4742 8732
rect 4742 8676 4798 8732
rect 4798 8676 4802 8732
rect 4738 8672 4802 8676
rect 4818 8732 4882 8736
rect 4818 8676 4822 8732
rect 4822 8676 4878 8732
rect 4878 8676 4882 8732
rect 4818 8672 4882 8676
rect 4898 8732 4962 8736
rect 4898 8676 4902 8732
rect 4902 8676 4958 8732
rect 4958 8676 4962 8732
rect 4898 8672 4962 8676
rect 7758 8732 7822 8736
rect 7758 8676 7762 8732
rect 7762 8676 7818 8732
rect 7818 8676 7822 8732
rect 7758 8672 7822 8676
rect 7838 8732 7902 8736
rect 7838 8676 7842 8732
rect 7842 8676 7898 8732
rect 7898 8676 7902 8732
rect 7838 8672 7902 8676
rect 7918 8732 7982 8736
rect 7918 8676 7922 8732
rect 7922 8676 7978 8732
rect 7978 8676 7982 8732
rect 7918 8672 7982 8676
rect 7998 8732 8062 8736
rect 7998 8676 8002 8732
rect 8002 8676 8058 8732
rect 8058 8676 8062 8732
rect 7998 8672 8062 8676
rect 10858 8732 10922 8736
rect 10858 8676 10862 8732
rect 10862 8676 10918 8732
rect 10918 8676 10922 8732
rect 10858 8672 10922 8676
rect 10938 8732 11002 8736
rect 10938 8676 10942 8732
rect 10942 8676 10998 8732
rect 10998 8676 11002 8732
rect 10938 8672 11002 8676
rect 11018 8732 11082 8736
rect 11018 8676 11022 8732
rect 11022 8676 11078 8732
rect 11078 8676 11082 8732
rect 11018 8672 11082 8676
rect 11098 8732 11162 8736
rect 11098 8676 11102 8732
rect 11102 8676 11158 8732
rect 11158 8676 11162 8732
rect 11098 8672 11162 8676
rect 13958 8732 14022 8736
rect 13958 8676 13962 8732
rect 13962 8676 14018 8732
rect 14018 8676 14022 8732
rect 13958 8672 14022 8676
rect 14038 8732 14102 8736
rect 14038 8676 14042 8732
rect 14042 8676 14098 8732
rect 14098 8676 14102 8732
rect 14038 8672 14102 8676
rect 14118 8732 14182 8736
rect 14118 8676 14122 8732
rect 14122 8676 14178 8732
rect 14178 8676 14182 8732
rect 14118 8672 14182 8676
rect 14198 8732 14262 8736
rect 14198 8676 14202 8732
rect 14202 8676 14258 8732
rect 14258 8676 14262 8732
rect 14198 8672 14262 8676
rect 17058 8732 17122 8736
rect 17058 8676 17062 8732
rect 17062 8676 17118 8732
rect 17118 8676 17122 8732
rect 17058 8672 17122 8676
rect 17138 8732 17202 8736
rect 17138 8676 17142 8732
rect 17142 8676 17198 8732
rect 17198 8676 17202 8732
rect 17138 8672 17202 8676
rect 17218 8732 17282 8736
rect 17218 8676 17222 8732
rect 17222 8676 17278 8732
rect 17278 8676 17282 8732
rect 17218 8672 17282 8676
rect 17298 8732 17362 8736
rect 17298 8676 17302 8732
rect 17302 8676 17358 8732
rect 17358 8676 17362 8732
rect 17298 8672 17362 8676
rect 3108 8188 3172 8192
rect 3108 8132 3112 8188
rect 3112 8132 3168 8188
rect 3168 8132 3172 8188
rect 3108 8128 3172 8132
rect 3188 8188 3252 8192
rect 3188 8132 3192 8188
rect 3192 8132 3248 8188
rect 3248 8132 3252 8188
rect 3188 8128 3252 8132
rect 3268 8188 3332 8192
rect 3268 8132 3272 8188
rect 3272 8132 3328 8188
rect 3328 8132 3332 8188
rect 3268 8128 3332 8132
rect 3348 8188 3412 8192
rect 3348 8132 3352 8188
rect 3352 8132 3408 8188
rect 3408 8132 3412 8188
rect 3348 8128 3412 8132
rect 6208 8188 6272 8192
rect 6208 8132 6212 8188
rect 6212 8132 6268 8188
rect 6268 8132 6272 8188
rect 6208 8128 6272 8132
rect 6288 8188 6352 8192
rect 6288 8132 6292 8188
rect 6292 8132 6348 8188
rect 6348 8132 6352 8188
rect 6288 8128 6352 8132
rect 6368 8188 6432 8192
rect 6368 8132 6372 8188
rect 6372 8132 6428 8188
rect 6428 8132 6432 8188
rect 6368 8128 6432 8132
rect 6448 8188 6512 8192
rect 6448 8132 6452 8188
rect 6452 8132 6508 8188
rect 6508 8132 6512 8188
rect 6448 8128 6512 8132
rect 9308 8188 9372 8192
rect 9308 8132 9312 8188
rect 9312 8132 9368 8188
rect 9368 8132 9372 8188
rect 9308 8128 9372 8132
rect 9388 8188 9452 8192
rect 9388 8132 9392 8188
rect 9392 8132 9448 8188
rect 9448 8132 9452 8188
rect 9388 8128 9452 8132
rect 9468 8188 9532 8192
rect 9468 8132 9472 8188
rect 9472 8132 9528 8188
rect 9528 8132 9532 8188
rect 9468 8128 9532 8132
rect 9548 8188 9612 8192
rect 9548 8132 9552 8188
rect 9552 8132 9608 8188
rect 9608 8132 9612 8188
rect 9548 8128 9612 8132
rect 12408 8188 12472 8192
rect 12408 8132 12412 8188
rect 12412 8132 12468 8188
rect 12468 8132 12472 8188
rect 12408 8128 12472 8132
rect 12488 8188 12552 8192
rect 12488 8132 12492 8188
rect 12492 8132 12548 8188
rect 12548 8132 12552 8188
rect 12488 8128 12552 8132
rect 12568 8188 12632 8192
rect 12568 8132 12572 8188
rect 12572 8132 12628 8188
rect 12628 8132 12632 8188
rect 12568 8128 12632 8132
rect 12648 8188 12712 8192
rect 12648 8132 12652 8188
rect 12652 8132 12708 8188
rect 12708 8132 12712 8188
rect 12648 8128 12712 8132
rect 15508 8188 15572 8192
rect 15508 8132 15512 8188
rect 15512 8132 15568 8188
rect 15568 8132 15572 8188
rect 15508 8128 15572 8132
rect 15588 8188 15652 8192
rect 15588 8132 15592 8188
rect 15592 8132 15648 8188
rect 15648 8132 15652 8188
rect 15588 8128 15652 8132
rect 15668 8188 15732 8192
rect 15668 8132 15672 8188
rect 15672 8132 15728 8188
rect 15728 8132 15732 8188
rect 15668 8128 15732 8132
rect 15748 8188 15812 8192
rect 15748 8132 15752 8188
rect 15752 8132 15808 8188
rect 15808 8132 15812 8188
rect 15748 8128 15812 8132
rect 18608 8188 18672 8192
rect 18608 8132 18612 8188
rect 18612 8132 18668 8188
rect 18668 8132 18672 8188
rect 18608 8128 18672 8132
rect 18688 8188 18752 8192
rect 18688 8132 18692 8188
rect 18692 8132 18748 8188
rect 18748 8132 18752 8188
rect 18688 8128 18752 8132
rect 18768 8188 18832 8192
rect 18768 8132 18772 8188
rect 18772 8132 18828 8188
rect 18828 8132 18832 8188
rect 18768 8128 18832 8132
rect 18848 8188 18912 8192
rect 18848 8132 18852 8188
rect 18852 8132 18908 8188
rect 18908 8132 18912 8188
rect 18848 8128 18912 8132
rect 1558 7644 1622 7648
rect 1558 7588 1562 7644
rect 1562 7588 1618 7644
rect 1618 7588 1622 7644
rect 1558 7584 1622 7588
rect 1638 7644 1702 7648
rect 1638 7588 1642 7644
rect 1642 7588 1698 7644
rect 1698 7588 1702 7644
rect 1638 7584 1702 7588
rect 1718 7644 1782 7648
rect 1718 7588 1722 7644
rect 1722 7588 1778 7644
rect 1778 7588 1782 7644
rect 1718 7584 1782 7588
rect 1798 7644 1862 7648
rect 1798 7588 1802 7644
rect 1802 7588 1858 7644
rect 1858 7588 1862 7644
rect 1798 7584 1862 7588
rect 4658 7644 4722 7648
rect 4658 7588 4662 7644
rect 4662 7588 4718 7644
rect 4718 7588 4722 7644
rect 4658 7584 4722 7588
rect 4738 7644 4802 7648
rect 4738 7588 4742 7644
rect 4742 7588 4798 7644
rect 4798 7588 4802 7644
rect 4738 7584 4802 7588
rect 4818 7644 4882 7648
rect 4818 7588 4822 7644
rect 4822 7588 4878 7644
rect 4878 7588 4882 7644
rect 4818 7584 4882 7588
rect 4898 7644 4962 7648
rect 4898 7588 4902 7644
rect 4902 7588 4958 7644
rect 4958 7588 4962 7644
rect 4898 7584 4962 7588
rect 7758 7644 7822 7648
rect 7758 7588 7762 7644
rect 7762 7588 7818 7644
rect 7818 7588 7822 7644
rect 7758 7584 7822 7588
rect 7838 7644 7902 7648
rect 7838 7588 7842 7644
rect 7842 7588 7898 7644
rect 7898 7588 7902 7644
rect 7838 7584 7902 7588
rect 7918 7644 7982 7648
rect 7918 7588 7922 7644
rect 7922 7588 7978 7644
rect 7978 7588 7982 7644
rect 7918 7584 7982 7588
rect 7998 7644 8062 7648
rect 7998 7588 8002 7644
rect 8002 7588 8058 7644
rect 8058 7588 8062 7644
rect 7998 7584 8062 7588
rect 10858 7644 10922 7648
rect 10858 7588 10862 7644
rect 10862 7588 10918 7644
rect 10918 7588 10922 7644
rect 10858 7584 10922 7588
rect 10938 7644 11002 7648
rect 10938 7588 10942 7644
rect 10942 7588 10998 7644
rect 10998 7588 11002 7644
rect 10938 7584 11002 7588
rect 11018 7644 11082 7648
rect 11018 7588 11022 7644
rect 11022 7588 11078 7644
rect 11078 7588 11082 7644
rect 11018 7584 11082 7588
rect 11098 7644 11162 7648
rect 11098 7588 11102 7644
rect 11102 7588 11158 7644
rect 11158 7588 11162 7644
rect 11098 7584 11162 7588
rect 13958 7644 14022 7648
rect 13958 7588 13962 7644
rect 13962 7588 14018 7644
rect 14018 7588 14022 7644
rect 13958 7584 14022 7588
rect 14038 7644 14102 7648
rect 14038 7588 14042 7644
rect 14042 7588 14098 7644
rect 14098 7588 14102 7644
rect 14038 7584 14102 7588
rect 14118 7644 14182 7648
rect 14118 7588 14122 7644
rect 14122 7588 14178 7644
rect 14178 7588 14182 7644
rect 14118 7584 14182 7588
rect 14198 7644 14262 7648
rect 14198 7588 14202 7644
rect 14202 7588 14258 7644
rect 14258 7588 14262 7644
rect 14198 7584 14262 7588
rect 17058 7644 17122 7648
rect 17058 7588 17062 7644
rect 17062 7588 17118 7644
rect 17118 7588 17122 7644
rect 17058 7584 17122 7588
rect 17138 7644 17202 7648
rect 17138 7588 17142 7644
rect 17142 7588 17198 7644
rect 17198 7588 17202 7644
rect 17138 7584 17202 7588
rect 17218 7644 17282 7648
rect 17218 7588 17222 7644
rect 17222 7588 17278 7644
rect 17278 7588 17282 7644
rect 17218 7584 17282 7588
rect 17298 7644 17362 7648
rect 17298 7588 17302 7644
rect 17302 7588 17358 7644
rect 17358 7588 17362 7644
rect 17298 7584 17362 7588
rect 3108 7100 3172 7104
rect 3108 7044 3112 7100
rect 3112 7044 3168 7100
rect 3168 7044 3172 7100
rect 3108 7040 3172 7044
rect 3188 7100 3252 7104
rect 3188 7044 3192 7100
rect 3192 7044 3248 7100
rect 3248 7044 3252 7100
rect 3188 7040 3252 7044
rect 3268 7100 3332 7104
rect 3268 7044 3272 7100
rect 3272 7044 3328 7100
rect 3328 7044 3332 7100
rect 3268 7040 3332 7044
rect 3348 7100 3412 7104
rect 3348 7044 3352 7100
rect 3352 7044 3408 7100
rect 3408 7044 3412 7100
rect 3348 7040 3412 7044
rect 6208 7100 6272 7104
rect 6208 7044 6212 7100
rect 6212 7044 6268 7100
rect 6268 7044 6272 7100
rect 6208 7040 6272 7044
rect 6288 7100 6352 7104
rect 6288 7044 6292 7100
rect 6292 7044 6348 7100
rect 6348 7044 6352 7100
rect 6288 7040 6352 7044
rect 6368 7100 6432 7104
rect 6368 7044 6372 7100
rect 6372 7044 6428 7100
rect 6428 7044 6432 7100
rect 6368 7040 6432 7044
rect 6448 7100 6512 7104
rect 6448 7044 6452 7100
rect 6452 7044 6508 7100
rect 6508 7044 6512 7100
rect 6448 7040 6512 7044
rect 9308 7100 9372 7104
rect 9308 7044 9312 7100
rect 9312 7044 9368 7100
rect 9368 7044 9372 7100
rect 9308 7040 9372 7044
rect 9388 7100 9452 7104
rect 9388 7044 9392 7100
rect 9392 7044 9448 7100
rect 9448 7044 9452 7100
rect 9388 7040 9452 7044
rect 9468 7100 9532 7104
rect 9468 7044 9472 7100
rect 9472 7044 9528 7100
rect 9528 7044 9532 7100
rect 9468 7040 9532 7044
rect 9548 7100 9612 7104
rect 9548 7044 9552 7100
rect 9552 7044 9608 7100
rect 9608 7044 9612 7100
rect 9548 7040 9612 7044
rect 12408 7100 12472 7104
rect 12408 7044 12412 7100
rect 12412 7044 12468 7100
rect 12468 7044 12472 7100
rect 12408 7040 12472 7044
rect 12488 7100 12552 7104
rect 12488 7044 12492 7100
rect 12492 7044 12548 7100
rect 12548 7044 12552 7100
rect 12488 7040 12552 7044
rect 12568 7100 12632 7104
rect 12568 7044 12572 7100
rect 12572 7044 12628 7100
rect 12628 7044 12632 7100
rect 12568 7040 12632 7044
rect 12648 7100 12712 7104
rect 12648 7044 12652 7100
rect 12652 7044 12708 7100
rect 12708 7044 12712 7100
rect 12648 7040 12712 7044
rect 15508 7100 15572 7104
rect 15508 7044 15512 7100
rect 15512 7044 15568 7100
rect 15568 7044 15572 7100
rect 15508 7040 15572 7044
rect 15588 7100 15652 7104
rect 15588 7044 15592 7100
rect 15592 7044 15648 7100
rect 15648 7044 15652 7100
rect 15588 7040 15652 7044
rect 15668 7100 15732 7104
rect 15668 7044 15672 7100
rect 15672 7044 15728 7100
rect 15728 7044 15732 7100
rect 15668 7040 15732 7044
rect 15748 7100 15812 7104
rect 15748 7044 15752 7100
rect 15752 7044 15808 7100
rect 15808 7044 15812 7100
rect 15748 7040 15812 7044
rect 18608 7100 18672 7104
rect 18608 7044 18612 7100
rect 18612 7044 18668 7100
rect 18668 7044 18672 7100
rect 18608 7040 18672 7044
rect 18688 7100 18752 7104
rect 18688 7044 18692 7100
rect 18692 7044 18748 7100
rect 18748 7044 18752 7100
rect 18688 7040 18752 7044
rect 18768 7100 18832 7104
rect 18768 7044 18772 7100
rect 18772 7044 18828 7100
rect 18828 7044 18832 7100
rect 18768 7040 18832 7044
rect 18848 7100 18912 7104
rect 18848 7044 18852 7100
rect 18852 7044 18908 7100
rect 18908 7044 18912 7100
rect 18848 7040 18912 7044
rect 1558 6556 1622 6560
rect 1558 6500 1562 6556
rect 1562 6500 1618 6556
rect 1618 6500 1622 6556
rect 1558 6496 1622 6500
rect 1638 6556 1702 6560
rect 1638 6500 1642 6556
rect 1642 6500 1698 6556
rect 1698 6500 1702 6556
rect 1638 6496 1702 6500
rect 1718 6556 1782 6560
rect 1718 6500 1722 6556
rect 1722 6500 1778 6556
rect 1778 6500 1782 6556
rect 1718 6496 1782 6500
rect 1798 6556 1862 6560
rect 1798 6500 1802 6556
rect 1802 6500 1858 6556
rect 1858 6500 1862 6556
rect 1798 6496 1862 6500
rect 4658 6556 4722 6560
rect 4658 6500 4662 6556
rect 4662 6500 4718 6556
rect 4718 6500 4722 6556
rect 4658 6496 4722 6500
rect 4738 6556 4802 6560
rect 4738 6500 4742 6556
rect 4742 6500 4798 6556
rect 4798 6500 4802 6556
rect 4738 6496 4802 6500
rect 4818 6556 4882 6560
rect 4818 6500 4822 6556
rect 4822 6500 4878 6556
rect 4878 6500 4882 6556
rect 4818 6496 4882 6500
rect 4898 6556 4962 6560
rect 4898 6500 4902 6556
rect 4902 6500 4958 6556
rect 4958 6500 4962 6556
rect 4898 6496 4962 6500
rect 7758 6556 7822 6560
rect 7758 6500 7762 6556
rect 7762 6500 7818 6556
rect 7818 6500 7822 6556
rect 7758 6496 7822 6500
rect 7838 6556 7902 6560
rect 7838 6500 7842 6556
rect 7842 6500 7898 6556
rect 7898 6500 7902 6556
rect 7838 6496 7902 6500
rect 7918 6556 7982 6560
rect 7918 6500 7922 6556
rect 7922 6500 7978 6556
rect 7978 6500 7982 6556
rect 7918 6496 7982 6500
rect 7998 6556 8062 6560
rect 7998 6500 8002 6556
rect 8002 6500 8058 6556
rect 8058 6500 8062 6556
rect 7998 6496 8062 6500
rect 10858 6556 10922 6560
rect 10858 6500 10862 6556
rect 10862 6500 10918 6556
rect 10918 6500 10922 6556
rect 10858 6496 10922 6500
rect 10938 6556 11002 6560
rect 10938 6500 10942 6556
rect 10942 6500 10998 6556
rect 10998 6500 11002 6556
rect 10938 6496 11002 6500
rect 11018 6556 11082 6560
rect 11018 6500 11022 6556
rect 11022 6500 11078 6556
rect 11078 6500 11082 6556
rect 11018 6496 11082 6500
rect 11098 6556 11162 6560
rect 11098 6500 11102 6556
rect 11102 6500 11158 6556
rect 11158 6500 11162 6556
rect 11098 6496 11162 6500
rect 13958 6556 14022 6560
rect 13958 6500 13962 6556
rect 13962 6500 14018 6556
rect 14018 6500 14022 6556
rect 13958 6496 14022 6500
rect 14038 6556 14102 6560
rect 14038 6500 14042 6556
rect 14042 6500 14098 6556
rect 14098 6500 14102 6556
rect 14038 6496 14102 6500
rect 14118 6556 14182 6560
rect 14118 6500 14122 6556
rect 14122 6500 14178 6556
rect 14178 6500 14182 6556
rect 14118 6496 14182 6500
rect 14198 6556 14262 6560
rect 14198 6500 14202 6556
rect 14202 6500 14258 6556
rect 14258 6500 14262 6556
rect 14198 6496 14262 6500
rect 17058 6556 17122 6560
rect 17058 6500 17062 6556
rect 17062 6500 17118 6556
rect 17118 6500 17122 6556
rect 17058 6496 17122 6500
rect 17138 6556 17202 6560
rect 17138 6500 17142 6556
rect 17142 6500 17198 6556
rect 17198 6500 17202 6556
rect 17138 6496 17202 6500
rect 17218 6556 17282 6560
rect 17218 6500 17222 6556
rect 17222 6500 17278 6556
rect 17278 6500 17282 6556
rect 17218 6496 17282 6500
rect 17298 6556 17362 6560
rect 17298 6500 17302 6556
rect 17302 6500 17358 6556
rect 17358 6500 17362 6556
rect 17298 6496 17362 6500
rect 3108 6012 3172 6016
rect 3108 5956 3112 6012
rect 3112 5956 3168 6012
rect 3168 5956 3172 6012
rect 3108 5952 3172 5956
rect 3188 6012 3252 6016
rect 3188 5956 3192 6012
rect 3192 5956 3248 6012
rect 3248 5956 3252 6012
rect 3188 5952 3252 5956
rect 3268 6012 3332 6016
rect 3268 5956 3272 6012
rect 3272 5956 3328 6012
rect 3328 5956 3332 6012
rect 3268 5952 3332 5956
rect 3348 6012 3412 6016
rect 3348 5956 3352 6012
rect 3352 5956 3408 6012
rect 3408 5956 3412 6012
rect 3348 5952 3412 5956
rect 6208 6012 6272 6016
rect 6208 5956 6212 6012
rect 6212 5956 6268 6012
rect 6268 5956 6272 6012
rect 6208 5952 6272 5956
rect 6288 6012 6352 6016
rect 6288 5956 6292 6012
rect 6292 5956 6348 6012
rect 6348 5956 6352 6012
rect 6288 5952 6352 5956
rect 6368 6012 6432 6016
rect 6368 5956 6372 6012
rect 6372 5956 6428 6012
rect 6428 5956 6432 6012
rect 6368 5952 6432 5956
rect 6448 6012 6512 6016
rect 6448 5956 6452 6012
rect 6452 5956 6508 6012
rect 6508 5956 6512 6012
rect 6448 5952 6512 5956
rect 9308 6012 9372 6016
rect 9308 5956 9312 6012
rect 9312 5956 9368 6012
rect 9368 5956 9372 6012
rect 9308 5952 9372 5956
rect 9388 6012 9452 6016
rect 9388 5956 9392 6012
rect 9392 5956 9448 6012
rect 9448 5956 9452 6012
rect 9388 5952 9452 5956
rect 9468 6012 9532 6016
rect 9468 5956 9472 6012
rect 9472 5956 9528 6012
rect 9528 5956 9532 6012
rect 9468 5952 9532 5956
rect 9548 6012 9612 6016
rect 9548 5956 9552 6012
rect 9552 5956 9608 6012
rect 9608 5956 9612 6012
rect 9548 5952 9612 5956
rect 12408 6012 12472 6016
rect 12408 5956 12412 6012
rect 12412 5956 12468 6012
rect 12468 5956 12472 6012
rect 12408 5952 12472 5956
rect 12488 6012 12552 6016
rect 12488 5956 12492 6012
rect 12492 5956 12548 6012
rect 12548 5956 12552 6012
rect 12488 5952 12552 5956
rect 12568 6012 12632 6016
rect 12568 5956 12572 6012
rect 12572 5956 12628 6012
rect 12628 5956 12632 6012
rect 12568 5952 12632 5956
rect 12648 6012 12712 6016
rect 12648 5956 12652 6012
rect 12652 5956 12708 6012
rect 12708 5956 12712 6012
rect 12648 5952 12712 5956
rect 15508 6012 15572 6016
rect 15508 5956 15512 6012
rect 15512 5956 15568 6012
rect 15568 5956 15572 6012
rect 15508 5952 15572 5956
rect 15588 6012 15652 6016
rect 15588 5956 15592 6012
rect 15592 5956 15648 6012
rect 15648 5956 15652 6012
rect 15588 5952 15652 5956
rect 15668 6012 15732 6016
rect 15668 5956 15672 6012
rect 15672 5956 15728 6012
rect 15728 5956 15732 6012
rect 15668 5952 15732 5956
rect 15748 6012 15812 6016
rect 15748 5956 15752 6012
rect 15752 5956 15808 6012
rect 15808 5956 15812 6012
rect 15748 5952 15812 5956
rect 18608 6012 18672 6016
rect 18608 5956 18612 6012
rect 18612 5956 18668 6012
rect 18668 5956 18672 6012
rect 18608 5952 18672 5956
rect 18688 6012 18752 6016
rect 18688 5956 18692 6012
rect 18692 5956 18748 6012
rect 18748 5956 18752 6012
rect 18688 5952 18752 5956
rect 18768 6012 18832 6016
rect 18768 5956 18772 6012
rect 18772 5956 18828 6012
rect 18828 5956 18832 6012
rect 18768 5952 18832 5956
rect 18848 6012 18912 6016
rect 18848 5956 18852 6012
rect 18852 5956 18908 6012
rect 18908 5956 18912 6012
rect 18848 5952 18912 5956
rect 1558 5468 1622 5472
rect 1558 5412 1562 5468
rect 1562 5412 1618 5468
rect 1618 5412 1622 5468
rect 1558 5408 1622 5412
rect 1638 5468 1702 5472
rect 1638 5412 1642 5468
rect 1642 5412 1698 5468
rect 1698 5412 1702 5468
rect 1638 5408 1702 5412
rect 1718 5468 1782 5472
rect 1718 5412 1722 5468
rect 1722 5412 1778 5468
rect 1778 5412 1782 5468
rect 1718 5408 1782 5412
rect 1798 5468 1862 5472
rect 1798 5412 1802 5468
rect 1802 5412 1858 5468
rect 1858 5412 1862 5468
rect 1798 5408 1862 5412
rect 4658 5468 4722 5472
rect 4658 5412 4662 5468
rect 4662 5412 4718 5468
rect 4718 5412 4722 5468
rect 4658 5408 4722 5412
rect 4738 5468 4802 5472
rect 4738 5412 4742 5468
rect 4742 5412 4798 5468
rect 4798 5412 4802 5468
rect 4738 5408 4802 5412
rect 4818 5468 4882 5472
rect 4818 5412 4822 5468
rect 4822 5412 4878 5468
rect 4878 5412 4882 5468
rect 4818 5408 4882 5412
rect 4898 5468 4962 5472
rect 4898 5412 4902 5468
rect 4902 5412 4958 5468
rect 4958 5412 4962 5468
rect 4898 5408 4962 5412
rect 7758 5468 7822 5472
rect 7758 5412 7762 5468
rect 7762 5412 7818 5468
rect 7818 5412 7822 5468
rect 7758 5408 7822 5412
rect 7838 5468 7902 5472
rect 7838 5412 7842 5468
rect 7842 5412 7898 5468
rect 7898 5412 7902 5468
rect 7838 5408 7902 5412
rect 7918 5468 7982 5472
rect 7918 5412 7922 5468
rect 7922 5412 7978 5468
rect 7978 5412 7982 5468
rect 7918 5408 7982 5412
rect 7998 5468 8062 5472
rect 7998 5412 8002 5468
rect 8002 5412 8058 5468
rect 8058 5412 8062 5468
rect 7998 5408 8062 5412
rect 10858 5468 10922 5472
rect 10858 5412 10862 5468
rect 10862 5412 10918 5468
rect 10918 5412 10922 5468
rect 10858 5408 10922 5412
rect 10938 5468 11002 5472
rect 10938 5412 10942 5468
rect 10942 5412 10998 5468
rect 10998 5412 11002 5468
rect 10938 5408 11002 5412
rect 11018 5468 11082 5472
rect 11018 5412 11022 5468
rect 11022 5412 11078 5468
rect 11078 5412 11082 5468
rect 11018 5408 11082 5412
rect 11098 5468 11162 5472
rect 11098 5412 11102 5468
rect 11102 5412 11158 5468
rect 11158 5412 11162 5468
rect 11098 5408 11162 5412
rect 13958 5468 14022 5472
rect 13958 5412 13962 5468
rect 13962 5412 14018 5468
rect 14018 5412 14022 5468
rect 13958 5408 14022 5412
rect 14038 5468 14102 5472
rect 14038 5412 14042 5468
rect 14042 5412 14098 5468
rect 14098 5412 14102 5468
rect 14038 5408 14102 5412
rect 14118 5468 14182 5472
rect 14118 5412 14122 5468
rect 14122 5412 14178 5468
rect 14178 5412 14182 5468
rect 14118 5408 14182 5412
rect 14198 5468 14262 5472
rect 14198 5412 14202 5468
rect 14202 5412 14258 5468
rect 14258 5412 14262 5468
rect 14198 5408 14262 5412
rect 17058 5468 17122 5472
rect 17058 5412 17062 5468
rect 17062 5412 17118 5468
rect 17118 5412 17122 5468
rect 17058 5408 17122 5412
rect 17138 5468 17202 5472
rect 17138 5412 17142 5468
rect 17142 5412 17198 5468
rect 17198 5412 17202 5468
rect 17138 5408 17202 5412
rect 17218 5468 17282 5472
rect 17218 5412 17222 5468
rect 17222 5412 17278 5468
rect 17278 5412 17282 5468
rect 17218 5408 17282 5412
rect 17298 5468 17362 5472
rect 17298 5412 17302 5468
rect 17302 5412 17358 5468
rect 17358 5412 17362 5468
rect 17298 5408 17362 5412
rect 3108 4924 3172 4928
rect 3108 4868 3112 4924
rect 3112 4868 3168 4924
rect 3168 4868 3172 4924
rect 3108 4864 3172 4868
rect 3188 4924 3252 4928
rect 3188 4868 3192 4924
rect 3192 4868 3248 4924
rect 3248 4868 3252 4924
rect 3188 4864 3252 4868
rect 3268 4924 3332 4928
rect 3268 4868 3272 4924
rect 3272 4868 3328 4924
rect 3328 4868 3332 4924
rect 3268 4864 3332 4868
rect 3348 4924 3412 4928
rect 3348 4868 3352 4924
rect 3352 4868 3408 4924
rect 3408 4868 3412 4924
rect 3348 4864 3412 4868
rect 6208 4924 6272 4928
rect 6208 4868 6212 4924
rect 6212 4868 6268 4924
rect 6268 4868 6272 4924
rect 6208 4864 6272 4868
rect 6288 4924 6352 4928
rect 6288 4868 6292 4924
rect 6292 4868 6348 4924
rect 6348 4868 6352 4924
rect 6288 4864 6352 4868
rect 6368 4924 6432 4928
rect 6368 4868 6372 4924
rect 6372 4868 6428 4924
rect 6428 4868 6432 4924
rect 6368 4864 6432 4868
rect 6448 4924 6512 4928
rect 6448 4868 6452 4924
rect 6452 4868 6508 4924
rect 6508 4868 6512 4924
rect 6448 4864 6512 4868
rect 9308 4924 9372 4928
rect 9308 4868 9312 4924
rect 9312 4868 9368 4924
rect 9368 4868 9372 4924
rect 9308 4864 9372 4868
rect 9388 4924 9452 4928
rect 9388 4868 9392 4924
rect 9392 4868 9448 4924
rect 9448 4868 9452 4924
rect 9388 4864 9452 4868
rect 9468 4924 9532 4928
rect 9468 4868 9472 4924
rect 9472 4868 9528 4924
rect 9528 4868 9532 4924
rect 9468 4864 9532 4868
rect 9548 4924 9612 4928
rect 9548 4868 9552 4924
rect 9552 4868 9608 4924
rect 9608 4868 9612 4924
rect 9548 4864 9612 4868
rect 12408 4924 12472 4928
rect 12408 4868 12412 4924
rect 12412 4868 12468 4924
rect 12468 4868 12472 4924
rect 12408 4864 12472 4868
rect 12488 4924 12552 4928
rect 12488 4868 12492 4924
rect 12492 4868 12548 4924
rect 12548 4868 12552 4924
rect 12488 4864 12552 4868
rect 12568 4924 12632 4928
rect 12568 4868 12572 4924
rect 12572 4868 12628 4924
rect 12628 4868 12632 4924
rect 12568 4864 12632 4868
rect 12648 4924 12712 4928
rect 12648 4868 12652 4924
rect 12652 4868 12708 4924
rect 12708 4868 12712 4924
rect 12648 4864 12712 4868
rect 15508 4924 15572 4928
rect 15508 4868 15512 4924
rect 15512 4868 15568 4924
rect 15568 4868 15572 4924
rect 15508 4864 15572 4868
rect 15588 4924 15652 4928
rect 15588 4868 15592 4924
rect 15592 4868 15648 4924
rect 15648 4868 15652 4924
rect 15588 4864 15652 4868
rect 15668 4924 15732 4928
rect 15668 4868 15672 4924
rect 15672 4868 15728 4924
rect 15728 4868 15732 4924
rect 15668 4864 15732 4868
rect 15748 4924 15812 4928
rect 15748 4868 15752 4924
rect 15752 4868 15808 4924
rect 15808 4868 15812 4924
rect 15748 4864 15812 4868
rect 18608 4924 18672 4928
rect 18608 4868 18612 4924
rect 18612 4868 18668 4924
rect 18668 4868 18672 4924
rect 18608 4864 18672 4868
rect 18688 4924 18752 4928
rect 18688 4868 18692 4924
rect 18692 4868 18748 4924
rect 18748 4868 18752 4924
rect 18688 4864 18752 4868
rect 18768 4924 18832 4928
rect 18768 4868 18772 4924
rect 18772 4868 18828 4924
rect 18828 4868 18832 4924
rect 18768 4864 18832 4868
rect 18848 4924 18912 4928
rect 18848 4868 18852 4924
rect 18852 4868 18908 4924
rect 18908 4868 18912 4924
rect 18848 4864 18912 4868
rect 1558 4380 1622 4384
rect 1558 4324 1562 4380
rect 1562 4324 1618 4380
rect 1618 4324 1622 4380
rect 1558 4320 1622 4324
rect 1638 4380 1702 4384
rect 1638 4324 1642 4380
rect 1642 4324 1698 4380
rect 1698 4324 1702 4380
rect 1638 4320 1702 4324
rect 1718 4380 1782 4384
rect 1718 4324 1722 4380
rect 1722 4324 1778 4380
rect 1778 4324 1782 4380
rect 1718 4320 1782 4324
rect 1798 4380 1862 4384
rect 1798 4324 1802 4380
rect 1802 4324 1858 4380
rect 1858 4324 1862 4380
rect 1798 4320 1862 4324
rect 4658 4380 4722 4384
rect 4658 4324 4662 4380
rect 4662 4324 4718 4380
rect 4718 4324 4722 4380
rect 4658 4320 4722 4324
rect 4738 4380 4802 4384
rect 4738 4324 4742 4380
rect 4742 4324 4798 4380
rect 4798 4324 4802 4380
rect 4738 4320 4802 4324
rect 4818 4380 4882 4384
rect 4818 4324 4822 4380
rect 4822 4324 4878 4380
rect 4878 4324 4882 4380
rect 4818 4320 4882 4324
rect 4898 4380 4962 4384
rect 4898 4324 4902 4380
rect 4902 4324 4958 4380
rect 4958 4324 4962 4380
rect 4898 4320 4962 4324
rect 7758 4380 7822 4384
rect 7758 4324 7762 4380
rect 7762 4324 7818 4380
rect 7818 4324 7822 4380
rect 7758 4320 7822 4324
rect 7838 4380 7902 4384
rect 7838 4324 7842 4380
rect 7842 4324 7898 4380
rect 7898 4324 7902 4380
rect 7838 4320 7902 4324
rect 7918 4380 7982 4384
rect 7918 4324 7922 4380
rect 7922 4324 7978 4380
rect 7978 4324 7982 4380
rect 7918 4320 7982 4324
rect 7998 4380 8062 4384
rect 7998 4324 8002 4380
rect 8002 4324 8058 4380
rect 8058 4324 8062 4380
rect 7998 4320 8062 4324
rect 10858 4380 10922 4384
rect 10858 4324 10862 4380
rect 10862 4324 10918 4380
rect 10918 4324 10922 4380
rect 10858 4320 10922 4324
rect 10938 4380 11002 4384
rect 10938 4324 10942 4380
rect 10942 4324 10998 4380
rect 10998 4324 11002 4380
rect 10938 4320 11002 4324
rect 11018 4380 11082 4384
rect 11018 4324 11022 4380
rect 11022 4324 11078 4380
rect 11078 4324 11082 4380
rect 11018 4320 11082 4324
rect 11098 4380 11162 4384
rect 11098 4324 11102 4380
rect 11102 4324 11158 4380
rect 11158 4324 11162 4380
rect 11098 4320 11162 4324
rect 13958 4380 14022 4384
rect 13958 4324 13962 4380
rect 13962 4324 14018 4380
rect 14018 4324 14022 4380
rect 13958 4320 14022 4324
rect 14038 4380 14102 4384
rect 14038 4324 14042 4380
rect 14042 4324 14098 4380
rect 14098 4324 14102 4380
rect 14038 4320 14102 4324
rect 14118 4380 14182 4384
rect 14118 4324 14122 4380
rect 14122 4324 14178 4380
rect 14178 4324 14182 4380
rect 14118 4320 14182 4324
rect 14198 4380 14262 4384
rect 14198 4324 14202 4380
rect 14202 4324 14258 4380
rect 14258 4324 14262 4380
rect 14198 4320 14262 4324
rect 17058 4380 17122 4384
rect 17058 4324 17062 4380
rect 17062 4324 17118 4380
rect 17118 4324 17122 4380
rect 17058 4320 17122 4324
rect 17138 4380 17202 4384
rect 17138 4324 17142 4380
rect 17142 4324 17198 4380
rect 17198 4324 17202 4380
rect 17138 4320 17202 4324
rect 17218 4380 17282 4384
rect 17218 4324 17222 4380
rect 17222 4324 17278 4380
rect 17278 4324 17282 4380
rect 17218 4320 17282 4324
rect 17298 4380 17362 4384
rect 17298 4324 17302 4380
rect 17302 4324 17358 4380
rect 17358 4324 17362 4380
rect 17298 4320 17362 4324
rect 3108 3836 3172 3840
rect 3108 3780 3112 3836
rect 3112 3780 3168 3836
rect 3168 3780 3172 3836
rect 3108 3776 3172 3780
rect 3188 3836 3252 3840
rect 3188 3780 3192 3836
rect 3192 3780 3248 3836
rect 3248 3780 3252 3836
rect 3188 3776 3252 3780
rect 3268 3836 3332 3840
rect 3268 3780 3272 3836
rect 3272 3780 3328 3836
rect 3328 3780 3332 3836
rect 3268 3776 3332 3780
rect 3348 3836 3412 3840
rect 3348 3780 3352 3836
rect 3352 3780 3408 3836
rect 3408 3780 3412 3836
rect 3348 3776 3412 3780
rect 6208 3836 6272 3840
rect 6208 3780 6212 3836
rect 6212 3780 6268 3836
rect 6268 3780 6272 3836
rect 6208 3776 6272 3780
rect 6288 3836 6352 3840
rect 6288 3780 6292 3836
rect 6292 3780 6348 3836
rect 6348 3780 6352 3836
rect 6288 3776 6352 3780
rect 6368 3836 6432 3840
rect 6368 3780 6372 3836
rect 6372 3780 6428 3836
rect 6428 3780 6432 3836
rect 6368 3776 6432 3780
rect 6448 3836 6512 3840
rect 6448 3780 6452 3836
rect 6452 3780 6508 3836
rect 6508 3780 6512 3836
rect 6448 3776 6512 3780
rect 9308 3836 9372 3840
rect 9308 3780 9312 3836
rect 9312 3780 9368 3836
rect 9368 3780 9372 3836
rect 9308 3776 9372 3780
rect 9388 3836 9452 3840
rect 9388 3780 9392 3836
rect 9392 3780 9448 3836
rect 9448 3780 9452 3836
rect 9388 3776 9452 3780
rect 9468 3836 9532 3840
rect 9468 3780 9472 3836
rect 9472 3780 9528 3836
rect 9528 3780 9532 3836
rect 9468 3776 9532 3780
rect 9548 3836 9612 3840
rect 9548 3780 9552 3836
rect 9552 3780 9608 3836
rect 9608 3780 9612 3836
rect 9548 3776 9612 3780
rect 12408 3836 12472 3840
rect 12408 3780 12412 3836
rect 12412 3780 12468 3836
rect 12468 3780 12472 3836
rect 12408 3776 12472 3780
rect 12488 3836 12552 3840
rect 12488 3780 12492 3836
rect 12492 3780 12548 3836
rect 12548 3780 12552 3836
rect 12488 3776 12552 3780
rect 12568 3836 12632 3840
rect 12568 3780 12572 3836
rect 12572 3780 12628 3836
rect 12628 3780 12632 3836
rect 12568 3776 12632 3780
rect 12648 3836 12712 3840
rect 12648 3780 12652 3836
rect 12652 3780 12708 3836
rect 12708 3780 12712 3836
rect 12648 3776 12712 3780
rect 15508 3836 15572 3840
rect 15508 3780 15512 3836
rect 15512 3780 15568 3836
rect 15568 3780 15572 3836
rect 15508 3776 15572 3780
rect 15588 3836 15652 3840
rect 15588 3780 15592 3836
rect 15592 3780 15648 3836
rect 15648 3780 15652 3836
rect 15588 3776 15652 3780
rect 15668 3836 15732 3840
rect 15668 3780 15672 3836
rect 15672 3780 15728 3836
rect 15728 3780 15732 3836
rect 15668 3776 15732 3780
rect 15748 3836 15812 3840
rect 15748 3780 15752 3836
rect 15752 3780 15808 3836
rect 15808 3780 15812 3836
rect 15748 3776 15812 3780
rect 18608 3836 18672 3840
rect 18608 3780 18612 3836
rect 18612 3780 18668 3836
rect 18668 3780 18672 3836
rect 18608 3776 18672 3780
rect 18688 3836 18752 3840
rect 18688 3780 18692 3836
rect 18692 3780 18748 3836
rect 18748 3780 18752 3836
rect 18688 3776 18752 3780
rect 18768 3836 18832 3840
rect 18768 3780 18772 3836
rect 18772 3780 18828 3836
rect 18828 3780 18832 3836
rect 18768 3776 18832 3780
rect 18848 3836 18912 3840
rect 18848 3780 18852 3836
rect 18852 3780 18908 3836
rect 18908 3780 18912 3836
rect 18848 3776 18912 3780
rect 1558 3292 1622 3296
rect 1558 3236 1562 3292
rect 1562 3236 1618 3292
rect 1618 3236 1622 3292
rect 1558 3232 1622 3236
rect 1638 3292 1702 3296
rect 1638 3236 1642 3292
rect 1642 3236 1698 3292
rect 1698 3236 1702 3292
rect 1638 3232 1702 3236
rect 1718 3292 1782 3296
rect 1718 3236 1722 3292
rect 1722 3236 1778 3292
rect 1778 3236 1782 3292
rect 1718 3232 1782 3236
rect 1798 3292 1862 3296
rect 1798 3236 1802 3292
rect 1802 3236 1858 3292
rect 1858 3236 1862 3292
rect 1798 3232 1862 3236
rect 4658 3292 4722 3296
rect 4658 3236 4662 3292
rect 4662 3236 4718 3292
rect 4718 3236 4722 3292
rect 4658 3232 4722 3236
rect 4738 3292 4802 3296
rect 4738 3236 4742 3292
rect 4742 3236 4798 3292
rect 4798 3236 4802 3292
rect 4738 3232 4802 3236
rect 4818 3292 4882 3296
rect 4818 3236 4822 3292
rect 4822 3236 4878 3292
rect 4878 3236 4882 3292
rect 4818 3232 4882 3236
rect 4898 3292 4962 3296
rect 4898 3236 4902 3292
rect 4902 3236 4958 3292
rect 4958 3236 4962 3292
rect 4898 3232 4962 3236
rect 7758 3292 7822 3296
rect 7758 3236 7762 3292
rect 7762 3236 7818 3292
rect 7818 3236 7822 3292
rect 7758 3232 7822 3236
rect 7838 3292 7902 3296
rect 7838 3236 7842 3292
rect 7842 3236 7898 3292
rect 7898 3236 7902 3292
rect 7838 3232 7902 3236
rect 7918 3292 7982 3296
rect 7918 3236 7922 3292
rect 7922 3236 7978 3292
rect 7978 3236 7982 3292
rect 7918 3232 7982 3236
rect 7998 3292 8062 3296
rect 7998 3236 8002 3292
rect 8002 3236 8058 3292
rect 8058 3236 8062 3292
rect 7998 3232 8062 3236
rect 10858 3292 10922 3296
rect 10858 3236 10862 3292
rect 10862 3236 10918 3292
rect 10918 3236 10922 3292
rect 10858 3232 10922 3236
rect 10938 3292 11002 3296
rect 10938 3236 10942 3292
rect 10942 3236 10998 3292
rect 10998 3236 11002 3292
rect 10938 3232 11002 3236
rect 11018 3292 11082 3296
rect 11018 3236 11022 3292
rect 11022 3236 11078 3292
rect 11078 3236 11082 3292
rect 11018 3232 11082 3236
rect 11098 3292 11162 3296
rect 11098 3236 11102 3292
rect 11102 3236 11158 3292
rect 11158 3236 11162 3292
rect 11098 3232 11162 3236
rect 13958 3292 14022 3296
rect 13958 3236 13962 3292
rect 13962 3236 14018 3292
rect 14018 3236 14022 3292
rect 13958 3232 14022 3236
rect 14038 3292 14102 3296
rect 14038 3236 14042 3292
rect 14042 3236 14098 3292
rect 14098 3236 14102 3292
rect 14038 3232 14102 3236
rect 14118 3292 14182 3296
rect 14118 3236 14122 3292
rect 14122 3236 14178 3292
rect 14178 3236 14182 3292
rect 14118 3232 14182 3236
rect 14198 3292 14262 3296
rect 14198 3236 14202 3292
rect 14202 3236 14258 3292
rect 14258 3236 14262 3292
rect 14198 3232 14262 3236
rect 17058 3292 17122 3296
rect 17058 3236 17062 3292
rect 17062 3236 17118 3292
rect 17118 3236 17122 3292
rect 17058 3232 17122 3236
rect 17138 3292 17202 3296
rect 17138 3236 17142 3292
rect 17142 3236 17198 3292
rect 17198 3236 17202 3292
rect 17138 3232 17202 3236
rect 17218 3292 17282 3296
rect 17218 3236 17222 3292
rect 17222 3236 17278 3292
rect 17278 3236 17282 3292
rect 17218 3232 17282 3236
rect 17298 3292 17362 3296
rect 17298 3236 17302 3292
rect 17302 3236 17358 3292
rect 17358 3236 17362 3292
rect 17298 3232 17362 3236
rect 3108 2748 3172 2752
rect 3108 2692 3112 2748
rect 3112 2692 3168 2748
rect 3168 2692 3172 2748
rect 3108 2688 3172 2692
rect 3188 2748 3252 2752
rect 3188 2692 3192 2748
rect 3192 2692 3248 2748
rect 3248 2692 3252 2748
rect 3188 2688 3252 2692
rect 3268 2748 3332 2752
rect 3268 2692 3272 2748
rect 3272 2692 3328 2748
rect 3328 2692 3332 2748
rect 3268 2688 3332 2692
rect 3348 2748 3412 2752
rect 3348 2692 3352 2748
rect 3352 2692 3408 2748
rect 3408 2692 3412 2748
rect 3348 2688 3412 2692
rect 6208 2748 6272 2752
rect 6208 2692 6212 2748
rect 6212 2692 6268 2748
rect 6268 2692 6272 2748
rect 6208 2688 6272 2692
rect 6288 2748 6352 2752
rect 6288 2692 6292 2748
rect 6292 2692 6348 2748
rect 6348 2692 6352 2748
rect 6288 2688 6352 2692
rect 6368 2748 6432 2752
rect 6368 2692 6372 2748
rect 6372 2692 6428 2748
rect 6428 2692 6432 2748
rect 6368 2688 6432 2692
rect 6448 2748 6512 2752
rect 6448 2692 6452 2748
rect 6452 2692 6508 2748
rect 6508 2692 6512 2748
rect 6448 2688 6512 2692
rect 9308 2748 9372 2752
rect 9308 2692 9312 2748
rect 9312 2692 9368 2748
rect 9368 2692 9372 2748
rect 9308 2688 9372 2692
rect 9388 2748 9452 2752
rect 9388 2692 9392 2748
rect 9392 2692 9448 2748
rect 9448 2692 9452 2748
rect 9388 2688 9452 2692
rect 9468 2748 9532 2752
rect 9468 2692 9472 2748
rect 9472 2692 9528 2748
rect 9528 2692 9532 2748
rect 9468 2688 9532 2692
rect 9548 2748 9612 2752
rect 9548 2692 9552 2748
rect 9552 2692 9608 2748
rect 9608 2692 9612 2748
rect 9548 2688 9612 2692
rect 12408 2748 12472 2752
rect 12408 2692 12412 2748
rect 12412 2692 12468 2748
rect 12468 2692 12472 2748
rect 12408 2688 12472 2692
rect 12488 2748 12552 2752
rect 12488 2692 12492 2748
rect 12492 2692 12548 2748
rect 12548 2692 12552 2748
rect 12488 2688 12552 2692
rect 12568 2748 12632 2752
rect 12568 2692 12572 2748
rect 12572 2692 12628 2748
rect 12628 2692 12632 2748
rect 12568 2688 12632 2692
rect 12648 2748 12712 2752
rect 12648 2692 12652 2748
rect 12652 2692 12708 2748
rect 12708 2692 12712 2748
rect 12648 2688 12712 2692
rect 15508 2748 15572 2752
rect 15508 2692 15512 2748
rect 15512 2692 15568 2748
rect 15568 2692 15572 2748
rect 15508 2688 15572 2692
rect 15588 2748 15652 2752
rect 15588 2692 15592 2748
rect 15592 2692 15648 2748
rect 15648 2692 15652 2748
rect 15588 2688 15652 2692
rect 15668 2748 15732 2752
rect 15668 2692 15672 2748
rect 15672 2692 15728 2748
rect 15728 2692 15732 2748
rect 15668 2688 15732 2692
rect 15748 2748 15812 2752
rect 15748 2692 15752 2748
rect 15752 2692 15808 2748
rect 15808 2692 15812 2748
rect 15748 2688 15812 2692
rect 18608 2748 18672 2752
rect 18608 2692 18612 2748
rect 18612 2692 18668 2748
rect 18668 2692 18672 2748
rect 18608 2688 18672 2692
rect 18688 2748 18752 2752
rect 18688 2692 18692 2748
rect 18692 2692 18748 2748
rect 18748 2692 18752 2748
rect 18688 2688 18752 2692
rect 18768 2748 18832 2752
rect 18768 2692 18772 2748
rect 18772 2692 18828 2748
rect 18828 2692 18832 2748
rect 18768 2688 18832 2692
rect 18848 2748 18912 2752
rect 18848 2692 18852 2748
rect 18852 2692 18908 2748
rect 18908 2692 18912 2748
rect 18848 2688 18912 2692
rect 1558 2204 1622 2208
rect 1558 2148 1562 2204
rect 1562 2148 1618 2204
rect 1618 2148 1622 2204
rect 1558 2144 1622 2148
rect 1638 2204 1702 2208
rect 1638 2148 1642 2204
rect 1642 2148 1698 2204
rect 1698 2148 1702 2204
rect 1638 2144 1702 2148
rect 1718 2204 1782 2208
rect 1718 2148 1722 2204
rect 1722 2148 1778 2204
rect 1778 2148 1782 2204
rect 1718 2144 1782 2148
rect 1798 2204 1862 2208
rect 1798 2148 1802 2204
rect 1802 2148 1858 2204
rect 1858 2148 1862 2204
rect 1798 2144 1862 2148
rect 4658 2204 4722 2208
rect 4658 2148 4662 2204
rect 4662 2148 4718 2204
rect 4718 2148 4722 2204
rect 4658 2144 4722 2148
rect 4738 2204 4802 2208
rect 4738 2148 4742 2204
rect 4742 2148 4798 2204
rect 4798 2148 4802 2204
rect 4738 2144 4802 2148
rect 4818 2204 4882 2208
rect 4818 2148 4822 2204
rect 4822 2148 4878 2204
rect 4878 2148 4882 2204
rect 4818 2144 4882 2148
rect 4898 2204 4962 2208
rect 4898 2148 4902 2204
rect 4902 2148 4958 2204
rect 4958 2148 4962 2204
rect 4898 2144 4962 2148
rect 7758 2204 7822 2208
rect 7758 2148 7762 2204
rect 7762 2148 7818 2204
rect 7818 2148 7822 2204
rect 7758 2144 7822 2148
rect 7838 2204 7902 2208
rect 7838 2148 7842 2204
rect 7842 2148 7898 2204
rect 7898 2148 7902 2204
rect 7838 2144 7902 2148
rect 7918 2204 7982 2208
rect 7918 2148 7922 2204
rect 7922 2148 7978 2204
rect 7978 2148 7982 2204
rect 7918 2144 7982 2148
rect 7998 2204 8062 2208
rect 7998 2148 8002 2204
rect 8002 2148 8058 2204
rect 8058 2148 8062 2204
rect 7998 2144 8062 2148
rect 10858 2204 10922 2208
rect 10858 2148 10862 2204
rect 10862 2148 10918 2204
rect 10918 2148 10922 2204
rect 10858 2144 10922 2148
rect 10938 2204 11002 2208
rect 10938 2148 10942 2204
rect 10942 2148 10998 2204
rect 10998 2148 11002 2204
rect 10938 2144 11002 2148
rect 11018 2204 11082 2208
rect 11018 2148 11022 2204
rect 11022 2148 11078 2204
rect 11078 2148 11082 2204
rect 11018 2144 11082 2148
rect 11098 2204 11162 2208
rect 11098 2148 11102 2204
rect 11102 2148 11158 2204
rect 11158 2148 11162 2204
rect 11098 2144 11162 2148
rect 13958 2204 14022 2208
rect 13958 2148 13962 2204
rect 13962 2148 14018 2204
rect 14018 2148 14022 2204
rect 13958 2144 14022 2148
rect 14038 2204 14102 2208
rect 14038 2148 14042 2204
rect 14042 2148 14098 2204
rect 14098 2148 14102 2204
rect 14038 2144 14102 2148
rect 14118 2204 14182 2208
rect 14118 2148 14122 2204
rect 14122 2148 14178 2204
rect 14178 2148 14182 2204
rect 14118 2144 14182 2148
rect 14198 2204 14262 2208
rect 14198 2148 14202 2204
rect 14202 2148 14258 2204
rect 14258 2148 14262 2204
rect 14198 2144 14262 2148
rect 17058 2204 17122 2208
rect 17058 2148 17062 2204
rect 17062 2148 17118 2204
rect 17118 2148 17122 2204
rect 17058 2144 17122 2148
rect 17138 2204 17202 2208
rect 17138 2148 17142 2204
rect 17142 2148 17198 2204
rect 17198 2148 17202 2204
rect 17138 2144 17202 2148
rect 17218 2204 17282 2208
rect 17218 2148 17222 2204
rect 17222 2148 17278 2204
rect 17278 2148 17282 2204
rect 17218 2144 17282 2148
rect 17298 2204 17362 2208
rect 17298 2148 17302 2204
rect 17302 2148 17358 2204
rect 17358 2148 17362 2204
rect 17298 2144 17362 2148
rect 3108 1660 3172 1664
rect 3108 1604 3112 1660
rect 3112 1604 3168 1660
rect 3168 1604 3172 1660
rect 3108 1600 3172 1604
rect 3188 1660 3252 1664
rect 3188 1604 3192 1660
rect 3192 1604 3248 1660
rect 3248 1604 3252 1660
rect 3188 1600 3252 1604
rect 3268 1660 3332 1664
rect 3268 1604 3272 1660
rect 3272 1604 3328 1660
rect 3328 1604 3332 1660
rect 3268 1600 3332 1604
rect 3348 1660 3412 1664
rect 3348 1604 3352 1660
rect 3352 1604 3408 1660
rect 3408 1604 3412 1660
rect 3348 1600 3412 1604
rect 6208 1660 6272 1664
rect 6208 1604 6212 1660
rect 6212 1604 6268 1660
rect 6268 1604 6272 1660
rect 6208 1600 6272 1604
rect 6288 1660 6352 1664
rect 6288 1604 6292 1660
rect 6292 1604 6348 1660
rect 6348 1604 6352 1660
rect 6288 1600 6352 1604
rect 6368 1660 6432 1664
rect 6368 1604 6372 1660
rect 6372 1604 6428 1660
rect 6428 1604 6432 1660
rect 6368 1600 6432 1604
rect 6448 1660 6512 1664
rect 6448 1604 6452 1660
rect 6452 1604 6508 1660
rect 6508 1604 6512 1660
rect 6448 1600 6512 1604
rect 9308 1660 9372 1664
rect 9308 1604 9312 1660
rect 9312 1604 9368 1660
rect 9368 1604 9372 1660
rect 9308 1600 9372 1604
rect 9388 1660 9452 1664
rect 9388 1604 9392 1660
rect 9392 1604 9448 1660
rect 9448 1604 9452 1660
rect 9388 1600 9452 1604
rect 9468 1660 9532 1664
rect 9468 1604 9472 1660
rect 9472 1604 9528 1660
rect 9528 1604 9532 1660
rect 9468 1600 9532 1604
rect 9548 1660 9612 1664
rect 9548 1604 9552 1660
rect 9552 1604 9608 1660
rect 9608 1604 9612 1660
rect 9548 1600 9612 1604
rect 12408 1660 12472 1664
rect 12408 1604 12412 1660
rect 12412 1604 12468 1660
rect 12468 1604 12472 1660
rect 12408 1600 12472 1604
rect 12488 1660 12552 1664
rect 12488 1604 12492 1660
rect 12492 1604 12548 1660
rect 12548 1604 12552 1660
rect 12488 1600 12552 1604
rect 12568 1660 12632 1664
rect 12568 1604 12572 1660
rect 12572 1604 12628 1660
rect 12628 1604 12632 1660
rect 12568 1600 12632 1604
rect 12648 1660 12712 1664
rect 12648 1604 12652 1660
rect 12652 1604 12708 1660
rect 12708 1604 12712 1660
rect 12648 1600 12712 1604
rect 15508 1660 15572 1664
rect 15508 1604 15512 1660
rect 15512 1604 15568 1660
rect 15568 1604 15572 1660
rect 15508 1600 15572 1604
rect 15588 1660 15652 1664
rect 15588 1604 15592 1660
rect 15592 1604 15648 1660
rect 15648 1604 15652 1660
rect 15588 1600 15652 1604
rect 15668 1660 15732 1664
rect 15668 1604 15672 1660
rect 15672 1604 15728 1660
rect 15728 1604 15732 1660
rect 15668 1600 15732 1604
rect 15748 1660 15812 1664
rect 15748 1604 15752 1660
rect 15752 1604 15808 1660
rect 15808 1604 15812 1660
rect 15748 1600 15812 1604
rect 18608 1660 18672 1664
rect 18608 1604 18612 1660
rect 18612 1604 18668 1660
rect 18668 1604 18672 1660
rect 18608 1600 18672 1604
rect 18688 1660 18752 1664
rect 18688 1604 18692 1660
rect 18692 1604 18748 1660
rect 18748 1604 18752 1660
rect 18688 1600 18752 1604
rect 18768 1660 18832 1664
rect 18768 1604 18772 1660
rect 18772 1604 18828 1660
rect 18828 1604 18832 1660
rect 18768 1600 18832 1604
rect 18848 1660 18912 1664
rect 18848 1604 18852 1660
rect 18852 1604 18908 1660
rect 18908 1604 18912 1660
rect 18848 1600 18912 1604
rect 1558 1116 1622 1120
rect 1558 1060 1562 1116
rect 1562 1060 1618 1116
rect 1618 1060 1622 1116
rect 1558 1056 1622 1060
rect 1638 1116 1702 1120
rect 1638 1060 1642 1116
rect 1642 1060 1698 1116
rect 1698 1060 1702 1116
rect 1638 1056 1702 1060
rect 1718 1116 1782 1120
rect 1718 1060 1722 1116
rect 1722 1060 1778 1116
rect 1778 1060 1782 1116
rect 1718 1056 1782 1060
rect 1798 1116 1862 1120
rect 1798 1060 1802 1116
rect 1802 1060 1858 1116
rect 1858 1060 1862 1116
rect 1798 1056 1862 1060
rect 4658 1116 4722 1120
rect 4658 1060 4662 1116
rect 4662 1060 4718 1116
rect 4718 1060 4722 1116
rect 4658 1056 4722 1060
rect 4738 1116 4802 1120
rect 4738 1060 4742 1116
rect 4742 1060 4798 1116
rect 4798 1060 4802 1116
rect 4738 1056 4802 1060
rect 4818 1116 4882 1120
rect 4818 1060 4822 1116
rect 4822 1060 4878 1116
rect 4878 1060 4882 1116
rect 4818 1056 4882 1060
rect 4898 1116 4962 1120
rect 4898 1060 4902 1116
rect 4902 1060 4958 1116
rect 4958 1060 4962 1116
rect 4898 1056 4962 1060
rect 7758 1116 7822 1120
rect 7758 1060 7762 1116
rect 7762 1060 7818 1116
rect 7818 1060 7822 1116
rect 7758 1056 7822 1060
rect 7838 1116 7902 1120
rect 7838 1060 7842 1116
rect 7842 1060 7898 1116
rect 7898 1060 7902 1116
rect 7838 1056 7902 1060
rect 7918 1116 7982 1120
rect 7918 1060 7922 1116
rect 7922 1060 7978 1116
rect 7978 1060 7982 1116
rect 7918 1056 7982 1060
rect 7998 1116 8062 1120
rect 7998 1060 8002 1116
rect 8002 1060 8058 1116
rect 8058 1060 8062 1116
rect 7998 1056 8062 1060
rect 10858 1116 10922 1120
rect 10858 1060 10862 1116
rect 10862 1060 10918 1116
rect 10918 1060 10922 1116
rect 10858 1056 10922 1060
rect 10938 1116 11002 1120
rect 10938 1060 10942 1116
rect 10942 1060 10998 1116
rect 10998 1060 11002 1116
rect 10938 1056 11002 1060
rect 11018 1116 11082 1120
rect 11018 1060 11022 1116
rect 11022 1060 11078 1116
rect 11078 1060 11082 1116
rect 11018 1056 11082 1060
rect 11098 1116 11162 1120
rect 11098 1060 11102 1116
rect 11102 1060 11158 1116
rect 11158 1060 11162 1116
rect 11098 1056 11162 1060
rect 13958 1116 14022 1120
rect 13958 1060 13962 1116
rect 13962 1060 14018 1116
rect 14018 1060 14022 1116
rect 13958 1056 14022 1060
rect 14038 1116 14102 1120
rect 14038 1060 14042 1116
rect 14042 1060 14098 1116
rect 14098 1060 14102 1116
rect 14038 1056 14102 1060
rect 14118 1116 14182 1120
rect 14118 1060 14122 1116
rect 14122 1060 14178 1116
rect 14178 1060 14182 1116
rect 14118 1056 14182 1060
rect 14198 1116 14262 1120
rect 14198 1060 14202 1116
rect 14202 1060 14258 1116
rect 14258 1060 14262 1116
rect 14198 1056 14262 1060
rect 17058 1116 17122 1120
rect 17058 1060 17062 1116
rect 17062 1060 17118 1116
rect 17118 1060 17122 1116
rect 17058 1056 17122 1060
rect 17138 1116 17202 1120
rect 17138 1060 17142 1116
rect 17142 1060 17198 1116
rect 17198 1060 17202 1116
rect 17138 1056 17202 1060
rect 17218 1116 17282 1120
rect 17218 1060 17222 1116
rect 17222 1060 17278 1116
rect 17278 1060 17282 1116
rect 17218 1056 17282 1060
rect 17298 1116 17362 1120
rect 17298 1060 17302 1116
rect 17302 1060 17358 1116
rect 17358 1060 17362 1116
rect 17298 1056 17362 1060
rect 3108 572 3172 576
rect 3108 516 3112 572
rect 3112 516 3168 572
rect 3168 516 3172 572
rect 3108 512 3172 516
rect 3188 572 3252 576
rect 3188 516 3192 572
rect 3192 516 3248 572
rect 3248 516 3252 572
rect 3188 512 3252 516
rect 3268 572 3332 576
rect 3268 516 3272 572
rect 3272 516 3328 572
rect 3328 516 3332 572
rect 3268 512 3332 516
rect 3348 572 3412 576
rect 3348 516 3352 572
rect 3352 516 3408 572
rect 3408 516 3412 572
rect 3348 512 3412 516
rect 6208 572 6272 576
rect 6208 516 6212 572
rect 6212 516 6268 572
rect 6268 516 6272 572
rect 6208 512 6272 516
rect 6288 572 6352 576
rect 6288 516 6292 572
rect 6292 516 6348 572
rect 6348 516 6352 572
rect 6288 512 6352 516
rect 6368 572 6432 576
rect 6368 516 6372 572
rect 6372 516 6428 572
rect 6428 516 6432 572
rect 6368 512 6432 516
rect 6448 572 6512 576
rect 6448 516 6452 572
rect 6452 516 6508 572
rect 6508 516 6512 572
rect 6448 512 6512 516
rect 9308 572 9372 576
rect 9308 516 9312 572
rect 9312 516 9368 572
rect 9368 516 9372 572
rect 9308 512 9372 516
rect 9388 572 9452 576
rect 9388 516 9392 572
rect 9392 516 9448 572
rect 9448 516 9452 572
rect 9388 512 9452 516
rect 9468 572 9532 576
rect 9468 516 9472 572
rect 9472 516 9528 572
rect 9528 516 9532 572
rect 9468 512 9532 516
rect 9548 572 9612 576
rect 9548 516 9552 572
rect 9552 516 9608 572
rect 9608 516 9612 572
rect 9548 512 9612 516
rect 12408 572 12472 576
rect 12408 516 12412 572
rect 12412 516 12468 572
rect 12468 516 12472 572
rect 12408 512 12472 516
rect 12488 572 12552 576
rect 12488 516 12492 572
rect 12492 516 12548 572
rect 12548 516 12552 572
rect 12488 512 12552 516
rect 12568 572 12632 576
rect 12568 516 12572 572
rect 12572 516 12628 572
rect 12628 516 12632 572
rect 12568 512 12632 516
rect 12648 572 12712 576
rect 12648 516 12652 572
rect 12652 516 12708 572
rect 12708 516 12712 572
rect 12648 512 12712 516
rect 15508 572 15572 576
rect 15508 516 15512 572
rect 15512 516 15568 572
rect 15568 516 15572 572
rect 15508 512 15572 516
rect 15588 572 15652 576
rect 15588 516 15592 572
rect 15592 516 15648 572
rect 15648 516 15652 572
rect 15588 512 15652 516
rect 15668 572 15732 576
rect 15668 516 15672 572
rect 15672 516 15728 572
rect 15728 516 15732 572
rect 15668 512 15732 516
rect 15748 572 15812 576
rect 15748 516 15752 572
rect 15752 516 15808 572
rect 15808 516 15812 572
rect 15748 512 15812 516
rect 18608 572 18672 576
rect 18608 516 18612 572
rect 18612 516 18668 572
rect 18668 516 18672 572
rect 18608 512 18672 516
rect 18688 572 18752 576
rect 18688 516 18692 572
rect 18692 516 18748 572
rect 18748 516 18752 572
rect 18688 512 18752 516
rect 18768 572 18832 576
rect 18768 516 18772 572
rect 18772 516 18828 572
rect 18828 516 18832 572
rect 18768 512 18832 516
rect 18848 572 18912 576
rect 18848 516 18852 572
rect 18852 516 18908 572
rect 18908 516 18912 572
rect 18848 512 18912 516
<< metal4 >>
rect 1550 18528 1870 18544
rect 1550 18464 1558 18528
rect 1622 18464 1638 18528
rect 1702 18464 1718 18528
rect 1782 18464 1798 18528
rect 1862 18464 1870 18528
rect 1550 17440 1870 18464
rect 1550 17376 1558 17440
rect 1622 17376 1638 17440
rect 1702 17376 1718 17440
rect 1782 17376 1798 17440
rect 1862 17376 1870 17440
rect 1550 16352 1870 17376
rect 1550 16288 1558 16352
rect 1622 16288 1638 16352
rect 1702 16288 1718 16352
rect 1782 16288 1798 16352
rect 1862 16288 1870 16352
rect 1550 15328 1870 16288
rect 1550 15264 1592 15328
rect 1828 15264 1870 15328
rect 1550 15200 1558 15264
rect 1862 15200 1870 15264
rect 1550 15092 1592 15200
rect 1828 15092 1870 15200
rect 1550 14176 1870 15092
rect 1550 14112 1558 14176
rect 1622 14112 1638 14176
rect 1702 14112 1718 14176
rect 1782 14112 1798 14176
rect 1862 14112 1870 14176
rect 1550 13088 1870 14112
rect 1550 13024 1558 13088
rect 1622 13024 1638 13088
rect 1702 13024 1718 13088
rect 1782 13024 1798 13088
rect 1862 13024 1870 13088
rect 1550 12000 1870 13024
rect 1550 11936 1558 12000
rect 1622 11948 1638 12000
rect 1702 11948 1718 12000
rect 1782 11948 1798 12000
rect 1862 11936 1870 12000
rect 1550 11712 1592 11936
rect 1828 11712 1870 11936
rect 1550 10912 1870 11712
rect 1550 10848 1558 10912
rect 1622 10848 1638 10912
rect 1702 10848 1718 10912
rect 1782 10848 1798 10912
rect 1862 10848 1870 10912
rect 1550 9824 1870 10848
rect 1550 9760 1558 9824
rect 1622 9760 1638 9824
rect 1702 9760 1718 9824
rect 1782 9760 1798 9824
rect 1862 9760 1870 9824
rect 1550 8736 1870 9760
rect 1550 8672 1558 8736
rect 1622 8672 1638 8736
rect 1702 8672 1718 8736
rect 1782 8672 1798 8736
rect 1862 8672 1870 8736
rect 1550 8568 1870 8672
rect 1550 8332 1592 8568
rect 1828 8332 1870 8568
rect 1550 7648 1870 8332
rect 1550 7584 1558 7648
rect 1622 7584 1638 7648
rect 1702 7584 1718 7648
rect 1782 7584 1798 7648
rect 1862 7584 1870 7648
rect 1550 6560 1870 7584
rect 1550 6496 1558 6560
rect 1622 6496 1638 6560
rect 1702 6496 1718 6560
rect 1782 6496 1798 6560
rect 1862 6496 1870 6560
rect 1550 5472 1870 6496
rect 1550 5408 1558 5472
rect 1622 5408 1638 5472
rect 1702 5408 1718 5472
rect 1782 5408 1798 5472
rect 1862 5408 1870 5472
rect 1550 5188 1870 5408
rect 1550 4952 1592 5188
rect 1828 4952 1870 5188
rect 1550 4384 1870 4952
rect 1550 4320 1558 4384
rect 1622 4320 1638 4384
rect 1702 4320 1718 4384
rect 1782 4320 1798 4384
rect 1862 4320 1870 4384
rect 1550 3296 1870 4320
rect 1550 3232 1558 3296
rect 1622 3232 1638 3296
rect 1702 3232 1718 3296
rect 1782 3232 1798 3296
rect 1862 3232 1870 3296
rect 1550 2208 1870 3232
rect 1550 2144 1558 2208
rect 1622 2144 1638 2208
rect 1702 2144 1718 2208
rect 1782 2144 1798 2208
rect 1862 2144 1870 2208
rect 1550 1808 1870 2144
rect 1550 1572 1592 1808
rect 1828 1572 1870 1808
rect 1550 1120 1870 1572
rect 1550 1056 1558 1120
rect 1622 1056 1638 1120
rect 1702 1056 1718 1120
rect 1782 1056 1798 1120
rect 1862 1056 1870 1120
rect 1550 496 1870 1056
rect 3100 17984 3420 18544
rect 3100 17920 3108 17984
rect 3172 17920 3188 17984
rect 3252 17920 3268 17984
rect 3332 17920 3348 17984
rect 3412 17920 3420 17984
rect 3100 17018 3420 17920
rect 3100 16896 3142 17018
rect 3378 16896 3420 17018
rect 3100 16832 3108 16896
rect 3412 16832 3420 16896
rect 3100 16782 3142 16832
rect 3378 16782 3420 16832
rect 3100 15808 3420 16782
rect 3100 15744 3108 15808
rect 3172 15744 3188 15808
rect 3252 15744 3268 15808
rect 3332 15744 3348 15808
rect 3412 15744 3420 15808
rect 3100 14720 3420 15744
rect 3100 14656 3108 14720
rect 3172 14656 3188 14720
rect 3252 14656 3268 14720
rect 3332 14656 3348 14720
rect 3412 14656 3420 14720
rect 3100 13638 3420 14656
rect 3100 13632 3142 13638
rect 3378 13632 3420 13638
rect 3100 13568 3108 13632
rect 3412 13568 3420 13632
rect 3100 13402 3142 13568
rect 3378 13402 3420 13568
rect 3100 12544 3420 13402
rect 3100 12480 3108 12544
rect 3172 12480 3188 12544
rect 3252 12480 3268 12544
rect 3332 12480 3348 12544
rect 3412 12480 3420 12544
rect 3100 11456 3420 12480
rect 3100 11392 3108 11456
rect 3172 11392 3188 11456
rect 3252 11392 3268 11456
rect 3332 11392 3348 11456
rect 3412 11392 3420 11456
rect 3100 10368 3420 11392
rect 3100 10304 3108 10368
rect 3172 10304 3188 10368
rect 3252 10304 3268 10368
rect 3332 10304 3348 10368
rect 3412 10304 3420 10368
rect 3100 10258 3420 10304
rect 3100 10022 3142 10258
rect 3378 10022 3420 10258
rect 3100 9280 3420 10022
rect 3100 9216 3108 9280
rect 3172 9216 3188 9280
rect 3252 9216 3268 9280
rect 3332 9216 3348 9280
rect 3412 9216 3420 9280
rect 3100 8192 3420 9216
rect 3100 8128 3108 8192
rect 3172 8128 3188 8192
rect 3252 8128 3268 8192
rect 3332 8128 3348 8192
rect 3412 8128 3420 8192
rect 3100 7104 3420 8128
rect 3100 7040 3108 7104
rect 3172 7040 3188 7104
rect 3252 7040 3268 7104
rect 3332 7040 3348 7104
rect 3412 7040 3420 7104
rect 3100 6878 3420 7040
rect 3100 6642 3142 6878
rect 3378 6642 3420 6878
rect 3100 6016 3420 6642
rect 3100 5952 3108 6016
rect 3172 5952 3188 6016
rect 3252 5952 3268 6016
rect 3332 5952 3348 6016
rect 3412 5952 3420 6016
rect 3100 4928 3420 5952
rect 3100 4864 3108 4928
rect 3172 4864 3188 4928
rect 3252 4864 3268 4928
rect 3332 4864 3348 4928
rect 3412 4864 3420 4928
rect 3100 3840 3420 4864
rect 3100 3776 3108 3840
rect 3172 3776 3188 3840
rect 3252 3776 3268 3840
rect 3332 3776 3348 3840
rect 3412 3776 3420 3840
rect 3100 3498 3420 3776
rect 3100 3262 3142 3498
rect 3378 3262 3420 3498
rect 3100 2752 3420 3262
rect 3100 2688 3108 2752
rect 3172 2688 3188 2752
rect 3252 2688 3268 2752
rect 3332 2688 3348 2752
rect 3412 2688 3420 2752
rect 3100 1664 3420 2688
rect 3100 1600 3108 1664
rect 3172 1600 3188 1664
rect 3252 1600 3268 1664
rect 3332 1600 3348 1664
rect 3412 1600 3420 1664
rect 3100 576 3420 1600
rect 3100 512 3108 576
rect 3172 512 3188 576
rect 3252 512 3268 576
rect 3332 512 3348 576
rect 3412 512 3420 576
rect 3100 496 3420 512
rect 4650 18528 4970 18544
rect 4650 18464 4658 18528
rect 4722 18464 4738 18528
rect 4802 18464 4818 18528
rect 4882 18464 4898 18528
rect 4962 18464 4970 18528
rect 4650 17440 4970 18464
rect 4650 17376 4658 17440
rect 4722 17376 4738 17440
rect 4802 17376 4818 17440
rect 4882 17376 4898 17440
rect 4962 17376 4970 17440
rect 4650 16352 4970 17376
rect 4650 16288 4658 16352
rect 4722 16288 4738 16352
rect 4802 16288 4818 16352
rect 4882 16288 4898 16352
rect 4962 16288 4970 16352
rect 4650 15328 4970 16288
rect 4650 15264 4692 15328
rect 4928 15264 4970 15328
rect 4650 15200 4658 15264
rect 4962 15200 4970 15264
rect 4650 15092 4692 15200
rect 4928 15092 4970 15200
rect 4650 14176 4970 15092
rect 4650 14112 4658 14176
rect 4722 14112 4738 14176
rect 4802 14112 4818 14176
rect 4882 14112 4898 14176
rect 4962 14112 4970 14176
rect 4650 13088 4970 14112
rect 4650 13024 4658 13088
rect 4722 13024 4738 13088
rect 4802 13024 4818 13088
rect 4882 13024 4898 13088
rect 4962 13024 4970 13088
rect 4650 12000 4970 13024
rect 4650 11936 4658 12000
rect 4722 11948 4738 12000
rect 4802 11948 4818 12000
rect 4882 11948 4898 12000
rect 4962 11936 4970 12000
rect 4650 11712 4692 11936
rect 4928 11712 4970 11936
rect 4650 10912 4970 11712
rect 4650 10848 4658 10912
rect 4722 10848 4738 10912
rect 4802 10848 4818 10912
rect 4882 10848 4898 10912
rect 4962 10848 4970 10912
rect 4650 9824 4970 10848
rect 4650 9760 4658 9824
rect 4722 9760 4738 9824
rect 4802 9760 4818 9824
rect 4882 9760 4898 9824
rect 4962 9760 4970 9824
rect 4650 8736 4970 9760
rect 4650 8672 4658 8736
rect 4722 8672 4738 8736
rect 4802 8672 4818 8736
rect 4882 8672 4898 8736
rect 4962 8672 4970 8736
rect 4650 8568 4970 8672
rect 4650 8332 4692 8568
rect 4928 8332 4970 8568
rect 4650 7648 4970 8332
rect 4650 7584 4658 7648
rect 4722 7584 4738 7648
rect 4802 7584 4818 7648
rect 4882 7584 4898 7648
rect 4962 7584 4970 7648
rect 4650 6560 4970 7584
rect 4650 6496 4658 6560
rect 4722 6496 4738 6560
rect 4802 6496 4818 6560
rect 4882 6496 4898 6560
rect 4962 6496 4970 6560
rect 4650 5472 4970 6496
rect 4650 5408 4658 5472
rect 4722 5408 4738 5472
rect 4802 5408 4818 5472
rect 4882 5408 4898 5472
rect 4962 5408 4970 5472
rect 4650 5188 4970 5408
rect 4650 4952 4692 5188
rect 4928 4952 4970 5188
rect 4650 4384 4970 4952
rect 4650 4320 4658 4384
rect 4722 4320 4738 4384
rect 4802 4320 4818 4384
rect 4882 4320 4898 4384
rect 4962 4320 4970 4384
rect 4650 3296 4970 4320
rect 4650 3232 4658 3296
rect 4722 3232 4738 3296
rect 4802 3232 4818 3296
rect 4882 3232 4898 3296
rect 4962 3232 4970 3296
rect 4650 2208 4970 3232
rect 4650 2144 4658 2208
rect 4722 2144 4738 2208
rect 4802 2144 4818 2208
rect 4882 2144 4898 2208
rect 4962 2144 4970 2208
rect 4650 1808 4970 2144
rect 4650 1572 4692 1808
rect 4928 1572 4970 1808
rect 4650 1120 4970 1572
rect 4650 1056 4658 1120
rect 4722 1056 4738 1120
rect 4802 1056 4818 1120
rect 4882 1056 4898 1120
rect 4962 1056 4970 1120
rect 4650 496 4970 1056
rect 6200 17984 6520 18544
rect 6200 17920 6208 17984
rect 6272 17920 6288 17984
rect 6352 17920 6368 17984
rect 6432 17920 6448 17984
rect 6512 17920 6520 17984
rect 6200 17018 6520 17920
rect 6200 16896 6242 17018
rect 6478 16896 6520 17018
rect 6200 16832 6208 16896
rect 6512 16832 6520 16896
rect 6200 16782 6242 16832
rect 6478 16782 6520 16832
rect 6200 15808 6520 16782
rect 6200 15744 6208 15808
rect 6272 15744 6288 15808
rect 6352 15744 6368 15808
rect 6432 15744 6448 15808
rect 6512 15744 6520 15808
rect 6200 14720 6520 15744
rect 6200 14656 6208 14720
rect 6272 14656 6288 14720
rect 6352 14656 6368 14720
rect 6432 14656 6448 14720
rect 6512 14656 6520 14720
rect 6200 13638 6520 14656
rect 6200 13632 6242 13638
rect 6478 13632 6520 13638
rect 6200 13568 6208 13632
rect 6512 13568 6520 13632
rect 6200 13402 6242 13568
rect 6478 13402 6520 13568
rect 6200 12544 6520 13402
rect 6200 12480 6208 12544
rect 6272 12480 6288 12544
rect 6352 12480 6368 12544
rect 6432 12480 6448 12544
rect 6512 12480 6520 12544
rect 6200 11456 6520 12480
rect 6200 11392 6208 11456
rect 6272 11392 6288 11456
rect 6352 11392 6368 11456
rect 6432 11392 6448 11456
rect 6512 11392 6520 11456
rect 6200 10368 6520 11392
rect 6200 10304 6208 10368
rect 6272 10304 6288 10368
rect 6352 10304 6368 10368
rect 6432 10304 6448 10368
rect 6512 10304 6520 10368
rect 6200 10258 6520 10304
rect 6200 10022 6242 10258
rect 6478 10022 6520 10258
rect 6200 9280 6520 10022
rect 6200 9216 6208 9280
rect 6272 9216 6288 9280
rect 6352 9216 6368 9280
rect 6432 9216 6448 9280
rect 6512 9216 6520 9280
rect 6200 8192 6520 9216
rect 6200 8128 6208 8192
rect 6272 8128 6288 8192
rect 6352 8128 6368 8192
rect 6432 8128 6448 8192
rect 6512 8128 6520 8192
rect 6200 7104 6520 8128
rect 6200 7040 6208 7104
rect 6272 7040 6288 7104
rect 6352 7040 6368 7104
rect 6432 7040 6448 7104
rect 6512 7040 6520 7104
rect 6200 6878 6520 7040
rect 6200 6642 6242 6878
rect 6478 6642 6520 6878
rect 6200 6016 6520 6642
rect 6200 5952 6208 6016
rect 6272 5952 6288 6016
rect 6352 5952 6368 6016
rect 6432 5952 6448 6016
rect 6512 5952 6520 6016
rect 6200 4928 6520 5952
rect 6200 4864 6208 4928
rect 6272 4864 6288 4928
rect 6352 4864 6368 4928
rect 6432 4864 6448 4928
rect 6512 4864 6520 4928
rect 6200 3840 6520 4864
rect 6200 3776 6208 3840
rect 6272 3776 6288 3840
rect 6352 3776 6368 3840
rect 6432 3776 6448 3840
rect 6512 3776 6520 3840
rect 6200 3498 6520 3776
rect 6200 3262 6242 3498
rect 6478 3262 6520 3498
rect 6200 2752 6520 3262
rect 6200 2688 6208 2752
rect 6272 2688 6288 2752
rect 6352 2688 6368 2752
rect 6432 2688 6448 2752
rect 6512 2688 6520 2752
rect 6200 1664 6520 2688
rect 6200 1600 6208 1664
rect 6272 1600 6288 1664
rect 6352 1600 6368 1664
rect 6432 1600 6448 1664
rect 6512 1600 6520 1664
rect 6200 576 6520 1600
rect 6200 512 6208 576
rect 6272 512 6288 576
rect 6352 512 6368 576
rect 6432 512 6448 576
rect 6512 512 6520 576
rect 6200 496 6520 512
rect 7750 18528 8070 18544
rect 7750 18464 7758 18528
rect 7822 18464 7838 18528
rect 7902 18464 7918 18528
rect 7982 18464 7998 18528
rect 8062 18464 8070 18528
rect 7750 17440 8070 18464
rect 7750 17376 7758 17440
rect 7822 17376 7838 17440
rect 7902 17376 7918 17440
rect 7982 17376 7998 17440
rect 8062 17376 8070 17440
rect 7750 16352 8070 17376
rect 7750 16288 7758 16352
rect 7822 16288 7838 16352
rect 7902 16288 7918 16352
rect 7982 16288 7998 16352
rect 8062 16288 8070 16352
rect 7750 15328 8070 16288
rect 7750 15264 7792 15328
rect 8028 15264 8070 15328
rect 7750 15200 7758 15264
rect 8062 15200 8070 15264
rect 7750 15092 7792 15200
rect 8028 15092 8070 15200
rect 7750 14176 8070 15092
rect 7750 14112 7758 14176
rect 7822 14112 7838 14176
rect 7902 14112 7918 14176
rect 7982 14112 7998 14176
rect 8062 14112 8070 14176
rect 7750 13088 8070 14112
rect 7750 13024 7758 13088
rect 7822 13024 7838 13088
rect 7902 13024 7918 13088
rect 7982 13024 7998 13088
rect 8062 13024 8070 13088
rect 7750 12000 8070 13024
rect 7750 11936 7758 12000
rect 7822 11948 7838 12000
rect 7902 11948 7918 12000
rect 7982 11948 7998 12000
rect 8062 11936 8070 12000
rect 7750 11712 7792 11936
rect 8028 11712 8070 11936
rect 7750 10912 8070 11712
rect 7750 10848 7758 10912
rect 7822 10848 7838 10912
rect 7902 10848 7918 10912
rect 7982 10848 7998 10912
rect 8062 10848 8070 10912
rect 7750 9824 8070 10848
rect 7750 9760 7758 9824
rect 7822 9760 7838 9824
rect 7902 9760 7918 9824
rect 7982 9760 7998 9824
rect 8062 9760 8070 9824
rect 7750 8736 8070 9760
rect 7750 8672 7758 8736
rect 7822 8672 7838 8736
rect 7902 8672 7918 8736
rect 7982 8672 7998 8736
rect 8062 8672 8070 8736
rect 7750 8568 8070 8672
rect 7750 8332 7792 8568
rect 8028 8332 8070 8568
rect 7750 7648 8070 8332
rect 7750 7584 7758 7648
rect 7822 7584 7838 7648
rect 7902 7584 7918 7648
rect 7982 7584 7998 7648
rect 8062 7584 8070 7648
rect 7750 6560 8070 7584
rect 7750 6496 7758 6560
rect 7822 6496 7838 6560
rect 7902 6496 7918 6560
rect 7982 6496 7998 6560
rect 8062 6496 8070 6560
rect 7750 5472 8070 6496
rect 7750 5408 7758 5472
rect 7822 5408 7838 5472
rect 7902 5408 7918 5472
rect 7982 5408 7998 5472
rect 8062 5408 8070 5472
rect 7750 5188 8070 5408
rect 7750 4952 7792 5188
rect 8028 4952 8070 5188
rect 7750 4384 8070 4952
rect 7750 4320 7758 4384
rect 7822 4320 7838 4384
rect 7902 4320 7918 4384
rect 7982 4320 7998 4384
rect 8062 4320 8070 4384
rect 7750 3296 8070 4320
rect 7750 3232 7758 3296
rect 7822 3232 7838 3296
rect 7902 3232 7918 3296
rect 7982 3232 7998 3296
rect 8062 3232 8070 3296
rect 7750 2208 8070 3232
rect 7750 2144 7758 2208
rect 7822 2144 7838 2208
rect 7902 2144 7918 2208
rect 7982 2144 7998 2208
rect 8062 2144 8070 2208
rect 7750 1808 8070 2144
rect 7750 1572 7792 1808
rect 8028 1572 8070 1808
rect 7750 1120 8070 1572
rect 7750 1056 7758 1120
rect 7822 1056 7838 1120
rect 7902 1056 7918 1120
rect 7982 1056 7998 1120
rect 8062 1056 8070 1120
rect 7750 496 8070 1056
rect 9300 17984 9620 18544
rect 9300 17920 9308 17984
rect 9372 17920 9388 17984
rect 9452 17920 9468 17984
rect 9532 17920 9548 17984
rect 9612 17920 9620 17984
rect 9300 17018 9620 17920
rect 9300 16896 9342 17018
rect 9578 16896 9620 17018
rect 9300 16832 9308 16896
rect 9612 16832 9620 16896
rect 9300 16782 9342 16832
rect 9578 16782 9620 16832
rect 9300 15808 9620 16782
rect 9300 15744 9308 15808
rect 9372 15744 9388 15808
rect 9452 15744 9468 15808
rect 9532 15744 9548 15808
rect 9612 15744 9620 15808
rect 9300 14720 9620 15744
rect 9300 14656 9308 14720
rect 9372 14656 9388 14720
rect 9452 14656 9468 14720
rect 9532 14656 9548 14720
rect 9612 14656 9620 14720
rect 9300 13638 9620 14656
rect 9300 13632 9342 13638
rect 9578 13632 9620 13638
rect 9300 13568 9308 13632
rect 9612 13568 9620 13632
rect 9300 13402 9342 13568
rect 9578 13402 9620 13568
rect 9300 12544 9620 13402
rect 9300 12480 9308 12544
rect 9372 12480 9388 12544
rect 9452 12480 9468 12544
rect 9532 12480 9548 12544
rect 9612 12480 9620 12544
rect 9300 11456 9620 12480
rect 9300 11392 9308 11456
rect 9372 11392 9388 11456
rect 9452 11392 9468 11456
rect 9532 11392 9548 11456
rect 9612 11392 9620 11456
rect 9300 10368 9620 11392
rect 9300 10304 9308 10368
rect 9372 10304 9388 10368
rect 9452 10304 9468 10368
rect 9532 10304 9548 10368
rect 9612 10304 9620 10368
rect 9300 10258 9620 10304
rect 9300 10022 9342 10258
rect 9578 10022 9620 10258
rect 9300 9280 9620 10022
rect 9300 9216 9308 9280
rect 9372 9216 9388 9280
rect 9452 9216 9468 9280
rect 9532 9216 9548 9280
rect 9612 9216 9620 9280
rect 9300 8192 9620 9216
rect 9300 8128 9308 8192
rect 9372 8128 9388 8192
rect 9452 8128 9468 8192
rect 9532 8128 9548 8192
rect 9612 8128 9620 8192
rect 9300 7104 9620 8128
rect 9300 7040 9308 7104
rect 9372 7040 9388 7104
rect 9452 7040 9468 7104
rect 9532 7040 9548 7104
rect 9612 7040 9620 7104
rect 9300 6878 9620 7040
rect 9300 6642 9342 6878
rect 9578 6642 9620 6878
rect 9300 6016 9620 6642
rect 9300 5952 9308 6016
rect 9372 5952 9388 6016
rect 9452 5952 9468 6016
rect 9532 5952 9548 6016
rect 9612 5952 9620 6016
rect 9300 4928 9620 5952
rect 9300 4864 9308 4928
rect 9372 4864 9388 4928
rect 9452 4864 9468 4928
rect 9532 4864 9548 4928
rect 9612 4864 9620 4928
rect 9300 3840 9620 4864
rect 9300 3776 9308 3840
rect 9372 3776 9388 3840
rect 9452 3776 9468 3840
rect 9532 3776 9548 3840
rect 9612 3776 9620 3840
rect 9300 3498 9620 3776
rect 9300 3262 9342 3498
rect 9578 3262 9620 3498
rect 9300 2752 9620 3262
rect 9300 2688 9308 2752
rect 9372 2688 9388 2752
rect 9452 2688 9468 2752
rect 9532 2688 9548 2752
rect 9612 2688 9620 2752
rect 9300 1664 9620 2688
rect 9300 1600 9308 1664
rect 9372 1600 9388 1664
rect 9452 1600 9468 1664
rect 9532 1600 9548 1664
rect 9612 1600 9620 1664
rect 9300 576 9620 1600
rect 9300 512 9308 576
rect 9372 512 9388 576
rect 9452 512 9468 576
rect 9532 512 9548 576
rect 9612 512 9620 576
rect 9300 496 9620 512
rect 10850 18528 11170 18544
rect 10850 18464 10858 18528
rect 10922 18464 10938 18528
rect 11002 18464 11018 18528
rect 11082 18464 11098 18528
rect 11162 18464 11170 18528
rect 10850 17440 11170 18464
rect 10850 17376 10858 17440
rect 10922 17376 10938 17440
rect 11002 17376 11018 17440
rect 11082 17376 11098 17440
rect 11162 17376 11170 17440
rect 10850 16352 11170 17376
rect 10850 16288 10858 16352
rect 10922 16288 10938 16352
rect 11002 16288 11018 16352
rect 11082 16288 11098 16352
rect 11162 16288 11170 16352
rect 10850 15328 11170 16288
rect 10850 15264 10892 15328
rect 11128 15264 11170 15328
rect 10850 15200 10858 15264
rect 11162 15200 11170 15264
rect 10850 15092 10892 15200
rect 11128 15092 11170 15200
rect 10850 14176 11170 15092
rect 10850 14112 10858 14176
rect 10922 14112 10938 14176
rect 11002 14112 11018 14176
rect 11082 14112 11098 14176
rect 11162 14112 11170 14176
rect 10850 13088 11170 14112
rect 10850 13024 10858 13088
rect 10922 13024 10938 13088
rect 11002 13024 11018 13088
rect 11082 13024 11098 13088
rect 11162 13024 11170 13088
rect 10850 12000 11170 13024
rect 10850 11936 10858 12000
rect 10922 11948 10938 12000
rect 11002 11948 11018 12000
rect 11082 11948 11098 12000
rect 11162 11936 11170 12000
rect 10850 11712 10892 11936
rect 11128 11712 11170 11936
rect 10850 10912 11170 11712
rect 10850 10848 10858 10912
rect 10922 10848 10938 10912
rect 11002 10848 11018 10912
rect 11082 10848 11098 10912
rect 11162 10848 11170 10912
rect 10850 9824 11170 10848
rect 10850 9760 10858 9824
rect 10922 9760 10938 9824
rect 11002 9760 11018 9824
rect 11082 9760 11098 9824
rect 11162 9760 11170 9824
rect 10850 8736 11170 9760
rect 10850 8672 10858 8736
rect 10922 8672 10938 8736
rect 11002 8672 11018 8736
rect 11082 8672 11098 8736
rect 11162 8672 11170 8736
rect 10850 8568 11170 8672
rect 10850 8332 10892 8568
rect 11128 8332 11170 8568
rect 10850 7648 11170 8332
rect 10850 7584 10858 7648
rect 10922 7584 10938 7648
rect 11002 7584 11018 7648
rect 11082 7584 11098 7648
rect 11162 7584 11170 7648
rect 10850 6560 11170 7584
rect 10850 6496 10858 6560
rect 10922 6496 10938 6560
rect 11002 6496 11018 6560
rect 11082 6496 11098 6560
rect 11162 6496 11170 6560
rect 10850 5472 11170 6496
rect 10850 5408 10858 5472
rect 10922 5408 10938 5472
rect 11002 5408 11018 5472
rect 11082 5408 11098 5472
rect 11162 5408 11170 5472
rect 10850 5188 11170 5408
rect 10850 4952 10892 5188
rect 11128 4952 11170 5188
rect 10850 4384 11170 4952
rect 10850 4320 10858 4384
rect 10922 4320 10938 4384
rect 11002 4320 11018 4384
rect 11082 4320 11098 4384
rect 11162 4320 11170 4384
rect 10850 3296 11170 4320
rect 10850 3232 10858 3296
rect 10922 3232 10938 3296
rect 11002 3232 11018 3296
rect 11082 3232 11098 3296
rect 11162 3232 11170 3296
rect 10850 2208 11170 3232
rect 10850 2144 10858 2208
rect 10922 2144 10938 2208
rect 11002 2144 11018 2208
rect 11082 2144 11098 2208
rect 11162 2144 11170 2208
rect 10850 1808 11170 2144
rect 10850 1572 10892 1808
rect 11128 1572 11170 1808
rect 10850 1120 11170 1572
rect 10850 1056 10858 1120
rect 10922 1056 10938 1120
rect 11002 1056 11018 1120
rect 11082 1056 11098 1120
rect 11162 1056 11170 1120
rect 10850 496 11170 1056
rect 12400 17984 12720 18544
rect 12400 17920 12408 17984
rect 12472 17920 12488 17984
rect 12552 17920 12568 17984
rect 12632 17920 12648 17984
rect 12712 17920 12720 17984
rect 12400 17018 12720 17920
rect 12400 16896 12442 17018
rect 12678 16896 12720 17018
rect 12400 16832 12408 16896
rect 12712 16832 12720 16896
rect 12400 16782 12442 16832
rect 12678 16782 12720 16832
rect 12400 15808 12720 16782
rect 12400 15744 12408 15808
rect 12472 15744 12488 15808
rect 12552 15744 12568 15808
rect 12632 15744 12648 15808
rect 12712 15744 12720 15808
rect 12400 14720 12720 15744
rect 12400 14656 12408 14720
rect 12472 14656 12488 14720
rect 12552 14656 12568 14720
rect 12632 14656 12648 14720
rect 12712 14656 12720 14720
rect 12400 13638 12720 14656
rect 12400 13632 12442 13638
rect 12678 13632 12720 13638
rect 12400 13568 12408 13632
rect 12712 13568 12720 13632
rect 12400 13402 12442 13568
rect 12678 13402 12720 13568
rect 12400 12544 12720 13402
rect 12400 12480 12408 12544
rect 12472 12480 12488 12544
rect 12552 12480 12568 12544
rect 12632 12480 12648 12544
rect 12712 12480 12720 12544
rect 12400 11456 12720 12480
rect 12400 11392 12408 11456
rect 12472 11392 12488 11456
rect 12552 11392 12568 11456
rect 12632 11392 12648 11456
rect 12712 11392 12720 11456
rect 12400 10368 12720 11392
rect 12400 10304 12408 10368
rect 12472 10304 12488 10368
rect 12552 10304 12568 10368
rect 12632 10304 12648 10368
rect 12712 10304 12720 10368
rect 12400 10258 12720 10304
rect 12400 10022 12442 10258
rect 12678 10022 12720 10258
rect 12400 9280 12720 10022
rect 12400 9216 12408 9280
rect 12472 9216 12488 9280
rect 12552 9216 12568 9280
rect 12632 9216 12648 9280
rect 12712 9216 12720 9280
rect 12400 8192 12720 9216
rect 12400 8128 12408 8192
rect 12472 8128 12488 8192
rect 12552 8128 12568 8192
rect 12632 8128 12648 8192
rect 12712 8128 12720 8192
rect 12400 7104 12720 8128
rect 12400 7040 12408 7104
rect 12472 7040 12488 7104
rect 12552 7040 12568 7104
rect 12632 7040 12648 7104
rect 12712 7040 12720 7104
rect 12400 6878 12720 7040
rect 12400 6642 12442 6878
rect 12678 6642 12720 6878
rect 12400 6016 12720 6642
rect 12400 5952 12408 6016
rect 12472 5952 12488 6016
rect 12552 5952 12568 6016
rect 12632 5952 12648 6016
rect 12712 5952 12720 6016
rect 12400 4928 12720 5952
rect 12400 4864 12408 4928
rect 12472 4864 12488 4928
rect 12552 4864 12568 4928
rect 12632 4864 12648 4928
rect 12712 4864 12720 4928
rect 12400 3840 12720 4864
rect 12400 3776 12408 3840
rect 12472 3776 12488 3840
rect 12552 3776 12568 3840
rect 12632 3776 12648 3840
rect 12712 3776 12720 3840
rect 12400 3498 12720 3776
rect 12400 3262 12442 3498
rect 12678 3262 12720 3498
rect 12400 2752 12720 3262
rect 12400 2688 12408 2752
rect 12472 2688 12488 2752
rect 12552 2688 12568 2752
rect 12632 2688 12648 2752
rect 12712 2688 12720 2752
rect 12400 1664 12720 2688
rect 12400 1600 12408 1664
rect 12472 1600 12488 1664
rect 12552 1600 12568 1664
rect 12632 1600 12648 1664
rect 12712 1600 12720 1664
rect 12400 576 12720 1600
rect 12400 512 12408 576
rect 12472 512 12488 576
rect 12552 512 12568 576
rect 12632 512 12648 576
rect 12712 512 12720 576
rect 12400 496 12720 512
rect 13950 18528 14270 18544
rect 13950 18464 13958 18528
rect 14022 18464 14038 18528
rect 14102 18464 14118 18528
rect 14182 18464 14198 18528
rect 14262 18464 14270 18528
rect 13950 17440 14270 18464
rect 13950 17376 13958 17440
rect 14022 17376 14038 17440
rect 14102 17376 14118 17440
rect 14182 17376 14198 17440
rect 14262 17376 14270 17440
rect 13950 16352 14270 17376
rect 13950 16288 13958 16352
rect 14022 16288 14038 16352
rect 14102 16288 14118 16352
rect 14182 16288 14198 16352
rect 14262 16288 14270 16352
rect 13950 15328 14270 16288
rect 13950 15264 13992 15328
rect 14228 15264 14270 15328
rect 13950 15200 13958 15264
rect 14262 15200 14270 15264
rect 13950 15092 13992 15200
rect 14228 15092 14270 15200
rect 13950 14176 14270 15092
rect 13950 14112 13958 14176
rect 14022 14112 14038 14176
rect 14102 14112 14118 14176
rect 14182 14112 14198 14176
rect 14262 14112 14270 14176
rect 13950 13088 14270 14112
rect 13950 13024 13958 13088
rect 14022 13024 14038 13088
rect 14102 13024 14118 13088
rect 14182 13024 14198 13088
rect 14262 13024 14270 13088
rect 13950 12000 14270 13024
rect 13950 11936 13958 12000
rect 14022 11948 14038 12000
rect 14102 11948 14118 12000
rect 14182 11948 14198 12000
rect 14262 11936 14270 12000
rect 13950 11712 13992 11936
rect 14228 11712 14270 11936
rect 13950 10912 14270 11712
rect 13950 10848 13958 10912
rect 14022 10848 14038 10912
rect 14102 10848 14118 10912
rect 14182 10848 14198 10912
rect 14262 10848 14270 10912
rect 13950 9824 14270 10848
rect 13950 9760 13958 9824
rect 14022 9760 14038 9824
rect 14102 9760 14118 9824
rect 14182 9760 14198 9824
rect 14262 9760 14270 9824
rect 13950 8736 14270 9760
rect 13950 8672 13958 8736
rect 14022 8672 14038 8736
rect 14102 8672 14118 8736
rect 14182 8672 14198 8736
rect 14262 8672 14270 8736
rect 13950 8568 14270 8672
rect 13950 8332 13992 8568
rect 14228 8332 14270 8568
rect 13950 7648 14270 8332
rect 13950 7584 13958 7648
rect 14022 7584 14038 7648
rect 14102 7584 14118 7648
rect 14182 7584 14198 7648
rect 14262 7584 14270 7648
rect 13950 6560 14270 7584
rect 13950 6496 13958 6560
rect 14022 6496 14038 6560
rect 14102 6496 14118 6560
rect 14182 6496 14198 6560
rect 14262 6496 14270 6560
rect 13950 5472 14270 6496
rect 13950 5408 13958 5472
rect 14022 5408 14038 5472
rect 14102 5408 14118 5472
rect 14182 5408 14198 5472
rect 14262 5408 14270 5472
rect 13950 5188 14270 5408
rect 13950 4952 13992 5188
rect 14228 4952 14270 5188
rect 13950 4384 14270 4952
rect 13950 4320 13958 4384
rect 14022 4320 14038 4384
rect 14102 4320 14118 4384
rect 14182 4320 14198 4384
rect 14262 4320 14270 4384
rect 13950 3296 14270 4320
rect 13950 3232 13958 3296
rect 14022 3232 14038 3296
rect 14102 3232 14118 3296
rect 14182 3232 14198 3296
rect 14262 3232 14270 3296
rect 13950 2208 14270 3232
rect 13950 2144 13958 2208
rect 14022 2144 14038 2208
rect 14102 2144 14118 2208
rect 14182 2144 14198 2208
rect 14262 2144 14270 2208
rect 13950 1808 14270 2144
rect 13950 1572 13992 1808
rect 14228 1572 14270 1808
rect 13950 1120 14270 1572
rect 13950 1056 13958 1120
rect 14022 1056 14038 1120
rect 14102 1056 14118 1120
rect 14182 1056 14198 1120
rect 14262 1056 14270 1120
rect 13950 496 14270 1056
rect 15500 17984 15820 18544
rect 15500 17920 15508 17984
rect 15572 17920 15588 17984
rect 15652 17920 15668 17984
rect 15732 17920 15748 17984
rect 15812 17920 15820 17984
rect 15500 17018 15820 17920
rect 15500 16896 15542 17018
rect 15778 16896 15820 17018
rect 15500 16832 15508 16896
rect 15812 16832 15820 16896
rect 15500 16782 15542 16832
rect 15778 16782 15820 16832
rect 15500 15808 15820 16782
rect 15500 15744 15508 15808
rect 15572 15744 15588 15808
rect 15652 15744 15668 15808
rect 15732 15744 15748 15808
rect 15812 15744 15820 15808
rect 15500 14720 15820 15744
rect 15500 14656 15508 14720
rect 15572 14656 15588 14720
rect 15652 14656 15668 14720
rect 15732 14656 15748 14720
rect 15812 14656 15820 14720
rect 15500 13638 15820 14656
rect 15500 13632 15542 13638
rect 15778 13632 15820 13638
rect 15500 13568 15508 13632
rect 15812 13568 15820 13632
rect 15500 13402 15542 13568
rect 15778 13402 15820 13568
rect 15500 12544 15820 13402
rect 15500 12480 15508 12544
rect 15572 12480 15588 12544
rect 15652 12480 15668 12544
rect 15732 12480 15748 12544
rect 15812 12480 15820 12544
rect 15500 11456 15820 12480
rect 15500 11392 15508 11456
rect 15572 11392 15588 11456
rect 15652 11392 15668 11456
rect 15732 11392 15748 11456
rect 15812 11392 15820 11456
rect 15500 10368 15820 11392
rect 15500 10304 15508 10368
rect 15572 10304 15588 10368
rect 15652 10304 15668 10368
rect 15732 10304 15748 10368
rect 15812 10304 15820 10368
rect 15500 10258 15820 10304
rect 15500 10022 15542 10258
rect 15778 10022 15820 10258
rect 15500 9280 15820 10022
rect 15500 9216 15508 9280
rect 15572 9216 15588 9280
rect 15652 9216 15668 9280
rect 15732 9216 15748 9280
rect 15812 9216 15820 9280
rect 15500 8192 15820 9216
rect 15500 8128 15508 8192
rect 15572 8128 15588 8192
rect 15652 8128 15668 8192
rect 15732 8128 15748 8192
rect 15812 8128 15820 8192
rect 15500 7104 15820 8128
rect 15500 7040 15508 7104
rect 15572 7040 15588 7104
rect 15652 7040 15668 7104
rect 15732 7040 15748 7104
rect 15812 7040 15820 7104
rect 15500 6878 15820 7040
rect 15500 6642 15542 6878
rect 15778 6642 15820 6878
rect 15500 6016 15820 6642
rect 15500 5952 15508 6016
rect 15572 5952 15588 6016
rect 15652 5952 15668 6016
rect 15732 5952 15748 6016
rect 15812 5952 15820 6016
rect 15500 4928 15820 5952
rect 15500 4864 15508 4928
rect 15572 4864 15588 4928
rect 15652 4864 15668 4928
rect 15732 4864 15748 4928
rect 15812 4864 15820 4928
rect 15500 3840 15820 4864
rect 15500 3776 15508 3840
rect 15572 3776 15588 3840
rect 15652 3776 15668 3840
rect 15732 3776 15748 3840
rect 15812 3776 15820 3840
rect 15500 3498 15820 3776
rect 15500 3262 15542 3498
rect 15778 3262 15820 3498
rect 15500 2752 15820 3262
rect 15500 2688 15508 2752
rect 15572 2688 15588 2752
rect 15652 2688 15668 2752
rect 15732 2688 15748 2752
rect 15812 2688 15820 2752
rect 15500 1664 15820 2688
rect 15500 1600 15508 1664
rect 15572 1600 15588 1664
rect 15652 1600 15668 1664
rect 15732 1600 15748 1664
rect 15812 1600 15820 1664
rect 15500 576 15820 1600
rect 15500 512 15508 576
rect 15572 512 15588 576
rect 15652 512 15668 576
rect 15732 512 15748 576
rect 15812 512 15820 576
rect 15500 496 15820 512
rect 17050 18528 17370 18544
rect 17050 18464 17058 18528
rect 17122 18464 17138 18528
rect 17202 18464 17218 18528
rect 17282 18464 17298 18528
rect 17362 18464 17370 18528
rect 17050 17440 17370 18464
rect 17050 17376 17058 17440
rect 17122 17376 17138 17440
rect 17202 17376 17218 17440
rect 17282 17376 17298 17440
rect 17362 17376 17370 17440
rect 17050 16352 17370 17376
rect 17050 16288 17058 16352
rect 17122 16288 17138 16352
rect 17202 16288 17218 16352
rect 17282 16288 17298 16352
rect 17362 16288 17370 16352
rect 17050 15328 17370 16288
rect 17050 15264 17092 15328
rect 17328 15264 17370 15328
rect 17050 15200 17058 15264
rect 17362 15200 17370 15264
rect 17050 15092 17092 15200
rect 17328 15092 17370 15200
rect 17050 14176 17370 15092
rect 17050 14112 17058 14176
rect 17122 14112 17138 14176
rect 17202 14112 17218 14176
rect 17282 14112 17298 14176
rect 17362 14112 17370 14176
rect 17050 13088 17370 14112
rect 17050 13024 17058 13088
rect 17122 13024 17138 13088
rect 17202 13024 17218 13088
rect 17282 13024 17298 13088
rect 17362 13024 17370 13088
rect 17050 12000 17370 13024
rect 17050 11936 17058 12000
rect 17122 11948 17138 12000
rect 17202 11948 17218 12000
rect 17282 11948 17298 12000
rect 17362 11936 17370 12000
rect 17050 11712 17092 11936
rect 17328 11712 17370 11936
rect 17050 10912 17370 11712
rect 17050 10848 17058 10912
rect 17122 10848 17138 10912
rect 17202 10848 17218 10912
rect 17282 10848 17298 10912
rect 17362 10848 17370 10912
rect 17050 9824 17370 10848
rect 17050 9760 17058 9824
rect 17122 9760 17138 9824
rect 17202 9760 17218 9824
rect 17282 9760 17298 9824
rect 17362 9760 17370 9824
rect 17050 8736 17370 9760
rect 17050 8672 17058 8736
rect 17122 8672 17138 8736
rect 17202 8672 17218 8736
rect 17282 8672 17298 8736
rect 17362 8672 17370 8736
rect 17050 8568 17370 8672
rect 17050 8332 17092 8568
rect 17328 8332 17370 8568
rect 17050 7648 17370 8332
rect 17050 7584 17058 7648
rect 17122 7584 17138 7648
rect 17202 7584 17218 7648
rect 17282 7584 17298 7648
rect 17362 7584 17370 7648
rect 17050 6560 17370 7584
rect 17050 6496 17058 6560
rect 17122 6496 17138 6560
rect 17202 6496 17218 6560
rect 17282 6496 17298 6560
rect 17362 6496 17370 6560
rect 17050 5472 17370 6496
rect 17050 5408 17058 5472
rect 17122 5408 17138 5472
rect 17202 5408 17218 5472
rect 17282 5408 17298 5472
rect 17362 5408 17370 5472
rect 17050 5188 17370 5408
rect 17050 4952 17092 5188
rect 17328 4952 17370 5188
rect 17050 4384 17370 4952
rect 17050 4320 17058 4384
rect 17122 4320 17138 4384
rect 17202 4320 17218 4384
rect 17282 4320 17298 4384
rect 17362 4320 17370 4384
rect 17050 3296 17370 4320
rect 17050 3232 17058 3296
rect 17122 3232 17138 3296
rect 17202 3232 17218 3296
rect 17282 3232 17298 3296
rect 17362 3232 17370 3296
rect 17050 2208 17370 3232
rect 17050 2144 17058 2208
rect 17122 2144 17138 2208
rect 17202 2144 17218 2208
rect 17282 2144 17298 2208
rect 17362 2144 17370 2208
rect 17050 1808 17370 2144
rect 17050 1572 17092 1808
rect 17328 1572 17370 1808
rect 17050 1120 17370 1572
rect 17050 1056 17058 1120
rect 17122 1056 17138 1120
rect 17202 1056 17218 1120
rect 17282 1056 17298 1120
rect 17362 1056 17370 1120
rect 17050 496 17370 1056
rect 18600 17984 18920 18544
rect 18600 17920 18608 17984
rect 18672 17920 18688 17984
rect 18752 17920 18768 17984
rect 18832 17920 18848 17984
rect 18912 17920 18920 17984
rect 18600 17018 18920 17920
rect 18600 16896 18642 17018
rect 18878 16896 18920 17018
rect 18600 16832 18608 16896
rect 18912 16832 18920 16896
rect 18600 16782 18642 16832
rect 18878 16782 18920 16832
rect 18600 15808 18920 16782
rect 18600 15744 18608 15808
rect 18672 15744 18688 15808
rect 18752 15744 18768 15808
rect 18832 15744 18848 15808
rect 18912 15744 18920 15808
rect 18600 14720 18920 15744
rect 18600 14656 18608 14720
rect 18672 14656 18688 14720
rect 18752 14656 18768 14720
rect 18832 14656 18848 14720
rect 18912 14656 18920 14720
rect 18600 13638 18920 14656
rect 18600 13632 18642 13638
rect 18878 13632 18920 13638
rect 18600 13568 18608 13632
rect 18912 13568 18920 13632
rect 18600 13402 18642 13568
rect 18878 13402 18920 13568
rect 18600 12544 18920 13402
rect 18600 12480 18608 12544
rect 18672 12480 18688 12544
rect 18752 12480 18768 12544
rect 18832 12480 18848 12544
rect 18912 12480 18920 12544
rect 18600 11456 18920 12480
rect 18600 11392 18608 11456
rect 18672 11392 18688 11456
rect 18752 11392 18768 11456
rect 18832 11392 18848 11456
rect 18912 11392 18920 11456
rect 18600 10368 18920 11392
rect 18600 10304 18608 10368
rect 18672 10304 18688 10368
rect 18752 10304 18768 10368
rect 18832 10304 18848 10368
rect 18912 10304 18920 10368
rect 18600 10258 18920 10304
rect 18600 10022 18642 10258
rect 18878 10022 18920 10258
rect 18600 9280 18920 10022
rect 18600 9216 18608 9280
rect 18672 9216 18688 9280
rect 18752 9216 18768 9280
rect 18832 9216 18848 9280
rect 18912 9216 18920 9280
rect 18600 8192 18920 9216
rect 18600 8128 18608 8192
rect 18672 8128 18688 8192
rect 18752 8128 18768 8192
rect 18832 8128 18848 8192
rect 18912 8128 18920 8192
rect 18600 7104 18920 8128
rect 18600 7040 18608 7104
rect 18672 7040 18688 7104
rect 18752 7040 18768 7104
rect 18832 7040 18848 7104
rect 18912 7040 18920 7104
rect 18600 6878 18920 7040
rect 18600 6642 18642 6878
rect 18878 6642 18920 6878
rect 18600 6016 18920 6642
rect 18600 5952 18608 6016
rect 18672 5952 18688 6016
rect 18752 5952 18768 6016
rect 18832 5952 18848 6016
rect 18912 5952 18920 6016
rect 18600 4928 18920 5952
rect 18600 4864 18608 4928
rect 18672 4864 18688 4928
rect 18752 4864 18768 4928
rect 18832 4864 18848 4928
rect 18912 4864 18920 4928
rect 18600 3840 18920 4864
rect 18600 3776 18608 3840
rect 18672 3776 18688 3840
rect 18752 3776 18768 3840
rect 18832 3776 18848 3840
rect 18912 3776 18920 3840
rect 18600 3498 18920 3776
rect 18600 3262 18642 3498
rect 18878 3262 18920 3498
rect 18600 2752 18920 3262
rect 18600 2688 18608 2752
rect 18672 2688 18688 2752
rect 18752 2688 18768 2752
rect 18832 2688 18848 2752
rect 18912 2688 18920 2752
rect 18600 1664 18920 2688
rect 18600 1600 18608 1664
rect 18672 1600 18688 1664
rect 18752 1600 18768 1664
rect 18832 1600 18848 1664
rect 18912 1600 18920 1664
rect 18600 576 18920 1600
rect 18600 512 18608 576
rect 18672 512 18688 576
rect 18752 512 18768 576
rect 18832 512 18848 576
rect 18912 512 18920 576
rect 18600 496 18920 512
<< via4 >>
rect 1592 15264 1828 15328
rect 1592 15200 1622 15264
rect 1622 15200 1638 15264
rect 1638 15200 1702 15264
rect 1702 15200 1718 15264
rect 1718 15200 1782 15264
rect 1782 15200 1798 15264
rect 1798 15200 1828 15264
rect 1592 15092 1828 15200
rect 1592 11936 1622 11948
rect 1622 11936 1638 11948
rect 1638 11936 1702 11948
rect 1702 11936 1718 11948
rect 1718 11936 1782 11948
rect 1782 11936 1798 11948
rect 1798 11936 1828 11948
rect 1592 11712 1828 11936
rect 1592 8332 1828 8568
rect 1592 4952 1828 5188
rect 1592 1572 1828 1808
rect 3142 16896 3378 17018
rect 3142 16832 3172 16896
rect 3172 16832 3188 16896
rect 3188 16832 3252 16896
rect 3252 16832 3268 16896
rect 3268 16832 3332 16896
rect 3332 16832 3348 16896
rect 3348 16832 3378 16896
rect 3142 16782 3378 16832
rect 3142 13632 3378 13638
rect 3142 13568 3172 13632
rect 3172 13568 3188 13632
rect 3188 13568 3252 13632
rect 3252 13568 3268 13632
rect 3268 13568 3332 13632
rect 3332 13568 3348 13632
rect 3348 13568 3378 13632
rect 3142 13402 3378 13568
rect 3142 10022 3378 10258
rect 3142 6642 3378 6878
rect 3142 3262 3378 3498
rect 4692 15264 4928 15328
rect 4692 15200 4722 15264
rect 4722 15200 4738 15264
rect 4738 15200 4802 15264
rect 4802 15200 4818 15264
rect 4818 15200 4882 15264
rect 4882 15200 4898 15264
rect 4898 15200 4928 15264
rect 4692 15092 4928 15200
rect 4692 11936 4722 11948
rect 4722 11936 4738 11948
rect 4738 11936 4802 11948
rect 4802 11936 4818 11948
rect 4818 11936 4882 11948
rect 4882 11936 4898 11948
rect 4898 11936 4928 11948
rect 4692 11712 4928 11936
rect 4692 8332 4928 8568
rect 4692 4952 4928 5188
rect 4692 1572 4928 1808
rect 6242 16896 6478 17018
rect 6242 16832 6272 16896
rect 6272 16832 6288 16896
rect 6288 16832 6352 16896
rect 6352 16832 6368 16896
rect 6368 16832 6432 16896
rect 6432 16832 6448 16896
rect 6448 16832 6478 16896
rect 6242 16782 6478 16832
rect 6242 13632 6478 13638
rect 6242 13568 6272 13632
rect 6272 13568 6288 13632
rect 6288 13568 6352 13632
rect 6352 13568 6368 13632
rect 6368 13568 6432 13632
rect 6432 13568 6448 13632
rect 6448 13568 6478 13632
rect 6242 13402 6478 13568
rect 6242 10022 6478 10258
rect 6242 6642 6478 6878
rect 6242 3262 6478 3498
rect 7792 15264 8028 15328
rect 7792 15200 7822 15264
rect 7822 15200 7838 15264
rect 7838 15200 7902 15264
rect 7902 15200 7918 15264
rect 7918 15200 7982 15264
rect 7982 15200 7998 15264
rect 7998 15200 8028 15264
rect 7792 15092 8028 15200
rect 7792 11936 7822 11948
rect 7822 11936 7838 11948
rect 7838 11936 7902 11948
rect 7902 11936 7918 11948
rect 7918 11936 7982 11948
rect 7982 11936 7998 11948
rect 7998 11936 8028 11948
rect 7792 11712 8028 11936
rect 7792 8332 8028 8568
rect 7792 4952 8028 5188
rect 7792 1572 8028 1808
rect 9342 16896 9578 17018
rect 9342 16832 9372 16896
rect 9372 16832 9388 16896
rect 9388 16832 9452 16896
rect 9452 16832 9468 16896
rect 9468 16832 9532 16896
rect 9532 16832 9548 16896
rect 9548 16832 9578 16896
rect 9342 16782 9578 16832
rect 9342 13632 9578 13638
rect 9342 13568 9372 13632
rect 9372 13568 9388 13632
rect 9388 13568 9452 13632
rect 9452 13568 9468 13632
rect 9468 13568 9532 13632
rect 9532 13568 9548 13632
rect 9548 13568 9578 13632
rect 9342 13402 9578 13568
rect 9342 10022 9578 10258
rect 9342 6642 9578 6878
rect 9342 3262 9578 3498
rect 10892 15264 11128 15328
rect 10892 15200 10922 15264
rect 10922 15200 10938 15264
rect 10938 15200 11002 15264
rect 11002 15200 11018 15264
rect 11018 15200 11082 15264
rect 11082 15200 11098 15264
rect 11098 15200 11128 15264
rect 10892 15092 11128 15200
rect 10892 11936 10922 11948
rect 10922 11936 10938 11948
rect 10938 11936 11002 11948
rect 11002 11936 11018 11948
rect 11018 11936 11082 11948
rect 11082 11936 11098 11948
rect 11098 11936 11128 11948
rect 10892 11712 11128 11936
rect 10892 8332 11128 8568
rect 10892 4952 11128 5188
rect 10892 1572 11128 1808
rect 12442 16896 12678 17018
rect 12442 16832 12472 16896
rect 12472 16832 12488 16896
rect 12488 16832 12552 16896
rect 12552 16832 12568 16896
rect 12568 16832 12632 16896
rect 12632 16832 12648 16896
rect 12648 16832 12678 16896
rect 12442 16782 12678 16832
rect 12442 13632 12678 13638
rect 12442 13568 12472 13632
rect 12472 13568 12488 13632
rect 12488 13568 12552 13632
rect 12552 13568 12568 13632
rect 12568 13568 12632 13632
rect 12632 13568 12648 13632
rect 12648 13568 12678 13632
rect 12442 13402 12678 13568
rect 12442 10022 12678 10258
rect 12442 6642 12678 6878
rect 12442 3262 12678 3498
rect 13992 15264 14228 15328
rect 13992 15200 14022 15264
rect 14022 15200 14038 15264
rect 14038 15200 14102 15264
rect 14102 15200 14118 15264
rect 14118 15200 14182 15264
rect 14182 15200 14198 15264
rect 14198 15200 14228 15264
rect 13992 15092 14228 15200
rect 13992 11936 14022 11948
rect 14022 11936 14038 11948
rect 14038 11936 14102 11948
rect 14102 11936 14118 11948
rect 14118 11936 14182 11948
rect 14182 11936 14198 11948
rect 14198 11936 14228 11948
rect 13992 11712 14228 11936
rect 13992 8332 14228 8568
rect 13992 4952 14228 5188
rect 13992 1572 14228 1808
rect 15542 16896 15778 17018
rect 15542 16832 15572 16896
rect 15572 16832 15588 16896
rect 15588 16832 15652 16896
rect 15652 16832 15668 16896
rect 15668 16832 15732 16896
rect 15732 16832 15748 16896
rect 15748 16832 15778 16896
rect 15542 16782 15778 16832
rect 15542 13632 15778 13638
rect 15542 13568 15572 13632
rect 15572 13568 15588 13632
rect 15588 13568 15652 13632
rect 15652 13568 15668 13632
rect 15668 13568 15732 13632
rect 15732 13568 15748 13632
rect 15748 13568 15778 13632
rect 15542 13402 15778 13568
rect 15542 10022 15778 10258
rect 15542 6642 15778 6878
rect 15542 3262 15778 3498
rect 17092 15264 17328 15328
rect 17092 15200 17122 15264
rect 17122 15200 17138 15264
rect 17138 15200 17202 15264
rect 17202 15200 17218 15264
rect 17218 15200 17282 15264
rect 17282 15200 17298 15264
rect 17298 15200 17328 15264
rect 17092 15092 17328 15200
rect 17092 11936 17122 11948
rect 17122 11936 17138 11948
rect 17138 11936 17202 11948
rect 17202 11936 17218 11948
rect 17218 11936 17282 11948
rect 17282 11936 17298 11948
rect 17298 11936 17328 11948
rect 17092 11712 17328 11936
rect 17092 8332 17328 8568
rect 17092 4952 17328 5188
rect 17092 1572 17328 1808
rect 18642 16896 18878 17018
rect 18642 16832 18672 16896
rect 18672 16832 18688 16896
rect 18688 16832 18752 16896
rect 18752 16832 18768 16896
rect 18768 16832 18832 16896
rect 18832 16832 18848 16896
rect 18848 16832 18878 16896
rect 18642 16782 18878 16832
rect 18642 13632 18878 13638
rect 18642 13568 18672 13632
rect 18672 13568 18688 13632
rect 18688 13568 18752 13632
rect 18752 13568 18768 13632
rect 18768 13568 18832 13632
rect 18832 13568 18848 13632
rect 18848 13568 18878 13632
rect 18642 13402 18878 13568
rect 18642 10022 18878 10258
rect 18642 6642 18878 6878
rect 18642 3262 18878 3498
<< metal5 >>
rect 136 17018 18920 17060
rect 136 16782 3142 17018
rect 3378 16782 6242 17018
rect 6478 16782 9342 17018
rect 9578 16782 12442 17018
rect 12678 16782 15542 17018
rect 15778 16782 18642 17018
rect 18878 16782 18920 17018
rect 136 16740 18920 16782
rect 136 15328 18908 15370
rect 136 15092 1592 15328
rect 1828 15092 4692 15328
rect 4928 15092 7792 15328
rect 8028 15092 10892 15328
rect 11128 15092 13992 15328
rect 14228 15092 17092 15328
rect 17328 15092 18908 15328
rect 136 15050 18908 15092
rect 136 13638 18920 13680
rect 136 13402 3142 13638
rect 3378 13402 6242 13638
rect 6478 13402 9342 13638
rect 9578 13402 12442 13638
rect 12678 13402 15542 13638
rect 15778 13402 18642 13638
rect 18878 13402 18920 13638
rect 136 13360 18920 13402
rect 136 11948 18908 11990
rect 136 11712 1592 11948
rect 1828 11712 4692 11948
rect 4928 11712 7792 11948
rect 8028 11712 10892 11948
rect 11128 11712 13992 11948
rect 14228 11712 17092 11948
rect 17328 11712 18908 11948
rect 136 11670 18908 11712
rect 136 10258 18920 10300
rect 136 10022 3142 10258
rect 3378 10022 6242 10258
rect 6478 10022 9342 10258
rect 9578 10022 12442 10258
rect 12678 10022 15542 10258
rect 15778 10022 18642 10258
rect 18878 10022 18920 10258
rect 136 9980 18920 10022
rect 136 8568 18908 8610
rect 136 8332 1592 8568
rect 1828 8332 4692 8568
rect 4928 8332 7792 8568
rect 8028 8332 10892 8568
rect 11128 8332 13992 8568
rect 14228 8332 17092 8568
rect 17328 8332 18908 8568
rect 136 8290 18908 8332
rect 136 6878 18920 6920
rect 136 6642 3142 6878
rect 3378 6642 6242 6878
rect 6478 6642 9342 6878
rect 9578 6642 12442 6878
rect 12678 6642 15542 6878
rect 15778 6642 18642 6878
rect 18878 6642 18920 6878
rect 136 6600 18920 6642
rect 136 5188 18908 5230
rect 136 4952 1592 5188
rect 1828 4952 4692 5188
rect 4928 4952 7792 5188
rect 8028 4952 10892 5188
rect 11128 4952 13992 5188
rect 14228 4952 17092 5188
rect 17328 4952 18908 5188
rect 136 4910 18908 4952
rect 136 3498 18920 3540
rect 136 3262 3142 3498
rect 3378 3262 6242 3498
rect 6478 3262 9342 3498
rect 9578 3262 12442 3498
rect 12678 3262 15542 3498
rect 15778 3262 18642 3498
rect 18878 3262 18920 3498
rect 136 3220 18920 3262
rect 136 1808 18908 1850
rect 136 1572 1592 1808
rect 1828 1572 4692 1808
rect 4928 1572 7792 1808
rect 8028 1572 10892 1808
rect 11128 1572 13992 1808
rect 14228 1572 17092 1808
rect 17328 1572 18908 1808
rect 136 1530 18908 1572
use sky130_fd_sc_hd__diode_2  ANTENNA__212__A1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 3956 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__213__A1
timestamp 1665323087
transform 1 0 1564 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__214__A1
timestamp 1665323087
transform 1 0 3956 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__215__A1
timestamp 1665323087
transform 1 0 2760 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__218__A1
timestamp 1665323087
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__219__A1
timestamp 1665323087
transform 1 0 6072 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__A1
timestamp 1665323087
transform 1 0 7820 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__221__A1
timestamp 1665323087
transform 1 0 8464 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__233__A1
timestamp 1665323087
transform 1 0 15732 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__234__A1
timestamp 1665323087
transform 1 0 14536 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__239__A1
timestamp 1665323087
transform 1 0 16652 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__A1
timestamp 1665323087
transform 1 0 16744 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__242__A0
timestamp 1665323087
transform 1 0 17572 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__A
timestamp 1665323087
transform 1 0 16376 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__265__A1
timestamp 1665323087
transform 1 0 14720 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__266__A1
timestamp 1665323087
transform 1 0 14720 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__A1
timestamp 1665323087
transform 1 0 14168 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__279__B
timestamp 1665323087
transform -1 0 6072 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__280__A2
timestamp 1665323087
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__280__B1
timestamp 1665323087
transform 1 0 4232 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__281__A2
timestamp 1665323087
transform -1 0 8372 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__281__B1
timestamp 1665323087
transform 1 0 5520 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__282__A2
timestamp 1665323087
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__282__B1
timestamp 1665323087
transform 1 0 5796 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__309__A
timestamp 1665323087
transform 1 0 2944 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__309__B
timestamp 1665323087
transform 1 0 2576 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__311__B
timestamp 1665323087
transform 1 0 4508 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__311__C
timestamp 1665323087
transform 1 0 5152 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__312__A1
timestamp 1665323087
transform 1 0 4692 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__312__A2
timestamp 1665323087
transform 1 0 4876 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__327__A
timestamp 1665323087
transform 1 0 14168 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__328__B1
timestamp 1665323087
transform -1 0 14076 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__342__A1
timestamp 1665323087
transform -1 0 18124 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__345__A_N
timestamp 1665323087
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__395__A2
timestamp 1665323087
transform 1 0 8280 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__395__B1
timestamp 1665323087
transform 1 0 8924 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__434__D
timestamp 1665323087
transform 1 0 11316 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__445__RESET_B
timestamp 1665323087
transform 1 0 16008 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__446__RESET_B
timestamp 1665323087
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__447__SET_B
timestamp 1665323087
transform 1 0 12052 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__448__RESET_B
timestamp 1665323087
transform 1 0 12420 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__450__RESET_B
timestamp 1665323087
transform 1 0 12328 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__451__SET_B
timestamp 1665323087
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__452__RESET_B
timestamp 1665323087
transform 1 0 12512 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__453__RESET_B
timestamp 1665323087
transform 1 0 13064 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__454__SET_B
timestamp 1665323087
transform 1 0 15456 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__455__RESET_B
timestamp 1665323087
transform -1 0 16100 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__459__RESET_B
timestamp 1665323087
transform 1 0 16008 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_ext_clk_A
timestamp 1665323087
transform -1 0 3680 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_pll_clk90_A
timestamp 1665323087
transform 1 0 17112 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_pll_clk_A
timestamp 1665323087
transform -1 0 8280 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout27_A
timestamp 1665323087
transform 1 0 10948 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1665323087
transform -1 0 18492 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1665323087
transform 1 0 18308 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1665323087
transform -1 0 1288 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1665323087
transform -1 0 18032 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1665323087
transform -1 0 18492 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1665323087
transform -1 0 18492 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1665323087
transform -1 0 18492 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1665323087
transform -1 0 18032 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1665323087
transform -1 0 18032 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 460 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 1196 0 1 544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 1472 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 2668 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 3404 0 1 544
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40
timestamp 1665323087
transform 1 0 3864 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53
timestamp 1665323087
transform 1 0 5060 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 5520 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64
timestamp 1665323087
transform 1 0 6072 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66
timestamp 1665323087
transform 1 0 6256 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79
timestamp 1665323087
transform 1 0 7452 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_92
timestamp 1665323087
transform 1 0 8648 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98
timestamp 1665323087
transform 1 0 9200 0 1 544
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105
timestamp 1665323087
transform 1 0 9844 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118
timestamp 1665323087
transform 1 0 11040 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_131
timestamp 1665323087
transform 1 0 12236 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_144
timestamp 1665323087
transform 1 0 13432 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_157
timestamp 1665323087
transform 1 0 14628 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_170
timestamp 1665323087
transform 1 0 15824 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_183
timestamp 1665323087
transform 1 0 17020 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_191
timestamp 1665323087
transform 1 0 17756 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_196
timestamp 1665323087
transform 1 0 18216 0 1 544
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1665323087
transform 1 0 460 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_15
timestamp 1665323087
transform 1 0 1564 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_25
timestamp 1665323087
transform 1 0 2484 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_27
timestamp 1665323087
transform 1 0 2668 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_37
timestamp 1665323087
transform 1 0 3588 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_41
timestamp 1665323087
transform 1 0 3956 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_51
timestamp 1665323087
transform 1 0 4876 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_53
timestamp 1665323087
transform 1 0 5060 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_60
timestamp 1665323087
transform 1 0 5704 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_68
timestamp 1665323087
transform 1 0 6440 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_77
timestamp 1665323087
transform 1 0 7268 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_79
timestamp 1665323087
transform 1 0 7452 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_87
timestamp 1665323087
transform 1 0 8188 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_93
timestamp 1665323087
transform 1 0 8740 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_99
timestamp 1665323087
transform 1 0 9292 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_103
timestamp 1665323087
transform 1 0 9660 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_105
timestamp 1665323087
transform 1 0 9844 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_110
timestamp 1665323087
transform 1 0 10304 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_114
timestamp 1665323087
transform 1 0 10672 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_122
timestamp 1665323087
transform 1 0 11408 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_127 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 11868 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_131
timestamp 1665323087
transform 1 0 12236 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_139
timestamp 1665323087
transform 1 0 12972 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_147
timestamp 1665323087
transform 1 0 13708 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_151
timestamp 1665323087
transform 1 0 14076 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_155
timestamp 1665323087
transform 1 0 14444 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_157
timestamp 1665323087
transform 1 0 14628 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_167
timestamp 1665323087
transform 1 0 15548 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_176
timestamp 1665323087
transform 1 0 16376 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_183
timestamp 1665323087
transform 1 0 17020 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_192
timestamp 1665323087
transform 1 0 17848 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_198
timestamp 1665323087
transform 1 0 18400 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3
timestamp 1665323087
transform 1 0 460 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_11
timestamp 1665323087
transform 1 0 1196 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_14
timestamp 1665323087
transform 1 0 1472 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_17
timestamp 1665323087
transform 1 0 1748 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_38
timestamp 1665323087
transform 1 0 3680 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_40
timestamp 1665323087
transform 1 0 3864 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_43
timestamp 1665323087
transform 1 0 4140 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_55
timestamp 1665323087
transform 1 0 5244 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_63
timestamp 1665323087
transform 1 0 5980 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_66
timestamp 1665323087
transform 1 0 6256 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_82
timestamp 1665323087
transform 1 0 7728 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_90
timestamp 1665323087
transform 1 0 8464 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_92
timestamp 1665323087
transform 1 0 8648 0 1 1632
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_105
timestamp 1665323087
transform 1 0 9844 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_118
timestamp 1665323087
transform 1 0 11040 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_128
timestamp 1665323087
transform 1 0 11960 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_139
timestamp 1665323087
transform 1 0 12972 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_144
timestamp 1665323087
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_152
timestamp 1665323087
transform 1 0 14168 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_168
timestamp 1665323087
transform 1 0 15640 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_170
timestamp 1665323087
transform 1 0 15824 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_180
timestamp 1665323087
transform 1 0 16744 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_194
timestamp 1665323087
transform 1 0 18032 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_196
timestamp 1665323087
transform 1 0 18216 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_199
timestamp 1665323087
transform 1 0 18492 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3
timestamp 1665323087
transform 1 0 460 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_13
timestamp 1665323087
transform 1 0 1380 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_24
timestamp 1665323087
transform 1 0 2392 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_27
timestamp 1665323087
transform 1 0 2668 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_30
timestamp 1665323087
transform 1 0 2944 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_42
timestamp 1665323087
transform 1 0 4048 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_50
timestamp 1665323087
transform 1 0 4784 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_53
timestamp 1665323087
transform 1 0 5060 0 -1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_65
timestamp 1665323087
transform 1 0 6164 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_77
timestamp 1665323087
transform 1 0 7268 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_79
timestamp 1665323087
transform 1 0 7452 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_85
timestamp 1665323087
transform 1 0 8004 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_96
timestamp 1665323087
transform 1 0 9016 0 -1 2720
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_105
timestamp 1665323087
transform 1 0 9844 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_117
timestamp 1665323087
transform 1 0 10948 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_129
timestamp 1665323087
transform 1 0 12052 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_131
timestamp 1665323087
transform 1 0 12236 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_139
timestamp 1665323087
transform 1 0 12972 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_145
timestamp 1665323087
transform 1 0 13524 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_150
timestamp 1665323087
transform 1 0 13984 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_154
timestamp 1665323087
transform 1 0 14352 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_157
timestamp 1665323087
transform 1 0 14628 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_172
timestamp 1665323087
transform 1 0 16008 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_178
timestamp 1665323087
transform 1 0 16560 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_181
timestamp 1665323087
transform 1 0 16836 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_183
timestamp 1665323087
transform 1 0 17020 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_194
timestamp 1665323087
transform 1 0 18032 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3
timestamp 1665323087
transform 1 0 460 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_9
timestamp 1665323087
transform 1 0 1012 0 1 2720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_14
timestamp 1665323087
transform 1 0 1472 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_26
timestamp 1665323087
transform 1 0 2576 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_38
timestamp 1665323087
transform 1 0 3680 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_40
timestamp 1665323087
transform 1 0 3864 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_61
timestamp 1665323087
transform 1 0 5796 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_66
timestamp 1665323087
transform 1 0 6256 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_71
timestamp 1665323087
transform 1 0 6716 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_82
timestamp 1665323087
transform 1 0 7728 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_90
timestamp 1665323087
transform 1 0 8464 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_92
timestamp 1665323087
transform 1 0 8648 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_102
timestamp 1665323087
transform 1 0 9568 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_116
timestamp 1665323087
transform 1 0 10856 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_118
timestamp 1665323087
transform 1 0 11040 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_125
timestamp 1665323087
transform 1 0 11684 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_142
timestamp 1665323087
transform 1 0 13248 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_144
timestamp 1665323087
transform 1 0 13432 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_156
timestamp 1665323087
transform 1 0 14536 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_168
timestamp 1665323087
transform 1 0 15640 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_170
timestamp 1665323087
transform 1 0 15824 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_178
timestamp 1665323087
transform 1 0 16560 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_182
timestamp 1665323087
transform 1 0 16928 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_193
timestamp 1665323087
transform 1 0 17940 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_196
timestamp 1665323087
transform 1 0 18216 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_199
timestamp 1665323087
transform 1 0 18492 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1665323087
transform 1 0 460 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_22
timestamp 1665323087
transform 1 0 2208 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_27
timestamp 1665323087
transform 1 0 2668 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_31
timestamp 1665323087
transform 1 0 3036 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_37
timestamp 1665323087
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_42
timestamp 1665323087
transform 1 0 4048 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_50
timestamp 1665323087
transform 1 0 4784 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_53
timestamp 1665323087
transform 1 0 5060 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_57
timestamp 1665323087
transform 1 0 5428 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_63
timestamp 1665323087
transform 1 0 5980 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_66
timestamp 1665323087
transform 1 0 6256 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_77
timestamp 1665323087
transform 1 0 7268 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_79
timestamp 1665323087
transform 1 0 7452 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_87
timestamp 1665323087
transform 1 0 8188 0 -1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_92
timestamp 1665323087
transform 1 0 8648 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_105
timestamp 1665323087
transform 1 0 9844 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_117
timestamp 1665323087
transform 1 0 10948 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_124
timestamp 1665323087
transform 1 0 11592 0 -1 3808
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_131
timestamp 1665323087
transform 1 0 12236 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_143
timestamp 1665323087
transform 1 0 13340 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_154
timestamp 1665323087
transform 1 0 14352 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_157
timestamp 1665323087
transform 1 0 14628 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_160
timestamp 1665323087
transform 1 0 14904 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_172
timestamp 1665323087
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_179
timestamp 1665323087
transform 1 0 16652 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_183
timestamp 1665323087
transform 1 0 17020 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_191
timestamp 1665323087
transform 1 0 17756 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_195
timestamp 1665323087
transform 1 0 18124 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_199
timestamp 1665323087
transform 1 0 18492 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_3
timestamp 1665323087
transform 1 0 460 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_10
timestamp 1665323087
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_14
timestamp 1665323087
transform 1 0 1472 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_26
timestamp 1665323087
transform 1 0 2576 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_38
timestamp 1665323087
transform 1 0 3680 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_40
timestamp 1665323087
transform 1 0 3864 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_44
timestamp 1665323087
transform 1 0 4232 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_51
timestamp 1665323087
transform 1 0 4876 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_63
timestamp 1665323087
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_66
timestamp 1665323087
transform 1 0 6256 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_78
timestamp 1665323087
transform 1 0 7360 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_90
timestamp 1665323087
transform 1 0 8464 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_92
timestamp 1665323087
transform 1 0 8648 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_102
timestamp 1665323087
transform 1 0 9568 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_114
timestamp 1665323087
transform 1 0 10672 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_118
timestamp 1665323087
transform 1 0 11040 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_128
timestamp 1665323087
transform 1 0 11960 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_140
timestamp 1665323087
transform 1 0 13064 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_144
timestamp 1665323087
transform 1 0 13432 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_152
timestamp 1665323087
transform 1 0 14168 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_159
timestamp 1665323087
transform 1 0 14812 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_167
timestamp 1665323087
transform 1 0 15548 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_170
timestamp 1665323087
transform 1 0 15824 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_180
timestamp 1665323087
transform 1 0 16744 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_190
timestamp 1665323087
transform 1 0 17664 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_194
timestamp 1665323087
transform 1 0 18032 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_196
timestamp 1665323087
transform 1 0 18216 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3
timestamp 1665323087
transform 1 0 460 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_24
timestamp 1665323087
transform 1 0 2392 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_27
timestamp 1665323087
transform 1 0 2668 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_31
timestamp 1665323087
transform 1 0 3036 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_38
timestamp 1665323087
transform 1 0 3680 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_46
timestamp 1665323087
transform 1 0 4416 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_51
timestamp 1665323087
transform 1 0 4876 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_53
timestamp 1665323087
transform 1 0 5060 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_65
timestamp 1665323087
transform 1 0 6164 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_73
timestamp 1665323087
transform 1 0 6900 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_77
timestamp 1665323087
transform 1 0 7268 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_79
timestamp 1665323087
transform 1 0 7452 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_91
timestamp 1665323087
transform 1 0 8556 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_103
timestamp 1665323087
transform 1 0 9660 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_105
timestamp 1665323087
transform 1 0 9844 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_127
timestamp 1665323087
transform 1 0 11868 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_131
timestamp 1665323087
transform 1 0 12236 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_152
timestamp 1665323087
transform 1 0 14168 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_157
timestamp 1665323087
transform 1 0 14628 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_162
timestamp 1665323087
transform 1 0 15088 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_170
timestamp 1665323087
transform 1 0 15824 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_173
timestamp 1665323087
transform 1 0 16100 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_181
timestamp 1665323087
transform 1 0 16836 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_183
timestamp 1665323087
transform 1 0 17020 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_195
timestamp 1665323087
transform 1 0 18124 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_199
timestamp 1665323087
transform 1 0 18492 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_3
timestamp 1665323087
transform 1 0 460 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_11
timestamp 1665323087
transform 1 0 1196 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_14
timestamp 1665323087
transform 1 0 1472 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_37
timestamp 1665323087
transform 1 0 3588 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_40
timestamp 1665323087
transform 1 0 3864 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_64
timestamp 1665323087
transform 1 0 6072 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_66
timestamp 1665323087
transform 1 0 6256 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_90
timestamp 1665323087
transform 1 0 8464 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_92
timestamp 1665323087
transform 1 0 8648 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_104
timestamp 1665323087
transform 1 0 9752 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_112
timestamp 1665323087
transform 1 0 10488 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_116
timestamp 1665323087
transform 1 0 10856 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_118
timestamp 1665323087
transform 1 0 11040 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_128
timestamp 1665323087
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_132
timestamp 1665323087
transform 1 0 12328 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_136
timestamp 1665323087
transform 1 0 12696 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_142
timestamp 1665323087
transform 1 0 13248 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_144
timestamp 1665323087
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_168
timestamp 1665323087
transform 1 0 15640 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_170
timestamp 1665323087
transform 1 0 15824 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_194
timestamp 1665323087
transform 1 0 18032 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_196
timestamp 1665323087
transform 1 0 18216 0 1 4896
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1665323087
transform 1 0 460 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_15
timestamp 1665323087
transform 1 0 1564 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_22
timestamp 1665323087
transform 1 0 2208 0 -1 5984
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1665323087
transform 1 0 2668 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_39
timestamp 1665323087
transform 1 0 3772 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_45
timestamp 1665323087
transform 1 0 4324 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_51
timestamp 1665323087
transform 1 0 4876 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_53
timestamp 1665323087
transform 1 0 5060 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_58
timestamp 1665323087
transform 1 0 5520 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_64
timestamp 1665323087
transform 1 0 6072 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_69
timestamp 1665323087
transform 1 0 6532 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_77
timestamp 1665323087
transform 1 0 7268 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_79
timestamp 1665323087
transform 1 0 7452 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_103
timestamp 1665323087
transform 1 0 9660 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_105
timestamp 1665323087
transform 1 0 9844 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_127
timestamp 1665323087
transform 1 0 11868 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_131
timestamp 1665323087
transform 1 0 12236 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_134
timestamp 1665323087
transform 1 0 12512 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_145
timestamp 1665323087
transform 1 0 13524 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_152
timestamp 1665323087
transform 1 0 14168 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_157
timestamp 1665323087
transform 1 0 14628 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_163
timestamp 1665323087
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_167
timestamp 1665323087
transform 1 0 15548 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_181
timestamp 1665323087
transform 1 0 16836 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_183
timestamp 1665323087
transform 1 0 17020 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_191
timestamp 1665323087
transform 1 0 17756 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_195
timestamp 1665323087
transform 1 0 18124 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_199
timestamp 1665323087
transform 1 0 18492 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3
timestamp 1665323087
transform 1 0 460 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_11
timestamp 1665323087
transform 1 0 1196 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_14
timestamp 1665323087
transform 1 0 1472 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_24
timestamp 1665323087
transform 1 0 2392 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_28
timestamp 1665323087
transform 1 0 2760 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_32
timestamp 1665323087
transform 1 0 3128 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_38
timestamp 1665323087
transform 1 0 3680 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_40
timestamp 1665323087
transform 1 0 3864 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_59
timestamp 1665323087
transform 1 0 5612 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_63
timestamp 1665323087
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_66
timestamp 1665323087
transform 1 0 6256 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_69
timestamp 1665323087
transform 1 0 6532 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_77
timestamp 1665323087
transform 1 0 7268 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_88
timestamp 1665323087
transform 1 0 8280 0 1 5984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_92
timestamp 1665323087
transform 1 0 8648 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_104
timestamp 1665323087
transform 1 0 9752 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_116
timestamp 1665323087
transform 1 0 10856 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_118
timestamp 1665323087
transform 1 0 11040 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_126
timestamp 1665323087
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_130
timestamp 1665323087
transform 1 0 12144 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_136
timestamp 1665323087
transform 1 0 12696 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_140
timestamp 1665323087
transform 1 0 13064 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_144
timestamp 1665323087
transform 1 0 13432 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_154
timestamp 1665323087
transform 1 0 14352 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_162
timestamp 1665323087
transform 1 0 15088 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_168
timestamp 1665323087
transform 1 0 15640 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_170
timestamp 1665323087
transform 1 0 15824 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_194
timestamp 1665323087
transform 1 0 18032 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_196
timestamp 1665323087
transform 1 0 18216 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1665323087
transform 1 0 460 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_24
timestamp 1665323087
transform 1 0 2392 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_27
timestamp 1665323087
transform 1 0 2668 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_37
timestamp 1665323087
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_48
timestamp 1665323087
transform 1 0 4600 0 -1 7072
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_53
timestamp 1665323087
transform 1 0 5060 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_65
timestamp 1665323087
transform 1 0 6164 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_73
timestamp 1665323087
transform 1 0 6900 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_77
timestamp 1665323087
transform 1 0 7268 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_79
timestamp 1665323087
transform 1 0 7452 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_88
timestamp 1665323087
transform 1 0 8280 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_93
timestamp 1665323087
transform 1 0 8740 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_97
timestamp 1665323087
transform 1 0 9108 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_103
timestamp 1665323087
transform 1 0 9660 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_105
timestamp 1665323087
transform 1 0 9844 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_128
timestamp 1665323087
transform 1 0 11960 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_131
timestamp 1665323087
transform 1 0 12236 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_152
timestamp 1665323087
transform 1 0 14168 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_157
timestamp 1665323087
transform 1 0 14628 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_167
timestamp 1665323087
transform 1 0 15548 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_179
timestamp 1665323087
transform 1 0 16652 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_183
timestamp 1665323087
transform 1 0 17020 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_190
timestamp 1665323087
transform 1 0 17664 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_194
timestamp 1665323087
transform 1 0 18032 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_199
timestamp 1665323087
transform 1 0 18492 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_3
timestamp 1665323087
transform 1 0 460 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_11
timestamp 1665323087
transform 1 0 1196 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_14
timestamp 1665323087
transform 1 0 1472 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_24
timestamp 1665323087
transform 1 0 2392 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_35
timestamp 1665323087
transform 1 0 3404 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_40
timestamp 1665323087
transform 1 0 3864 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_46
timestamp 1665323087
transform 1 0 4416 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_52
timestamp 1665323087
transform 1 0 4968 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_60
timestamp 1665323087
transform 1 0 5704 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_64
timestamp 1665323087
transform 1 0 6072 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_66
timestamp 1665323087
transform 1 0 6256 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_72
timestamp 1665323087
transform 1 0 6808 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_76
timestamp 1665323087
transform 1 0 7176 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_84
timestamp 1665323087
transform 1 0 7912 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_90
timestamp 1665323087
transform 1 0 8464 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_92
timestamp 1665323087
transform 1 0 8648 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_100
timestamp 1665323087
transform 1 0 9384 0 1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_105
timestamp 1665323087
transform 1 0 9844 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_118
timestamp 1665323087
transform 1 0 11040 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_123
timestamp 1665323087
transform 1 0 11500 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_133
timestamp 1665323087
transform 1 0 12420 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1665323087
transform 1 0 13156 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_144
timestamp 1665323087
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_148
timestamp 1665323087
transform 1 0 13800 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_160
timestamp 1665323087
transform 1 0 14904 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_168
timestamp 1665323087
transform 1 0 15640 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_170
timestamp 1665323087
transform 1 0 15824 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_12_192
timestamp 1665323087
transform 1 0 17848 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_196
timestamp 1665323087
transform 1 0 18216 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 1665323087
transform 1 0 460 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_24
timestamp 1665323087
transform 1 0 2392 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_27
timestamp 1665323087
transform 1 0 2668 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_48
timestamp 1665323087
transform 1 0 4600 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_53
timestamp 1665323087
transform 1 0 5060 0 -1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_63
timestamp 1665323087
transform 1 0 5980 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_75
timestamp 1665323087
transform 1 0 7084 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_79
timestamp 1665323087
transform 1 0 7452 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_101
timestamp 1665323087
transform 1 0 9476 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_105
timestamp 1665323087
transform 1 0 9844 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_113
timestamp 1665323087
transform 1 0 10580 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_118
timestamp 1665323087
transform 1 0 11040 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_131
timestamp 1665323087
transform 1 0 12236 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_155
timestamp 1665323087
transform 1 0 14444 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_157
timestamp 1665323087
transform 1 0 14628 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_167
timestamp 1665323087
transform 1 0 15548 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_171
timestamp 1665323087
transform 1 0 15916 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_179
timestamp 1665323087
transform 1 0 16652 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_183
timestamp 1665323087
transform 1 0 17020 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_189
timestamp 1665323087
transform 1 0 17572 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_197
timestamp 1665323087
transform 1 0 18308 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_3
timestamp 1665323087
transform 1 0 460 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_11
timestamp 1665323087
transform 1 0 1196 0 1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_14
timestamp 1665323087
transform 1 0 1472 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_26
timestamp 1665323087
transform 1 0 2576 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_36
timestamp 1665323087
transform 1 0 3496 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_40
timestamp 1665323087
transform 1 0 3864 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_47
timestamp 1665323087
transform 1 0 4508 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_53
timestamp 1665323087
transform 1 0 5060 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_58
timestamp 1665323087
transform 1 0 5520 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_64
timestamp 1665323087
transform 1 0 6072 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_66
timestamp 1665323087
transform 1 0 6256 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_74
timestamp 1665323087
transform 1 0 6992 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_86
timestamp 1665323087
transform 1 0 8096 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_90
timestamp 1665323087
transform 1 0 8464 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_92
timestamp 1665323087
transform 1 0 8648 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_104
timestamp 1665323087
transform 1 0 9752 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_116
timestamp 1665323087
transform 1 0 10856 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_118
timestamp 1665323087
transform 1 0 11040 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_123
timestamp 1665323087
transform 1 0 11500 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_134
timestamp 1665323087
transform 1 0 12512 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_142
timestamp 1665323087
transform 1 0 13248 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_144
timestamp 1665323087
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_154
timestamp 1665323087
transform 1 0 14352 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_158
timestamp 1665323087
transform 1 0 14720 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_166
timestamp 1665323087
transform 1 0 15456 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_170
timestamp 1665323087
transform 1 0 15824 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_176
timestamp 1665323087
transform 1 0 16376 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_194
timestamp 1665323087
transform 1 0 18032 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_196
timestamp 1665323087
transform 1 0 18216 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_3
timestamp 1665323087
transform 1 0 460 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_11
timestamp 1665323087
transform 1 0 1196 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_21
timestamp 1665323087
transform 1 0 2116 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_25
timestamp 1665323087
transform 1 0 2484 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_27
timestamp 1665323087
transform 1 0 2668 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_31
timestamp 1665323087
transform 1 0 3036 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_41
timestamp 1665323087
transform 1 0 3956 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_49
timestamp 1665323087
transform 1 0 4692 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_53
timestamp 1665323087
transform 1 0 5060 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_76
timestamp 1665323087
transform 1 0 7176 0 -1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_79
timestamp 1665323087
transform 1 0 7452 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_91
timestamp 1665323087
transform 1 0 8556 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_103
timestamp 1665323087
transform 1 0 9660 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_105
timestamp 1665323087
transform 1 0 9844 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_129
timestamp 1665323087
transform 1 0 12052 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_131
timestamp 1665323087
transform 1 0 12236 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_138
timestamp 1665323087
transform 1 0 12880 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_150
timestamp 1665323087
transform 1 0 13984 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_155
timestamp 1665323087
transform 1 0 14444 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_157
timestamp 1665323087
transform 1 0 14628 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_163
timestamp 1665323087
transform 1 0 15180 0 -1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1665323087
transform 1 0 15732 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_181
timestamp 1665323087
transform 1 0 16836 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_183
timestamp 1665323087
transform 1 0 17020 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_188
timestamp 1665323087
transform 1 0 17480 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_194
timestamp 1665323087
transform 1 0 18032 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_199
timestamp 1665323087
transform 1 0 18492 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_3
timestamp 1665323087
transform 1 0 460 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_11
timestamp 1665323087
transform 1 0 1196 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_14
timestamp 1665323087
transform 1 0 1472 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_16_26
timestamp 1665323087
transform 1 0 2576 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_38
timestamp 1665323087
transform 1 0 3680 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_40
timestamp 1665323087
transform 1 0 3864 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_48
timestamp 1665323087
transform 1 0 4600 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_51
timestamp 1665323087
transform 1 0 4876 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_55
timestamp 1665323087
transform 1 0 5244 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_61
timestamp 1665323087
transform 1 0 5796 0 1 9248
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_66
timestamp 1665323087
transform 1 0 6256 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_78
timestamp 1665323087
transform 1 0 7360 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_90
timestamp 1665323087
transform 1 0 8464 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_92
timestamp 1665323087
transform 1 0 8648 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1665323087
transform 1 0 9108 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_109
timestamp 1665323087
transform 1 0 10212 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_118
timestamp 1665323087
transform 1 0 11040 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_126
timestamp 1665323087
transform 1 0 11776 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_131
timestamp 1665323087
transform 1 0 12236 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_135
timestamp 1665323087
transform 1 0 12604 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_144
timestamp 1665323087
transform 1 0 13432 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_152
timestamp 1665323087
transform 1 0 14168 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_163
timestamp 1665323087
transform 1 0 15180 0 1 9248
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_170
timestamp 1665323087
transform 1 0 15824 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_182
timestamp 1665323087
transform 1 0 16928 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_194
timestamp 1665323087
transform 1 0 18032 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_196
timestamp 1665323087
transform 1 0 18216 0 1 9248
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1665323087
transform 1 0 460 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_24
timestamp 1665323087
transform 1 0 2392 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_27
timestamp 1665323087
transform 1 0 2668 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_48
timestamp 1665323087
transform 1 0 4600 0 -1 10336
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_53
timestamp 1665323087
transform 1 0 5060 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_65
timestamp 1665323087
transform 1 0 6164 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_70
timestamp 1665323087
transform 1 0 6624 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_77
timestamp 1665323087
transform 1 0 7268 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_79
timestamp 1665323087
transform 1 0 7452 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_101
timestamp 1665323087
transform 1 0 9476 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_105
timestamp 1665323087
transform 1 0 9844 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_129
timestamp 1665323087
transform 1 0 12052 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_131
timestamp 1665323087
transform 1 0 12236 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_138
timestamp 1665323087
transform 1 0 12880 0 -1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_143
timestamp 1665323087
transform 1 0 13340 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_155
timestamp 1665323087
transform 1 0 14444 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_157
timestamp 1665323087
transform 1 0 14628 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_169
timestamp 1665323087
transform 1 0 15732 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_174
timestamp 1665323087
transform 1 0 16192 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_183
timestamp 1665323087
transform 1 0 17020 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_191
timestamp 1665323087
transform 1 0 17756 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_199
timestamp 1665323087
transform 1 0 18492 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1665323087
transform 1 0 460 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_12
timestamp 1665323087
transform 1 0 1288 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_14
timestamp 1665323087
transform 1 0 1472 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_36
timestamp 1665323087
transform 1 0 3496 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_40
timestamp 1665323087
transform 1 0 3864 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_47
timestamp 1665323087
transform 1 0 4508 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_52
timestamp 1665323087
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_56
timestamp 1665323087
transform 1 0 5336 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_64
timestamp 1665323087
transform 1 0 6072 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_66
timestamp 1665323087
transform 1 0 6256 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_69
timestamp 1665323087
transform 1 0 6532 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_81
timestamp 1665323087
transform 1 0 7636 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_89
timestamp 1665323087
transform 1 0 8372 0 1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_92
timestamp 1665323087
transform 1 0 8648 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_104
timestamp 1665323087
transform 1 0 9752 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_108
timestamp 1665323087
transform 1 0 10120 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_114
timestamp 1665323087
transform 1 0 10672 0 1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_118
timestamp 1665323087
transform 1 0 11040 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_130
timestamp 1665323087
transform 1 0 12144 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_140
timestamp 1665323087
transform 1 0 13064 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_144
timestamp 1665323087
transform 1 0 13432 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_152
timestamp 1665323087
transform 1 0 14168 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_160
timestamp 1665323087
transform 1 0 14904 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_168
timestamp 1665323087
transform 1 0 15640 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_170
timestamp 1665323087
transform 1 0 15824 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_194
timestamp 1665323087
transform 1 0 18032 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_196
timestamp 1665323087
transform 1 0 18216 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_3
timestamp 1665323087
transform 1 0 460 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_20
timestamp 1665323087
transform 1 0 2024 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_27
timestamp 1665323087
transform 1 0 2668 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_35
timestamp 1665323087
transform 1 0 3404 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_49
timestamp 1665323087
transform 1 0 4692 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_53
timestamp 1665323087
transform 1 0 5060 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_74
timestamp 1665323087
transform 1 0 6992 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_79
timestamp 1665323087
transform 1 0 7452 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_103
timestamp 1665323087
transform 1 0 9660 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_105
timestamp 1665323087
transform 1 0 9844 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_113
timestamp 1665323087
transform 1 0 10580 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_123
timestamp 1665323087
transform 1 0 11500 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_129
timestamp 1665323087
transform 1 0 12052 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_131
timestamp 1665323087
transform 1 0 12236 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_152
timestamp 1665323087
transform 1 0 14168 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_157
timestamp 1665323087
transform 1 0 14628 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_167
timestamp 1665323087
transform 1 0 15548 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_174
timestamp 1665323087
transform 1 0 16192 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_180
timestamp 1665323087
transform 1 0 16744 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_183
timestamp 1665323087
transform 1 0 17020 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_190
timestamp 1665323087
transform 1 0 17664 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_194
timestamp 1665323087
transform 1 0 18032 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_199
timestamp 1665323087
transform 1 0 18492 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3
timestamp 1665323087
transform 1 0 460 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_11
timestamp 1665323087
transform 1 0 1196 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_14
timestamp 1665323087
transform 1 0 1472 0 1 11424
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_27
timestamp 1665323087
transform 1 0 2668 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_40
timestamp 1665323087
transform 1 0 3864 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_46
timestamp 1665323087
transform 1 0 4416 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_55
timestamp 1665323087
transform 1 0 5244 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_64
timestamp 1665323087
transform 1 0 6072 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_66
timestamp 1665323087
transform 1 0 6256 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_73
timestamp 1665323087
transform 1 0 6900 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_84
timestamp 1665323087
transform 1 0 7912 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_88
timestamp 1665323087
transform 1 0 8280 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_92
timestamp 1665323087
transform 1 0 8648 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_113
timestamp 1665323087
transform 1 0 10580 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_118
timestamp 1665323087
transform 1 0 11040 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_126
timestamp 1665323087
transform 1 0 11776 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_138
timestamp 1665323087
transform 1 0 12880 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_142
timestamp 1665323087
transform 1 0 13248 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_144
timestamp 1665323087
transform 1 0 13432 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_168
timestamp 1665323087
transform 1 0 15640 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_170
timestamp 1665323087
transform 1 0 15824 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_194
timestamp 1665323087
transform 1 0 18032 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_196
timestamp 1665323087
transform 1 0 18216 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_3
timestamp 1665323087
transform 1 0 460 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_25
timestamp 1665323087
transform 1 0 2484 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_27
timestamp 1665323087
transform 1 0 2668 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_33
timestamp 1665323087
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1665323087
transform 1 0 3772 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_51
timestamp 1665323087
transform 1 0 4876 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_53
timestamp 1665323087
transform 1 0 5060 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_74
timestamp 1665323087
transform 1 0 6992 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_79
timestamp 1665323087
transform 1 0 7452 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_103
timestamp 1665323087
transform 1 0 9660 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_105
timestamp 1665323087
transform 1 0 9844 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_116
timestamp 1665323087
transform 1 0 10856 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_125
timestamp 1665323087
transform 1 0 11684 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_129
timestamp 1665323087
transform 1 0 12052 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_131
timestamp 1665323087
transform 1 0 12236 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_139
timestamp 1665323087
transform 1 0 12972 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_152
timestamp 1665323087
transform 1 0 14168 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_157
timestamp 1665323087
transform 1 0 14628 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_160
timestamp 1665323087
transform 1 0 14904 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1665323087
transform 1 0 15456 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_173
timestamp 1665323087
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_179
timestamp 1665323087
transform 1 0 16652 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_183
timestamp 1665323087
transform 1 0 17020 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_186
timestamp 1665323087
transform 1 0 17296 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_198
timestamp 1665323087
transform 1 0 18400 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_3
timestamp 1665323087
transform 1 0 460 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_11
timestamp 1665323087
transform 1 0 1196 0 1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_14
timestamp 1665323087
transform 1 0 1472 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_26
timestamp 1665323087
transform 1 0 2576 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_38
timestamp 1665323087
transform 1 0 3680 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_40
timestamp 1665323087
transform 1 0 3864 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_46
timestamp 1665323087
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_53
timestamp 1665323087
transform 1 0 5060 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_61
timestamp 1665323087
transform 1 0 5796 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_66
timestamp 1665323087
transform 1 0 6256 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_80
timestamp 1665323087
transform 1 0 7544 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_86
timestamp 1665323087
transform 1 0 8096 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_90
timestamp 1665323087
transform 1 0 8464 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_92
timestamp 1665323087
transform 1 0 8648 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_113
timestamp 1665323087
transform 1 0 10580 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_118
timestamp 1665323087
transform 1 0 11040 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_140
timestamp 1665323087
transform 1 0 13064 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_144
timestamp 1665323087
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_150
timestamp 1665323087
transform 1 0 13984 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_168
timestamp 1665323087
transform 1 0 15640 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_170
timestamp 1665323087
transform 1 0 15824 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_194
timestamp 1665323087
transform 1 0 18032 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_196
timestamp 1665323087
transform 1 0 18216 0 1 12512
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1665323087
transform 1 0 460 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_15
timestamp 1665323087
transform 1 0 1564 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_23
timestamp 1665323087
transform 1 0 2300 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_27
timestamp 1665323087
transform 1 0 2668 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_51
timestamp 1665323087
transform 1 0 4876 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_53
timestamp 1665323087
transform 1 0 5060 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_61
timestamp 1665323087
transform 1 0 5796 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_68
timestamp 1665323087
transform 1 0 6440 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_77
timestamp 1665323087
transform 1 0 7268 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_79
timestamp 1665323087
transform 1 0 7452 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_103
timestamp 1665323087
transform 1 0 9660 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_105
timestamp 1665323087
transform 1 0 9844 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_129
timestamp 1665323087
transform 1 0 12052 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_131
timestamp 1665323087
transform 1 0 12236 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_155
timestamp 1665323087
transform 1 0 14444 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_157
timestamp 1665323087
transform 1 0 14628 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_165
timestamp 1665323087
transform 1 0 15364 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_170
timestamp 1665323087
transform 1 0 15824 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_174
timestamp 1665323087
transform 1 0 16192 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_178
timestamp 1665323087
transform 1 0 16560 0 -1 13600
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_183
timestamp 1665323087
transform 1 0 17020 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_195
timestamp 1665323087
transform 1 0 18124 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_199
timestamp 1665323087
transform 1 0 18492 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_3
timestamp 1665323087
transform 1 0 460 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_11
timestamp 1665323087
transform 1 0 1196 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_14
timestamp 1665323087
transform 1 0 1472 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_29
timestamp 1665323087
transform 1 0 2852 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_37
timestamp 1665323087
transform 1 0 3588 0 1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_40
timestamp 1665323087
transform 1 0 3864 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_52
timestamp 1665323087
transform 1 0 4968 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_60
timestamp 1665323087
transform 1 0 5704 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_64
timestamp 1665323087
transform 1 0 6072 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_66
timestamp 1665323087
transform 1 0 6256 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_77
timestamp 1665323087
transform 1 0 7268 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1665323087
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_89
timestamp 1665323087
transform 1 0 8372 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_92
timestamp 1665323087
transform 1 0 8648 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_113
timestamp 1665323087
transform 1 0 10580 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_118
timestamp 1665323087
transform 1 0 11040 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_129
timestamp 1665323087
transform 1 0 12052 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1665323087
transform 1 0 13156 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_144
timestamp 1665323087
transform 1 0 13432 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_157
timestamp 1665323087
transform 1 0 14628 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_165
timestamp 1665323087
transform 1 0 15364 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_170
timestamp 1665323087
transform 1 0 15824 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_177
timestamp 1665323087
transform 1 0 16468 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_183
timestamp 1665323087
transform 1 0 17020 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_189
timestamp 1665323087
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_194
timestamp 1665323087
transform 1 0 18032 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_196
timestamp 1665323087
transform 1 0 18216 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_199
timestamp 1665323087
transform 1 0 18492 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_3
timestamp 1665323087
transform 1 0 460 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_25
timestamp 1665323087
transform 1 0 2484 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_27
timestamp 1665323087
transform 1 0 2668 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_42
timestamp 1665323087
transform 1 0 4048 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_50
timestamp 1665323087
transform 1 0 4784 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1665323087
transform 1 0 5060 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_77
timestamp 1665323087
transform 1 0 7268 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_79
timestamp 1665323087
transform 1 0 7452 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_103
timestamp 1665323087
transform 1 0 9660 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_105
timestamp 1665323087
transform 1 0 9844 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_115
timestamp 1665323087
transform 1 0 10764 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_119
timestamp 1665323087
transform 1 0 11132 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_123
timestamp 1665323087
transform 1 0 11500 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_129
timestamp 1665323087
transform 1 0 12052 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_131
timestamp 1665323087
transform 1 0 12236 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_153
timestamp 1665323087
transform 1 0 14260 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_157
timestamp 1665323087
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_163
timestamp 1665323087
transform 1 0 15180 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_174
timestamp 1665323087
transform 1 0 16192 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_183
timestamp 1665323087
transform 1 0 17020 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_190
timestamp 1665323087
transform 1 0 17664 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_197
timestamp 1665323087
transform 1 0 18308 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_3
timestamp 1665323087
transform 1 0 460 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_11
timestamp 1665323087
transform 1 0 1196 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_14
timestamp 1665323087
transform 1 0 1472 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_24
timestamp 1665323087
transform 1 0 2392 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_30
timestamp 1665323087
transform 1 0 2944 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_34
timestamp 1665323087
transform 1 0 3312 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_38
timestamp 1665323087
transform 1 0 3680 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_40
timestamp 1665323087
transform 1 0 3864 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_51
timestamp 1665323087
transform 1 0 4876 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_57
timestamp 1665323087
transform 1 0 5428 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_62
timestamp 1665323087
transform 1 0 5888 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_66
timestamp 1665323087
transform 1 0 6256 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_69
timestamp 1665323087
transform 1 0 6532 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_77
timestamp 1665323087
transform 1 0 7268 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_89
timestamp 1665323087
transform 1 0 8372 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_92
timestamp 1665323087
transform 1 0 8648 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_116
timestamp 1665323087
transform 1 0 10856 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_118
timestamp 1665323087
transform 1 0 11040 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_140
timestamp 1665323087
transform 1 0 13064 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_144
timestamp 1665323087
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_161
timestamp 1665323087
transform 1 0 14996 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_170
timestamp 1665323087
transform 1 0 15824 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_180
timestamp 1665323087
transform 1 0 16744 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_186
timestamp 1665323087
transform 1 0 17296 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_190
timestamp 1665323087
transform 1 0 17664 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_194
timestamp 1665323087
transform 1 0 18032 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_196
timestamp 1665323087
transform 1 0 18216 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_3
timestamp 1665323087
transform 1 0 460 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_24
timestamp 1665323087
transform 1 0 2392 0 -1 15776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1665323087
transform 1 0 2668 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_39
timestamp 1665323087
transform 1 0 3772 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_51
timestamp 1665323087
transform 1 0 4876 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_53
timestamp 1665323087
transform 1 0 5060 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_77
timestamp 1665323087
transform 1 0 7268 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_79
timestamp 1665323087
transform 1 0 7452 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_103
timestamp 1665323087
transform 1 0 9660 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_105
timestamp 1665323087
transform 1 0 9844 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_129
timestamp 1665323087
transform 1 0 12052 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_131
timestamp 1665323087
transform 1 0 12236 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_152
timestamp 1665323087
transform 1 0 14168 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_157
timestamp 1665323087
transform 1 0 14628 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_167
timestamp 1665323087
transform 1 0 15548 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_175
timestamp 1665323087
transform 1 0 16284 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_180
timestamp 1665323087
transform 1 0 16744 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_183
timestamp 1665323087
transform 1 0 17020 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_187
timestamp 1665323087
transform 1 0 17388 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_191
timestamp 1665323087
transform 1 0 17756 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_199
timestamp 1665323087
transform 1 0 18492 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_3
timestamp 1665323087
transform 1 0 460 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_11
timestamp 1665323087
transform 1 0 1196 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_14
timestamp 1665323087
transform 1 0 1472 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_24
timestamp 1665323087
transform 1 0 2392 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_34
timestamp 1665323087
transform 1 0 3312 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_38
timestamp 1665323087
transform 1 0 3680 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_40
timestamp 1665323087
transform 1 0 3864 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_64
timestamp 1665323087
transform 1 0 6072 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_66
timestamp 1665323087
transform 1 0 6256 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_87
timestamp 1665323087
transform 1 0 8188 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_92
timestamp 1665323087
transform 1 0 8648 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_113
timestamp 1665323087
transform 1 0 10580 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_118
timestamp 1665323087
transform 1 0 11040 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_139
timestamp 1665323087
transform 1 0 12972 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_144
timestamp 1665323087
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_165
timestamp 1665323087
transform 1 0 15364 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_170
timestamp 1665323087
transform 1 0 15824 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_175
timestamp 1665323087
transform 1 0 16284 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_181
timestamp 1665323087
transform 1 0 16836 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_191
timestamp 1665323087
transform 1 0 17756 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_196
timestamp 1665323087
transform 1 0 18216 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_199
timestamp 1665323087
transform 1 0 18492 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1665323087
transform 1 0 460 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_20
timestamp 1665323087
transform 1 0 2024 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_29_27
timestamp 1665323087
transform 1 0 2668 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_33
timestamp 1665323087
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_51
timestamp 1665323087
transform 1 0 4876 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_53
timestamp 1665323087
transform 1 0 5060 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_75
timestamp 1665323087
transform 1 0 7084 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_79
timestamp 1665323087
transform 1 0 7452 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_103
timestamp 1665323087
transform 1 0 9660 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_105
timestamp 1665323087
transform 1 0 9844 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_129
timestamp 1665323087
transform 1 0 12052 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_131
timestamp 1665323087
transform 1 0 12236 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_152
timestamp 1665323087
transform 1 0 14168 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_157
timestamp 1665323087
transform 1 0 14628 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_178
timestamp 1665323087
transform 1 0 16560 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_183
timestamp 1665323087
transform 1 0 17020 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_194
timestamp 1665323087
transform 1 0 18032 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_199
timestamp 1665323087
transform 1 0 18492 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1665323087
transform 1 0 460 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_11
timestamp 1665323087
transform 1 0 1196 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_14
timestamp 1665323087
transform 1 0 1472 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_21
timestamp 1665323087
transform 1 0 2116 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_29
timestamp 1665323087
transform 1 0 2852 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_35
timestamp 1665323087
transform 1 0 3404 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_38
timestamp 1665323087
transform 1 0 3680 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_40
timestamp 1665323087
transform 1 0 3864 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_62
timestamp 1665323087
transform 1 0 5888 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_66
timestamp 1665323087
transform 1 0 6256 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_90
timestamp 1665323087
transform 1 0 8464 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_92
timestamp 1665323087
transform 1 0 8648 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_114
timestamp 1665323087
transform 1 0 10672 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_118
timestamp 1665323087
transform 1 0 11040 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_139
timestamp 1665323087
transform 1 0 12972 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_144
timestamp 1665323087
transform 1 0 13432 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_168
timestamp 1665323087
transform 1 0 15640 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_170
timestamp 1665323087
transform 1 0 15824 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_194
timestamp 1665323087
transform 1 0 18032 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_196
timestamp 1665323087
transform 1 0 18216 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1665323087
transform 1 0 460 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_25
timestamp 1665323087
transform 1 0 2484 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_27
timestamp 1665323087
transform 1 0 2668 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_48
timestamp 1665323087
transform 1 0 4600 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_53
timestamp 1665323087
transform 1 0 5060 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_74
timestamp 1665323087
transform 1 0 6992 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_79
timestamp 1665323087
transform 1 0 7452 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_103
timestamp 1665323087
transform 1 0 9660 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_105
timestamp 1665323087
transform 1 0 9844 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_127
timestamp 1665323087
transform 1 0 11868 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_131
timestamp 1665323087
transform 1 0 12236 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_152
timestamp 1665323087
transform 1 0 14168 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_157
timestamp 1665323087
transform 1 0 14628 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_179
timestamp 1665323087
transform 1 0 16652 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_183
timestamp 1665323087
transform 1 0 17020 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_193
timestamp 1665323087
transform 1 0 17940 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_199
timestamp 1665323087
transform 1 0 18492 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_3
timestamp 1665323087
transform 1 0 460 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_9
timestamp 1665323087
transform 1 0 1012 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_12
timestamp 1665323087
transform 1 0 1288 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_14
timestamp 1665323087
transform 1 0 1472 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_20
timestamp 1665323087
transform 1 0 2024 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_25
timestamp 1665323087
transform 1 0 2484 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1665323087
transform 1 0 2668 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_32
timestamp 1665323087
transform 1 0 3128 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_38
timestamp 1665323087
transform 1 0 3680 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_40
timestamp 1665323087
transform 1 0 3864 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_51
timestamp 1665323087
transform 1 0 4876 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_53
timestamp 1665323087
transform 1 0 5060 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_64
timestamp 1665323087
transform 1 0 6072 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_66
timestamp 1665323087
transform 1 0 6256 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_75
timestamp 1665323087
transform 1 0 7084 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_79
timestamp 1665323087
transform 1 0 7452 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_83
timestamp 1665323087
transform 1 0 7820 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_90
timestamp 1665323087
transform 1 0 8464 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_92
timestamp 1665323087
transform 1 0 8648 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_103
timestamp 1665323087
transform 1 0 9660 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_105
timestamp 1665323087
transform 1 0 9844 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_115
timestamp 1665323087
transform 1 0 10764 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_118
timestamp 1665323087
transform 1 0 11040 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_125
timestamp 1665323087
transform 1 0 11684 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_129
timestamp 1665323087
transform 1 0 12052 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_131
timestamp 1665323087
transform 1 0 12236 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_136
timestamp 1665323087
transform 1 0 12696 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_142
timestamp 1665323087
transform 1 0 13248 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_144
timestamp 1665323087
transform 1 0 13432 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_157
timestamp 1665323087
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_170
timestamp 1665323087
transform 1 0 15824 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_183
timestamp 1665323087
transform 1 0 17020 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_194
timestamp 1665323087
transform 1 0 18032 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_196
timestamp 1665323087
transform 1 0 18216 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_199
timestamp 1665323087
transform 1 0 18492 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1665323087
transform 1 0 184 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1665323087
transform -1 0 18860 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1665323087
transform 1 0 184 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1665323087
transform -1 0 18860 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1665323087
transform 1 0 184 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1665323087
transform -1 0 18860 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1665323087
transform 1 0 184 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1665323087
transform -1 0 18860 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1665323087
transform 1 0 184 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1665323087
transform -1 0 18860 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1665323087
transform 1 0 184 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1665323087
transform -1 0 18860 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1665323087
transform 1 0 184 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1665323087
transform -1 0 18860 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1665323087
transform 1 0 184 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1665323087
transform -1 0 18860 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1665323087
transform 1 0 184 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1665323087
transform -1 0 18860 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1665323087
transform 1 0 184 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1665323087
transform -1 0 18860 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1665323087
transform 1 0 184 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1665323087
transform -1 0 18860 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1665323087
transform 1 0 184 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1665323087
transform -1 0 18860 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1665323087
transform 1 0 184 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1665323087
transform -1 0 18860 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1665323087
transform 1 0 184 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1665323087
transform -1 0 18860 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1665323087
transform 1 0 184 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1665323087
transform -1 0 18860 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1665323087
transform 1 0 184 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1665323087
transform -1 0 18860 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1665323087
transform 1 0 184 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1665323087
transform -1 0 18860 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1665323087
transform 1 0 184 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1665323087
transform -1 0 18860 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1665323087
transform 1 0 184 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1665323087
transform -1 0 18860 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1665323087
transform 1 0 184 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1665323087
transform -1 0 18860 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1665323087
transform 1 0 184 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1665323087
transform -1 0 18860 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1665323087
transform 1 0 184 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1665323087
transform -1 0 18860 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1665323087
transform 1 0 184 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1665323087
transform -1 0 18860 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1665323087
transform 1 0 184 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1665323087
transform -1 0 18860 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1665323087
transform 1 0 184 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1665323087
transform -1 0 18860 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1665323087
transform 1 0 184 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1665323087
transform -1 0 18860 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1665323087
transform 1 0 184 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1665323087
transform -1 0 18860 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1665323087
transform 1 0 184 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1665323087
transform -1 0 18860 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1665323087
transform 1 0 184 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1665323087
transform -1 0 18860 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1665323087
transform 1 0 184 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1665323087
transform -1 0 18860 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1665323087
transform 1 0 184 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1665323087
transform -1 0 18860 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1665323087
transform 1 0 184 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1665323087
transform -1 0 18860 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1665323087
transform 1 0 184 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1665323087
transform -1 0 18860 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 1380 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1665323087
transform 1 0 2576 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1665323087
transform 1 0 3772 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1665323087
transform 1 0 4968 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1665323087
transform 1 0 6164 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1665323087
transform 1 0 7360 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1665323087
transform 1 0 8556 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1665323087
transform 1 0 9752 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1665323087
transform 1 0 10948 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1665323087
transform 1 0 12144 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1665323087
transform 1 0 13340 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1665323087
transform 1 0 14536 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1665323087
transform 1 0 15732 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1665323087
transform 1 0 16928 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1665323087
transform 1 0 18124 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1665323087
transform 1 0 2576 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1665323087
transform 1 0 4968 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1665323087
transform 1 0 7360 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1665323087
transform 1 0 9752 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1665323087
transform 1 0 12144 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1665323087
transform 1 0 14536 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1665323087
transform 1 0 16928 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1665323087
transform 1 0 1380 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1665323087
transform 1 0 3772 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1665323087
transform 1 0 6164 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1665323087
transform 1 0 8556 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1665323087
transform 1 0 10948 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1665323087
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1665323087
transform 1 0 15732 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1665323087
transform 1 0 18124 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1665323087
transform 1 0 2576 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1665323087
transform 1 0 4968 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1665323087
transform 1 0 7360 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1665323087
transform 1 0 9752 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1665323087
transform 1 0 12144 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1665323087
transform 1 0 14536 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1665323087
transform 1 0 16928 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1665323087
transform 1 0 1380 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1665323087
transform 1 0 3772 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1665323087
transform 1 0 6164 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1665323087
transform 1 0 8556 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1665323087
transform 1 0 10948 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1665323087
transform 1 0 13340 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1665323087
transform 1 0 15732 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1665323087
transform 1 0 18124 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1665323087
transform 1 0 2576 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1665323087
transform 1 0 4968 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1665323087
transform 1 0 7360 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1665323087
transform 1 0 9752 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1665323087
transform 1 0 12144 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1665323087
transform 1 0 14536 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1665323087
transform 1 0 16928 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1665323087
transform 1 0 1380 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1665323087
transform 1 0 3772 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1665323087
transform 1 0 6164 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1665323087
transform 1 0 8556 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1665323087
transform 1 0 10948 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1665323087
transform 1 0 13340 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1665323087
transform 1 0 15732 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1665323087
transform 1 0 18124 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1665323087
transform 1 0 2576 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1665323087
transform 1 0 4968 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1665323087
transform 1 0 7360 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1665323087
transform 1 0 9752 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1665323087
transform 1 0 12144 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1665323087
transform 1 0 14536 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1665323087
transform 1 0 16928 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1665323087
transform 1 0 1380 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1665323087
transform 1 0 3772 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1665323087
transform 1 0 6164 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1665323087
transform 1 0 8556 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1665323087
transform 1 0 10948 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1665323087
transform 1 0 13340 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1665323087
transform 1 0 15732 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1665323087
transform 1 0 18124 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1665323087
transform 1 0 2576 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1665323087
transform 1 0 4968 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1665323087
transform 1 0 7360 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1665323087
transform 1 0 9752 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1665323087
transform 1 0 12144 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1665323087
transform 1 0 14536 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1665323087
transform 1 0 16928 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1665323087
transform 1 0 1380 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1665323087
transform 1 0 3772 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1665323087
transform 1 0 6164 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1665323087
transform 1 0 8556 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1665323087
transform 1 0 10948 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1665323087
transform 1 0 13340 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1665323087
transform 1 0 15732 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1665323087
transform 1 0 18124 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1665323087
transform 1 0 2576 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1665323087
transform 1 0 4968 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1665323087
transform 1 0 7360 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1665323087
transform 1 0 9752 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1665323087
transform 1 0 12144 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1665323087
transform 1 0 14536 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1665323087
transform 1 0 16928 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1665323087
transform 1 0 1380 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1665323087
transform 1 0 3772 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1665323087
transform 1 0 6164 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1665323087
transform 1 0 8556 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1665323087
transform 1 0 10948 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1665323087
transform 1 0 13340 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1665323087
transform 1 0 15732 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1665323087
transform 1 0 18124 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1665323087
transform 1 0 2576 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1665323087
transform 1 0 4968 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1665323087
transform 1 0 7360 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1665323087
transform 1 0 9752 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1665323087
transform 1 0 12144 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1665323087
transform 1 0 14536 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1665323087
transform 1 0 16928 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1665323087
transform 1 0 1380 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1665323087
transform 1 0 3772 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1665323087
transform 1 0 6164 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1665323087
transform 1 0 8556 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1665323087
transform 1 0 10948 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1665323087
transform 1 0 13340 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1665323087
transform 1 0 15732 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1665323087
transform 1 0 18124 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1665323087
transform 1 0 2576 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1665323087
transform 1 0 4968 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1665323087
transform 1 0 7360 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1665323087
transform 1 0 9752 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1665323087
transform 1 0 12144 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1665323087
transform 1 0 14536 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1665323087
transform 1 0 16928 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1665323087
transform 1 0 1380 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1665323087
transform 1 0 3772 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1665323087
transform 1 0 6164 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1665323087
transform 1 0 8556 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1665323087
transform 1 0 10948 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1665323087
transform 1 0 13340 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1665323087
transform 1 0 15732 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1665323087
transform 1 0 18124 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1665323087
transform 1 0 2576 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1665323087
transform 1 0 4968 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1665323087
transform 1 0 7360 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1665323087
transform 1 0 9752 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1665323087
transform 1 0 12144 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1665323087
transform 1 0 14536 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1665323087
transform 1 0 16928 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1665323087
transform 1 0 1380 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1665323087
transform 1 0 3772 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1665323087
transform 1 0 6164 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1665323087
transform 1 0 8556 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1665323087
transform 1 0 10948 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1665323087
transform 1 0 13340 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1665323087
transform 1 0 15732 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1665323087
transform 1 0 18124 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1665323087
transform 1 0 2576 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1665323087
transform 1 0 4968 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1665323087
transform 1 0 7360 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1665323087
transform 1 0 9752 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1665323087
transform 1 0 12144 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1665323087
transform 1 0 14536 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1665323087
transform 1 0 16928 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1665323087
transform 1 0 1380 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1665323087
transform 1 0 3772 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1665323087
transform 1 0 6164 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1665323087
transform 1 0 8556 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1665323087
transform 1 0 10948 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1665323087
transform 1 0 13340 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1665323087
transform 1 0 15732 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1665323087
transform 1 0 18124 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1665323087
transform 1 0 2576 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1665323087
transform 1 0 4968 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1665323087
transform 1 0 7360 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1665323087
transform 1 0 9752 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1665323087
transform 1 0 12144 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1665323087
transform 1 0 14536 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1665323087
transform 1 0 16928 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1665323087
transform 1 0 1380 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1665323087
transform 1 0 3772 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1665323087
transform 1 0 6164 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1665323087
transform 1 0 8556 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1665323087
transform 1 0 10948 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1665323087
transform 1 0 13340 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1665323087
transform 1 0 15732 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1665323087
transform 1 0 18124 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1665323087
transform 1 0 2576 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1665323087
transform 1 0 4968 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1665323087
transform 1 0 7360 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1665323087
transform 1 0 9752 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1665323087
transform 1 0 12144 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1665323087
transform 1 0 14536 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1665323087
transform 1 0 16928 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1665323087
transform 1 0 1380 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1665323087
transform 1 0 3772 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1665323087
transform 1 0 6164 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1665323087
transform 1 0 8556 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1665323087
transform 1 0 10948 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1665323087
transform 1 0 13340 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1665323087
transform 1 0 15732 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1665323087
transform 1 0 18124 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1665323087
transform 1 0 2576 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1665323087
transform 1 0 4968 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1665323087
transform 1 0 7360 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1665323087
transform 1 0 9752 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1665323087
transform 1 0 12144 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1665323087
transform 1 0 14536 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1665323087
transform 1 0 16928 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1665323087
transform 1 0 1380 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1665323087
transform 1 0 3772 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1665323087
transform 1 0 6164 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1665323087
transform 1 0 8556 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1665323087
transform 1 0 10948 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1665323087
transform 1 0 13340 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1665323087
transform 1 0 15732 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1665323087
transform 1 0 18124 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1665323087
transform 1 0 2576 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1665323087
transform 1 0 4968 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1665323087
transform 1 0 7360 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1665323087
transform 1 0 9752 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1665323087
transform 1 0 12144 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1665323087
transform 1 0 14536 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1665323087
transform 1 0 16928 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1665323087
transform 1 0 1380 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1665323087
transform 1 0 3772 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1665323087
transform 1 0 6164 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1665323087
transform 1 0 8556 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1665323087
transform 1 0 10948 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1665323087
transform 1 0 13340 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1665323087
transform 1 0 15732 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1665323087
transform 1 0 18124 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1665323087
transform 1 0 2576 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1665323087
transform 1 0 4968 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1665323087
transform 1 0 7360 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1665323087
transform 1 0 9752 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1665323087
transform 1 0 12144 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1665323087
transform 1 0 14536 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1665323087
transform 1 0 16928 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1665323087
transform 1 0 1380 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1665323087
transform 1 0 3772 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1665323087
transform 1 0 6164 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1665323087
transform 1 0 8556 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1665323087
transform 1 0 10948 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1665323087
transform 1 0 13340 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1665323087
transform 1 0 15732 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1665323087
transform 1 0 18124 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1665323087
transform 1 0 2576 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1665323087
transform 1 0 4968 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1665323087
transform 1 0 7360 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1665323087
transform 1 0 9752 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1665323087
transform 1 0 12144 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1665323087
transform 1 0 14536 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1665323087
transform 1 0 16928 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1665323087
transform 1 0 1380 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1665323087
transform 1 0 2576 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1665323087
transform 1 0 3772 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1665323087
transform 1 0 4968 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1665323087
transform 1 0 6164 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1665323087
transform 1 0 7360 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1665323087
transform 1 0 8556 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1665323087
transform 1 0 9752 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1665323087
transform 1 0 10948 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1665323087
transform 1 0 12144 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1665323087
transform 1 0 13340 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1665323087
transform 1 0 14536 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1665323087
transform 1 0 15732 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1665323087
transform 1 0 16928 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1665323087
transform 1 0 18124 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _202_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 3772 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _203_
timestamp 1665323087
transform 1 0 12696 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _204_
timestamp 1665323087
transform 1 0 7084 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _205_
timestamp 1665323087
transform -1 0 6072 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _206_
timestamp 1665323087
transform -1 0 8372 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _207_
timestamp 1665323087
transform -1 0 14628 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _208_
timestamp 1665323087
transform -1 0 10764 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _209_
timestamp 1665323087
transform 1 0 2760 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _210_
timestamp 1665323087
transform 1 0 2852 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _211_
timestamp 1665323087
transform 1 0 3128 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _212_
timestamp 1665323087
transform 1 0 2760 0 -1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _213_
timestamp 1665323087
transform 1 0 552 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _214_
timestamp 1665323087
transform 1 0 2852 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _215_
timestamp 1665323087
transform 1 0 1564 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _216_
timestamp 1665323087
transform 1 0 5336 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _217_
timestamp 1665323087
transform 1 0 4968 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _218_
timestamp 1665323087
transform 1 0 6900 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _219_
timestamp 1665323087
transform 1 0 6440 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _220_
timestamp 1665323087
transform 1 0 8188 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _221_
timestamp 1665323087
transform 1 0 7636 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _222_
timestamp 1665323087
transform 1 0 8740 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _223_
timestamp 1665323087
transform 1 0 8740 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _224_
timestamp 1665323087
transform 1 0 2024 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _225_
timestamp 1665323087
transform 1 0 3220 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _226_
timestamp 1665323087
transform -1 0 11960 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _227_
timestamp 1665323087
transform 1 0 12144 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _228_
timestamp 1665323087
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _229_
timestamp 1665323087
transform 1 0 14720 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _230_
timestamp 1665323087
transform 1 0 14076 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _231_
timestamp 1665323087
transform 1 0 14720 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _232_
timestamp 1665323087
transform 1 0 13340 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _233_
timestamp 1665323087
transform 1 0 14720 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _234_
timestamp 1665323087
transform 1 0 13524 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _235_
timestamp 1665323087
transform 1 0 15180 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _236_
timestamp 1665323087
transform 1 0 14812 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _237_
timestamp 1665323087
transform -1 0 16744 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _238_
timestamp 1665323087
transform 1 0 15916 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _239_
timestamp 1665323087
transform 1 0 17204 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _240_
timestamp 1665323087
transform 1 0 17112 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _241_
timestamp 1665323087
transform 1 0 15916 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _242_
timestamp 1665323087
transform 1 0 17204 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_4  _243_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 12328 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  _244_
timestamp 1665323087
transform 1 0 6348 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  _245_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 2944 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _246_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 3128 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _247_
timestamp 1665323087
transform -1 0 2484 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_4  _248_
timestamp 1665323087
transform 1 0 7544 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  _249_
timestamp 1665323087
transform -1 0 15180 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _250_
timestamp 1665323087
transform -1 0 11868 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _251_
timestamp 1665323087
transform 1 0 14720 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_4  _252_
timestamp 1665323087
transform 1 0 15732 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  _253_
timestamp 1665323087
transform -1 0 9844 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__inv_4  _254__7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 9200 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _255_
timestamp 1665323087
transform 1 0 736 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  _256__4
timestamp 1665323087
transform -1 0 2208 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _257_
timestamp 1665323087
transform 1 0 5152 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _258_
timestamp 1665323087
transform -1 0 13800 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  _259__1
timestamp 1665323087
transform -1 0 10672 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _260_
timestamp 1665323087
transform -1 0 12512 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _261_
timestamp 1665323087
transform 1 0 11132 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__nor3b_2  _262_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 15180 0 1 9248
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_2  _263_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 11132 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _264_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 15548 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_2  _265_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 14352 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _266_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 13524 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_4  _267_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 14168 0 -1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _268_
timestamp 1665323087
transform 1 0 12788 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _269_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 11132 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__a41oi_1  _270_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 10856 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _271_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 10580 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _272_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 11040 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _273_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 12880 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _274_
timestamp 1665323087
transform -1 0 13340 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2ai_1  _275_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 12420 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _276_
timestamp 1665323087
transform 1 0 1564 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__nor3b_2  _277_
timestamp 1665323087
transform 1 0 4324 0 1 1632
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_2  _278_
timestamp 1665323087
transform 1 0 3956 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _279_
timestamp 1665323087
transform -1 0 6440 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _280_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 5520 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _281_
timestamp 1665323087
transform -1 0 7268 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_4  _282_
timestamp 1665323087
transform -1 0 5612 0 1 5984
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _283_
timestamp 1665323087
transform -1 0 4324 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _284_
timestamp 1665323087
transform 1 0 5336 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__a41oi_1  _285_
timestamp 1665323087
transform -1 0 5704 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _286_
timestamp 1665323087
transform -1 0 5520 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _287_
timestamp 1665323087
transform 1 0 5152 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _288_
timestamp 1665323087
transform -1 0 3588 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _289_
timestamp 1665323087
transform -1 0 4048 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2ai_1  _290_
timestamp 1665323087
transform 1 0 1564 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _291_
timestamp 1665323087
transform -1 0 3220 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _292_
timestamp 1665323087
transform 1 0 3404 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _293_
timestamp 1665323087
transform -1 0 6900 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _294_
timestamp 1665323087
transform 1 0 9568 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _295_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 7728 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _296_
timestamp 1665323087
transform 1 0 17388 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _297_
timestamp 1665323087
transform -1 0 17388 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _298_
timestamp 1665323087
transform 1 0 13708 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _299_
timestamp 1665323087
transform -1 0 15548 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _300_
timestamp 1665323087
transform 1 0 14904 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_2  _301_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 6624 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _302_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 6808 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _303_
timestamp 1665323087
transform -1 0 6624 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_2  _304_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 6624 0 1 12512
box -38 -48 958 592
use sky130_fd_sc_hd__nand2b_2  _305_
timestamp 1665323087
transform -1 0 15364 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _306_
timestamp 1665323087
transform -1 0 13984 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _307_
timestamp 1665323087
transform -1 0 12052 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_2  _308_
timestamp 1665323087
transform 1 0 12236 0 1 13600
box -38 -48 958 592
use sky130_fd_sc_hd__xnor2_1  _309_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 1748 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _310_
timestamp 1665323087
transform 1 0 2760 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _311_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 4508 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _312_
timestamp 1665323087
transform 1 0 4140 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _313_
timestamp 1665323087
transform 1 0 4692 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _314_
timestamp 1665323087
transform -1 0 3496 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _315_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 3956 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _316_
timestamp 1665323087
transform 1 0 2760 0 1 544
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _317_
timestamp 1665323087
transform -1 0 5520 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _318_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 4508 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _319_
timestamp 1665323087
transform 1 0 5244 0 -1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _320_
timestamp 1665323087
transform 1 0 6624 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _321_
timestamp 1665323087
transform 1 0 9936 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _322_
timestamp 1665323087
transform -1 0 9200 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _323_
timestamp 1665323087
transform -1 0 9292 0 -1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _324_
timestamp 1665323087
transform 1 0 2668 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _325_
timestamp 1665323087
transform -1 0 14168 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _326_
timestamp 1665323087
transform 1 0 10764 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _327_
timestamp 1665323087
transform 1 0 13156 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _328_
timestamp 1665323087
transform 1 0 13156 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _329_
timestamp 1665323087
transform 1 0 13708 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _330_
timestamp 1665323087
transform 1 0 11132 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _331_
timestamp 1665323087
transform 1 0 10304 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _332_
timestamp 1665323087
transform 1 0 14260 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _333_
timestamp 1665323087
transform -1 0 14444 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _334_
timestamp 1665323087
transform -1 0 15732 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _335_
timestamp 1665323087
transform 1 0 14720 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _336_
timestamp 1665323087
transform 1 0 14904 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _337_
timestamp 1665323087
transform 1 0 18032 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _338_
timestamp 1665323087
transform -1 0 17756 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _339_
timestamp 1665323087
transform -1 0 17848 0 -1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _340_
timestamp 1665323087
transform 1 0 17112 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _341_
timestamp 1665323087
transform 1 0 12420 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__o2111ai_2  _342_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 15732 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__a21oi_1  _343_
timestamp 1665323087
transform 1 0 16376 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _344_
timestamp 1665323087
transform 1 0 15824 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nand4bb_1  _345_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 4876 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _346_
timestamp 1665323087
transform 1 0 5060 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _347_
timestamp 1665323087
transform -1 0 5888 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _348_
timestamp 1665323087
transform 1 0 2208 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _349_
timestamp 1665323087
transform 1 0 2760 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _350_
timestamp 1665323087
transform -1 0 4416 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _351_
timestamp 1665323087
transform 1 0 4600 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _352_
timestamp 1665323087
transform 1 0 5428 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _353_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 3404 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _354_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 5244 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _355_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 3680 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _356_
timestamp 1665323087
transform 1 0 736 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_1  _357_
timestamp 1665323087
transform 1 0 4324 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _358_
timestamp 1665323087
transform -1 0 4876 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _359_
timestamp 1665323087
transform 1 0 1564 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _360_
timestamp 1665323087
transform 1 0 1288 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _361_
timestamp 1665323087
transform 1 0 6164 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _362_
timestamp 1665323087
transform -1 0 6900 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _363_
timestamp 1665323087
transform 1 0 6900 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _364_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 8280 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _365_
timestamp 1665323087
transform -1 0 8740 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _366_
timestamp 1665323087
transform 1 0 7544 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _367_
timestamp 1665323087
transform 1 0 1564 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _368_
timestamp 1665323087
transform 1 0 1564 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__nor4_1  _369_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 1564 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__o31ai_1  _370_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 2116 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _371_
timestamp 1665323087
transform 1 0 1564 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _372_
timestamp 1665323087
transform 1 0 4048 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__nand4bb_1  _373_
timestamp 1665323087
transform -1 0 16192 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _374_
timestamp 1665323087
transform -1 0 16284 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _375_
timestamp 1665323087
transform -1 0 16744 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _376_
timestamp 1665323087
transform 1 0 15916 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _377_
timestamp 1665323087
transform 1 0 17112 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _378_
timestamp 1665323087
transform -1 0 17480 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _379_
timestamp 1665323087
transform -1 0 15456 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _380_
timestamp 1665323087
transform 1 0 15640 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _381_
timestamp 1665323087
transform 1 0 16284 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _382_
timestamp 1665323087
transform 1 0 17112 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _383_
timestamp 1665323087
transform -1 0 12420 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _384_
timestamp 1665323087
transform -1 0 11500 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_1  _385_
timestamp 1665323087
transform -1 0 12880 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _386_
timestamp 1665323087
transform -1 0 11500 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _387_
timestamp 1665323087
transform 1 0 11132 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _388_
timestamp 1665323087
transform -1 0 13064 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _389_
timestamp 1665323087
transform 1 0 14444 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _390_
timestamp 1665323087
transform -1 0 15088 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _391_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 16100 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _392_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 17112 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _393_
timestamp 1665323087
transform 1 0 17204 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _394_
timestamp 1665323087
transform 1 0 17020 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__o2111ai_1  _395_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 9384 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _396_
timestamp 1665323087
transform 1 0 8740 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _397_
timestamp 1665323087
transform 1 0 8096 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _398_
timestamp 1665323087
transform 1 0 14720 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _399_
timestamp 1665323087
transform 1 0 17112 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__nor4_1  _400_
timestamp 1665323087
transform -1 0 18308 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__o31ai_1  _401_
timestamp 1665323087
transform -1 0 17664 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _402_
timestamp 1665323087
transform -1 0 17572 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _403__8
timestamp 1665323087
transform 1 0 8004 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _404__9
timestamp 1665323087
transform -1 0 7084 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _405__5
timestamp 1665323087
transform -1 0 5796 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _406__6
timestamp 1665323087
transform 1 0 828 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _407__2
timestamp 1665323087
transform -1 0 11684 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _408__3
timestamp 1665323087
transform -1 0 10488 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__dfstp_1  _409_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 9936 0 -1 17952
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _410_
timestamp 1665323087
transform 1 0 8740 0 1 16864
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _411__30 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 7820 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _411_
timestamp 1665323087
transform 1 0 6532 0 1 16864
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _412_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 9660 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _413_
timestamp 1665323087
transform 1 0 5428 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _414_
timestamp 1665323087
transform 1 0 16100 0 1 11424
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _415_
timestamp 1665323087
transform 1 0 4048 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _416_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 552 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _417_
timestamp 1665323087
transform 1 0 1012 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _418_
timestamp 1665323087
transform 1 0 3404 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfstp_1  _419_
timestamp 1665323087
transform 1 0 5336 0 -1 14688
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _420_
timestamp 1665323087
transform 1 0 5152 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtn_1  _421_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 552 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _422_
timestamp 1665323087
transform 1 0 1656 0 1 4896
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtn_1  _423_
timestamp 1665323087
transform 1 0 4232 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _424_
timestamp 1665323087
transform 1 0 5244 0 -1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtn_1  _425_
timestamp 1665323087
transform 1 0 552 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _426_
timestamp 1665323087
transform 1 0 1564 0 1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtn_1  _427_
timestamp 1665323087
transform 1 0 552 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _428_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 6348 0 1 4896
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_2  _429_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 7544 0 -1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _430_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 7728 0 -1 5984
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _431_
timestamp 1665323087
transform 1 0 552 0 -1 14688
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _432_
timestamp 1665323087
transform 1 0 552 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _433_
timestamp 1665323087
transform 1 0 644 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _434_
timestamp 1665323087
transform 1 0 7820 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _435_
timestamp 1665323087
transform -1 0 9660 0 -1 13600
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _436_
timestamp 1665323087
transform -1 0 10580 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _437_
timestamp 1665323087
transform -1 0 10580 0 1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _438_
timestamp 1665323087
transform 1 0 7728 0 -1 14688
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _439_
timestamp 1665323087
transform -1 0 10580 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _440_
timestamp 1665323087
transform 1 0 3404 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _441_
timestamp 1665323087
transform 1 0 16560 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _442_
timestamp 1665323087
transform 1 0 16376 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _443_
timestamp 1665323087
transform 1 0 14168 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfstp_1  _444_
timestamp 1665323087
transform -1 0 15640 0 1 16864
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _445_
timestamp 1665323087
transform 1 0 16192 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtn_1  _446_
timestamp 1665323087
transform 1 0 10120 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _447_
timestamp 1665323087
transform 1 0 10120 0 -1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtn_1  _448_
timestamp 1665323087
transform 1 0 10212 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _449_
timestamp 1665323087
transform 1 0 11132 0 1 12512
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtn_1  _450_
timestamp 1665323087
transform 1 0 10028 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _451_
timestamp 1665323087
transform 1 0 9936 0 -1 4896
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtn_1  _452_
timestamp 1665323087
transform -1 0 14168 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _453_
timestamp 1665323087
transform 1 0 13524 0 1 4896
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_2  _454_
timestamp 1665323087
transform 1 0 16100 0 1 5984
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _455_
timestamp 1665323087
transform 1 0 16100 0 1 4896
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _456_
timestamp 1665323087
transform 1 0 7544 0 -1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _457_
timestamp 1665323087
transform 1 0 14720 0 -1 17952
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _458_
timestamp 1665323087
transform 1 0 16192 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _459_
timestamp 1665323087
transform 1 0 16192 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _460_
timestamp 1665323087
transform -1 0 14168 0 -1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _461_
timestamp 1665323087
transform 1 0 11132 0 1 14688
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _462_
timestamp 1665323087
transform 1 0 10212 0 -1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _463_
timestamp 1665323087
transform 1 0 12328 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _464_
timestamp 1665323087
transform 1 0 12328 0 -1 14688
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _465_
timestamp 1665323087
transform 1 0 13524 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__037_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 7820 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_divider.out
timestamp 1665323087
transform 1 0 9016 0 1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_divider2.out
timestamp 1665323087
transform 1 0 12328 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_ext_clk
timestamp 1665323087
transform 1 0 5152 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_net10
timestamp 1665323087
transform 1 0 8740 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_pll_clk
timestamp 1665323087
transform -1 0 6992 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_pll_clk90
timestamp 1665323087
transform -1 0 15640 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__037_
timestamp 1665323087
transform -1 0 7084 0 -1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_divider.out
timestamp 1665323087
transform -1 0 9660 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_divider2.out
timestamp 1665323087
transform -1 0 12052 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_ext_clk
timestamp 1665323087
transform -1 0 4600 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_net10
timestamp 1665323087
transform -1 0 8188 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_pll_clk90
timestamp 1665323087
transform -1 0 14444 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_pll_clk
timestamp 1665323087
transform -1 0 4600 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__037_
timestamp 1665323087
transform 1 0 14720 0 -1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_divider.out
timestamp 1665323087
transform -1 0 9660 0 -1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_divider2.out
timestamp 1665323087
transform -1 0 12052 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_ext_clk
timestamp 1665323087
transform 1 0 4232 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_net10
timestamp 1665323087
transform 1 0 11132 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_pll_clk90
timestamp 1665323087
transform -1 0 14444 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_pll_clk
timestamp 1665323087
transform -1 0 4600 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_4  fanout13 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 15916 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout14
timestamp 1665323087
transform -1 0 16284 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout15
timestamp 1665323087
transform -1 0 15364 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 16468 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout17
timestamp 1665323087
transform -1 0 6900 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout18
timestamp 1665323087
transform 1 0 7452 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout19
timestamp 1665323087
transform -1 0 4876 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout20
timestamp 1665323087
transform -1 0 8096 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 17112 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout22
timestamp 1665323087
transform -1 0 17664 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout23
timestamp 1665323087
transform -1 0 7912 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout24
timestamp 1665323087
transform -1 0 5796 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout25
timestamp 1665323087
transform 1 0 2300 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout26
timestamp 1665323087
transform -1 0 2576 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout27
timestamp 1665323087
transform -1 0 10764 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout28
timestamp 1665323087
transform 1 0 11132 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 2760 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 18032 0 1 1632
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 17756 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1665323087
transform -1 0 2484 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1665323087
transform 1 0 18216 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1665323087
transform 1 0 17756 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1665323087
transform 1 0 18216 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1665323087
transform 1 0 18216 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1665323087
transform 1 0 18216 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1665323087
transform 1 0 18216 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  output11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 13524 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  user_clk_out_buffer
timestamp 1665323087
transform 1 0 11132 0 1 16864
box -38 -48 1878 592
<< labels >>
flabel metal4 s 3100 496 3420 18544 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 6200 496 6520 18544 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 9300 496 9620 18544 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 12400 496 12720 18544 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 15500 496 15820 18544 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 18600 496 18920 18544 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 136 3220 18920 3540 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 136 6600 18920 6920 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 136 9980 18920 10300 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 136 13360 18920 13680 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 136 16740 18920 17060 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 1550 496 1870 18544 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 4650 496 4970 18544 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 7750 496 8070 18544 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 10850 496 11170 18544 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 13950 496 14270 18544 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 17050 496 17370 18544 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 136 1530 18908 1850 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 136 4910 18908 5230 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 136 8290 18908 8610 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 136 11670 18908 11990 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 136 15050 18908 15370 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 7102 19200 7158 20000 0 FreeSans 224 90 0 0 core_clk
port 2 nsew signal tristate
flabel metal2 s 4250 19200 4306 20000 0 FreeSans 224 90 0 0 ext_clk
port 3 nsew signal input
flabel metal3 s 19200 1368 20000 1488 0 FreeSans 480 0 0 0 ext_clk_sel
port 4 nsew signal input
flabel metal3 s 19200 18504 20000 18624 0 FreeSans 480 0 0 0 ext_reset
port 5 nsew signal input
flabel metal2 s 15658 19200 15714 20000 0 FreeSans 224 90 0 0 pll_clk
port 6 nsew signal input
flabel metal2 s 18510 19200 18566 20000 0 FreeSans 224 90 0 0 pll_clk90
port 7 nsew signal input
flabel metal2 s 1398 19200 1454 20000 0 FreeSans 224 90 0 0 resetb
port 8 nsew signal input
flabel metal2 s 12806 19200 12862 20000 0 FreeSans 224 90 0 0 resetb_sync
port 9 nsew signal tristate
flabel metal3 s 19200 11160 20000 11280 0 FreeSans 480 0 0 0 sel2[0]
port 10 nsew signal input
flabel metal3 s 19200 13608 20000 13728 0 FreeSans 480 0 0 0 sel2[1]
port 11 nsew signal input
flabel metal3 s 19200 16056 20000 16176 0 FreeSans 480 0 0 0 sel2[2]
port 12 nsew signal input
flabel metal3 s 19200 3816 20000 3936 0 FreeSans 480 0 0 0 sel[0]
port 13 nsew signal input
flabel metal3 s 19200 6264 20000 6384 0 FreeSans 480 0 0 0 sel[1]
port 14 nsew signal input
flabel metal3 s 19200 8712 20000 8832 0 FreeSans 480 0 0 0 sel[2]
port 15 nsew signal input
flabel metal2 s 9954 19200 10010 20000 0 FreeSans 224 90 0 0 user_clk
port 16 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 20000 20000
<< end >>
