VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO chip_io_alt
  CLASS BLOCK ;
  FOREIGN chip_io_alt ;
  ORIGIN 0.000 0.000 ;
  SIZE 3588.000 BY 5188.000 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 938.200 32.990 1000.800 95.440 ;
    END
  END clock
  PIN clock_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.635 208.565 936.915 210.965 ;
    END
  END clock_core
  PIN por
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.215 208.565 970.495 210.965 ;
    END
  END por
  PIN flash_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1755.200 32.990 1817.800 95.440 ;
    END
  END flash_clk
  PIN flash_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1481.200 32.990 1543.800 95.440 ;
    END
  END flash_csb
  PIN flash_io0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2029.200 32.990 2091.800 95.440 ;
    END
  END flash_io0
  PIN flash_io0_di_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2027.635 208.565 2027.915 210.965 ;
    END
  END flash_io0_di_core
  PIN flash_io0_do_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2082.835 208.565 2083.115 210.965 ;
    END
  END flash_io0_do_core
  PIN flash_io0_ieb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2046.020 212.985 2077.220 213.265 ;
        RECT 2076.825 212.965 2077.165 212.985 ;
      LAYER via ;
        RECT 2046.050 212.985 2046.330 213.265 ;
        RECT 2061.215 212.985 2061.495 213.265 ;
        RECT 2076.855 212.965 2077.135 213.245 ;
      LAYER met2 ;
        RECT 2046.035 213.295 2046.315 213.360 ;
        RECT 2046.035 212.955 2046.330 213.295 ;
        RECT 2046.035 208.565 2046.315 212.955 ;
        RECT 2061.215 208.565 2061.495 213.390 ;
        RECT 2076.855 208.565 2077.135 213.335 ;
    END
  END flash_io0_ieb_core
  PIN flash_io0_oeb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2055.045 213.460 2098.785 213.740 ;
        RECT 2055.200 213.425 2055.555 213.460 ;
      LAYER via ;
        RECT 2055.230 213.425 2055.525 213.720 ;
        RECT 2098.475 213.460 2098.755 213.740 ;
      LAYER met2 ;
        RECT 2055.230 210.155 2055.525 213.750 ;
        RECT 2055.235 208.565 2055.515 210.155 ;
        RECT 2098.475 208.565 2098.755 213.770 ;
    END
  END flash_io0_oeb_core
  PIN flash_io1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2303.200 32.990 2365.800 95.440 ;
    END
  END flash_io1
  PIN flash_io1_di_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2301.635 208.565 2301.915 210.965 ;
    END
  END flash_io1_di_core
  PIN flash_io1_do_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2356.835 208.565 2357.115 210.965 ;
    END
  END flash_io1_do_core
  PIN flash_io1_ieb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2335.215 213.770 2335.495 213.800 ;
        RECT 2320.000 213.490 2351.155 213.770 ;
        RECT 2335.215 213.460 2335.495 213.490 ;
      LAYER via ;
        RECT 2320.030 213.490 2320.310 213.770 ;
        RECT 2335.215 213.490 2335.495 213.770 ;
        RECT 2350.845 213.490 2351.125 213.770 ;
      LAYER met2 ;
        RECT 2320.035 213.800 2320.315 213.840 ;
        RECT 2320.030 213.460 2320.315 213.800 ;
        RECT 2350.845 213.790 2351.125 213.800 ;
        RECT 2335.185 213.490 2335.525 213.770 ;
        RECT 2320.035 208.565 2320.315 213.460 ;
        RECT 2335.215 208.565 2335.495 213.490 ;
        RECT 2350.845 213.460 2351.135 213.790 ;
        RECT 2350.855 208.565 2351.135 213.460 ;
    END
  END flash_io1_ieb_core
  PIN flash_io1_oeb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2329.195 212.820 2372.785 213.100 ;
      LAYER via ;
        RECT 2329.225 212.820 2329.505 213.100 ;
        RECT 2372.475 212.820 2372.755 213.100 ;
      LAYER met2 ;
        RECT 2329.235 213.130 2329.515 213.170 ;
        RECT 2329.225 212.790 2329.515 213.130 ;
        RECT 2329.235 208.565 2329.515 212.790 ;
        RECT 2372.475 208.565 2372.755 213.130 ;
    END
  END flash_io1_oeb_core
  PIN gpio
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2577.200 32.990 2639.800 95.440 ;
    END
  END gpio
  PIN gpio_in_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2575.635 208.565 2575.915 210.965 ;
    END
  END gpio_in_core
  PIN gpio_inenb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2609.215 208.565 2609.495 210.965 ;
    END
  END gpio_inenb_core
  PIN gpio_mode0_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2603.235 208.565 2603.515 210.965 ;
    END
  END gpio_mode0_core
  PIN gpio_mode1_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2593.990 213.555 2594.310 213.615 ;
        RECT 2624.730 213.555 2625.050 213.615 ;
        RECT 2593.990 213.415 2625.050 213.555 ;
        RECT 2593.990 213.355 2594.310 213.415 ;
        RECT 2624.730 213.355 2625.050 213.415 ;
      LAYER via ;
        RECT 2594.020 213.355 2594.280 213.615 ;
        RECT 2624.760 213.355 2625.020 213.615 ;
      LAYER met2 ;
        RECT 2594.080 213.645 2594.220 213.735 ;
        RECT 2594.020 213.325 2594.280 213.645 ;
        RECT 2624.760 213.325 2625.020 213.645 ;
        RECT 2594.080 210.965 2594.220 213.325 ;
        RECT 2624.820 210.975 2624.960 213.325 ;
        RECT 2594.035 208.565 2594.315 210.965 ;
        RECT 2624.820 210.510 2625.135 210.975 ;
        RECT 2624.855 208.565 2625.135 210.510 ;
    END
  END gpio_mode1_core
  PIN gpio_out_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2630.835 208.565 2631.115 210.965 ;
    END
  END gpio_out_core
  PIN gpio_outenb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2646.475 208.565 2646.755 210.965 ;
    END
  END gpio_outenb_core
  PIN vccd_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 30.835 350.270 98.100 404.670 ;
    END
  END vccd_pad
  PIN vdda_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3121.110 34.055 3181.950 94.880 ;
    END
  END vdda_pad
  PIN vddio_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 34.055 558.050 94.880 618.890 ;
    END
  END vddio_pad
  PIN vddio_pad2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 34.055 4356.050 94.880 4416.890 ;
    END
  END vddio_pad2
  PIN vssa_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 401.110 34.055 461.950 94.880 ;
    END
  END vssa_pad
  PIN vssd_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1216.330 30.835 1270.730 98.100 ;
    END
  END vssd_pad
  PIN vssio_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2852.110 34.055 2912.950 94.880 ;
    END
  END vssio_pad
  PIN vssio_pad2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1674.050 5093.120 1734.890 5153.945 ;
    END
  END vssio_pad2
  PIN mprj_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 506.200 3555.010 568.800 ;
    END
  END mprj_io[0]
  PIN mprj_io_analog_en[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 529.015 3379.435 529.295 ;
    END
  END mprj_io_analog_en[0]
  PIN mprj_io_analog_pol[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 535.455 3379.435 535.735 ;
    END
  END mprj_io_analog_pol[0]
  PIN mprj_io_analog_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 550.635 3379.435 550.915 ;
    END
  END mprj_io_analog_sel[0]
  PIN mprj_io_dm[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 532.235 3379.435 532.515 ;
    END
  END mprj_io_dm[0]
  PIN mprj_io_dm[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 523.035 3379.435 523.315 ;
    END
  END mprj_io_dm[1]
  PIN mprj_io_dm[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 553.855 3379.435 554.135 ;
    END
  END mprj_io_dm[2]
  PIN mprj_io_holdover[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 557.075 3379.435 557.355 ;
    END
  END mprj_io_holdover[0]
  PIN mprj_io_ib_mode_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 572.255 3379.435 572.535 ;
    END
  END mprj_io_ib_mode_sel[0]
  PIN mprj_io_inp_dis[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 538.215 3379.435 538.495 ;
    END
  END mprj_io_inp_dis[0]
  PIN mprj_io_oeb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 575.475 3379.435 575.755 ;
    END
  END mprj_io_oeb[0]
  PIN mprj_io_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 559.835 3379.435 560.115 ;
    END
  END mprj_io_out[0]
  PIN mprj_io_slow_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 513.835 3379.435 514.115 ;
    END
  END mprj_io_slow_sel[0]
  PIN mprj_io_vtrip_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 569.035 3379.435 569.315 ;
    END
  END mprj_io_vtrip_sel[0]
  PIN mprj_io_in[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 504.635 3379.435 504.915 ;
    END
  END mprj_io_in[0]
  PIN mprj_io_in_3v3[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 578.235 3379.435 578.515 ;
    END
  END mprj_io_in_3v3[0]
  PIN mprj_gpio_analog[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3433.055 3379.435 3433.335 ;
    END
  END mprj_gpio_analog[3]
  PIN mprj_gpio_noesd[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3442.255 3379.435 3442.535 ;
    END
  END mprj_gpio_noesd[3]
  PIN mprj_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 3422.200 3555.010 3484.800 ;
    END
  END mprj_io[10]
  PIN mprj_io_analog_en[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3445.015 3379.435 3445.295 ;
    END
  END mprj_io_analog_en[10]
  PIN mprj_io_analog_pol[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3451.455 3379.435 3451.735 ;
    END
  END mprj_io_analog_pol[10]
  PIN mprj_io_analog_sel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3466.635 3379.435 3466.915 ;
    END
  END mprj_io_analog_sel[10]
  PIN mprj_io_dm[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3448.235 3379.435 3448.515 ;
    END
  END mprj_io_dm[30]
  PIN mprj_io_dm[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3439.035 3379.435 3439.315 ;
    END
  END mprj_io_dm[31]
  PIN mprj_io_dm[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3469.855 3379.435 3470.135 ;
    END
  END mprj_io_dm[32]
  PIN mprj_io_holdover[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3473.075 3379.435 3473.355 ;
    END
  END mprj_io_holdover[10]
  PIN mprj_io_ib_mode_sel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3488.255 3379.435 3488.535 ;
    END
  END mprj_io_ib_mode_sel[10]
  PIN mprj_io_inp_dis[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3454.215 3379.435 3454.495 ;
    END
  END mprj_io_inp_dis[10]
  PIN mprj_io_oeb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3491.475 3379.435 3491.755 ;
    END
  END mprj_io_oeb[10]
  PIN mprj_io_out[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3475.835 3379.435 3476.115 ;
    END
  END mprj_io_out[10]
  PIN mprj_io_slow_sel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3429.835 3379.435 3430.115 ;
    END
  END mprj_io_slow_sel[10]
  PIN mprj_io_vtrip_sel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3485.035 3379.435 3485.315 ;
    END
  END mprj_io_vtrip_sel[10]
  PIN mprj_io_in[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3420.635 3379.435 3420.915 ;
    END
  END mprj_io_in[10]
  PIN mprj_io_in_3v3[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3494.235 3379.435 3494.515 ;
    END
  END mprj_io_in_3v3[10]
  PIN mprj_gpio_analog[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3658.055 3379.435 3658.335 ;
    END
  END mprj_gpio_analog[4]
  PIN mprj_gpio_noesd[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3667.255 3379.435 3667.535 ;
    END
  END mprj_gpio_noesd[4]
  PIN mprj_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 3647.200 3555.010 3709.800 ;
    END
  END mprj_io[11]
  PIN mprj_io_analog_en[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3670.015 3379.435 3670.295 ;
    END
  END mprj_io_analog_en[11]
  PIN mprj_io_analog_pol[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3676.455 3379.435 3676.735 ;
    END
  END mprj_io_analog_pol[11]
  PIN mprj_io_analog_sel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3691.635 3379.435 3691.915 ;
    END
  END mprj_io_analog_sel[11]
  PIN mprj_io_dm[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3673.235 3379.435 3673.515 ;
    END
  END mprj_io_dm[33]
  PIN mprj_io_dm[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3664.035 3379.435 3664.315 ;
    END
  END mprj_io_dm[34]
  PIN mprj_io_dm[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3694.855 3379.435 3695.135 ;
    END
  END mprj_io_dm[35]
  PIN mprj_io_holdover[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3698.075 3379.435 3698.355 ;
    END
  END mprj_io_holdover[11]
  PIN mprj_io_ib_mode_sel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3713.255 3379.435 3713.535 ;
    END
  END mprj_io_ib_mode_sel[11]
  PIN mprj_io_inp_dis[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3679.215 3379.435 3679.495 ;
    END
  END mprj_io_inp_dis[11]
  PIN mprj_io_oeb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3716.475 3379.435 3716.755 ;
    END
  END mprj_io_oeb[11]
  PIN mprj_io_out[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3700.835 3379.435 3701.115 ;
    END
  END mprj_io_out[11]
  PIN mprj_io_slow_sel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3654.835 3379.435 3655.115 ;
    END
  END mprj_io_slow_sel[11]
  PIN mprj_io_vtrip_sel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3710.035 3379.435 3710.315 ;
    END
  END mprj_io_vtrip_sel[11]
  PIN mprj_io_in[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3645.635 3379.435 3645.915 ;
    END
  END mprj_io_in[11]
  PIN mprj_io_in_3v3[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3719.235 3379.435 3719.515 ;
    END
  END mprj_io_in_3v3[11]
  PIN mprj_gpio_analog[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3883.055 3379.435 3883.335 ;
    END
  END mprj_gpio_analog[5]
  PIN mprj_gpio_noesd[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3892.255 3379.435 3892.535 ;
    END
  END mprj_gpio_noesd[5]
  PIN mprj_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 3872.200 3555.010 3934.800 ;
    END
  END mprj_io[12]
  PIN mprj_io_analog_en[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3895.015 3379.435 3895.295 ;
    END
  END mprj_io_analog_en[12]
  PIN mprj_io_analog_pol[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3901.455 3379.435 3901.735 ;
    END
  END mprj_io_analog_pol[12]
  PIN mprj_io_analog_sel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3916.635 3379.435 3916.915 ;
    END
  END mprj_io_analog_sel[12]
  PIN mprj_io_dm[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3898.235 3379.435 3898.515 ;
    END
  END mprj_io_dm[36]
  PIN mprj_io_dm[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3889.035 3379.435 3889.315 ;
    END
  END mprj_io_dm[37]
  PIN mprj_io_dm[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3919.855 3379.435 3920.135 ;
    END
  END mprj_io_dm[38]
  PIN mprj_io_holdover[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3923.075 3379.435 3923.355 ;
    END
  END mprj_io_holdover[12]
  PIN mprj_io_ib_mode_sel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3938.255 3379.435 3938.535 ;
    END
  END mprj_io_ib_mode_sel[12]
  PIN mprj_io_inp_dis[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3904.215 3379.435 3904.495 ;
    END
  END mprj_io_inp_dis[12]
  PIN mprj_io_oeb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3941.475 3379.435 3941.755 ;
    END
  END mprj_io_oeb[12]
  PIN mprj_io_out[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3925.835 3379.435 3926.115 ;
    END
  END mprj_io_out[12]
  PIN mprj_io_slow_sel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3879.835 3379.435 3880.115 ;
    END
  END mprj_io_slow_sel[12]
  PIN mprj_io_vtrip_sel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3935.035 3379.435 3935.315 ;
    END
  END mprj_io_vtrip_sel[12]
  PIN mprj_io_in[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3870.635 3379.435 3870.915 ;
    END
  END mprj_io_in[12]
  PIN mprj_io_in_3v3[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3944.235 3379.435 3944.515 ;
    END
  END mprj_io_in_3v3[12]
  PIN mprj_gpio_analog[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4329.055 3379.435 4329.335 ;
    END
  END mprj_gpio_analog[6]
  PIN mprj_gpio_noesd[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4338.255 3379.435 4338.535 ;
    END
  END mprj_gpio_noesd[6]
  PIN mprj_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 4318.200 3555.010 4380.800 ;
    END
  END mprj_io[13]
  PIN mprj_io_analog_en[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4341.015 3379.435 4341.295 ;
    END
  END mprj_io_analog_en[13]
  PIN mprj_io_analog_pol[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4347.455 3379.435 4347.735 ;
    END
  END mprj_io_analog_pol[13]
  PIN mprj_io_analog_sel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4362.635 3379.435 4362.915 ;
    END
  END mprj_io_analog_sel[13]
  PIN mprj_io_dm[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4344.235 3379.435 4344.515 ;
    END
  END mprj_io_dm[39]
  PIN mprj_io_dm[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4335.035 3379.435 4335.315 ;
    END
  END mprj_io_dm[40]
  PIN mprj_io_dm[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4365.855 3379.435 4366.135 ;
    END
  END mprj_io_dm[41]
  PIN mprj_io_holdover[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4369.075 3379.435 4369.355 ;
    END
  END mprj_io_holdover[13]
  PIN mprj_io_ib_mode_sel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4384.255 3379.435 4384.535 ;
    END
  END mprj_io_ib_mode_sel[13]
  PIN mprj_io_inp_dis[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4350.215 3379.435 4350.495 ;
    END
  END mprj_io_inp_dis[13]
  PIN mprj_io_oeb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4387.475 3379.435 4387.755 ;
    END
  END mprj_io_oeb[13]
  PIN mprj_io_out[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4371.835 3379.435 4372.115 ;
    END
  END mprj_io_out[13]
  PIN mprj_io_slow_sel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4325.835 3379.435 4326.115 ;
    END
  END mprj_io_slow_sel[13]
  PIN mprj_io_vtrip_sel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4381.035 3379.435 4381.315 ;
    END
  END mprj_io_vtrip_sel[13]
  PIN mprj_io_in[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4316.635 3379.435 4316.915 ;
    END
  END mprj_io_in[13]
  PIN mprj_io_in_3v3[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4390.235 3379.435 4390.515 ;
    END
  END mprj_io_in_3v3[13]
  PIN mprj_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 732.200 3555.010 794.800 ;
    END
  END mprj_io[1]
  PIN mprj_io_analog_en[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 755.015 3379.435 755.295 ;
    END
  END mprj_io_analog_en[1]
  PIN mprj_io_analog_pol[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 761.455 3379.435 761.735 ;
    END
  END mprj_io_analog_pol[1]
  PIN mprj_io_analog_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 776.635 3379.435 776.915 ;
    END
  END mprj_io_analog_sel[1]
  PIN mprj_io_dm[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 758.235 3379.435 758.515 ;
    END
  END mprj_io_dm[3]
  PIN mprj_io_dm[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 749.035 3379.435 749.315 ;
    END
  END mprj_io_dm[4]
  PIN mprj_io_dm[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 779.855 3379.435 780.135 ;
    END
  END mprj_io_dm[5]
  PIN mprj_io_holdover[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 783.075 3379.435 783.355 ;
    END
  END mprj_io_holdover[1]
  PIN mprj_io_ib_mode_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 798.255 3379.435 798.535 ;
    END
  END mprj_io_ib_mode_sel[1]
  PIN mprj_io_inp_dis[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 764.215 3379.435 764.495 ;
    END
  END mprj_io_inp_dis[1]
  PIN mprj_io_oeb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 801.475 3379.435 801.755 ;
    END
  END mprj_io_oeb[1]
  PIN mprj_io_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 785.835 3379.435 786.115 ;
    END
  END mprj_io_out[1]
  PIN mprj_io_slow_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 739.835 3379.435 740.115 ;
    END
  END mprj_io_slow_sel[1]
  PIN mprj_io_vtrip_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 795.035 3379.435 795.315 ;
    END
  END mprj_io_vtrip_sel[1]
  PIN mprj_io_in[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 730.635 3379.435 730.915 ;
    END
  END mprj_io_in[1]
  PIN mprj_io_in_3v3[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 804.235 3379.435 804.515 ;
    END
  END mprj_io_in_3v3[1]
  PIN mprj_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 957.200 3555.010 1019.800 ;
    END
  END mprj_io[2]
  PIN mprj_io_analog_en[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 980.015 3379.435 980.295 ;
    END
  END mprj_io_analog_en[2]
  PIN mprj_io_analog_pol[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 986.455 3379.435 986.735 ;
    END
  END mprj_io_analog_pol[2]
  PIN mprj_io_analog_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1001.635 3379.435 1001.915 ;
    END
  END mprj_io_analog_sel[2]
  PIN mprj_io_dm[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 983.235 3379.435 983.515 ;
    END
  END mprj_io_dm[6]
  PIN mprj_io_dm[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 974.035 3379.435 974.315 ;
    END
  END mprj_io_dm[7]
  PIN mprj_io_dm[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1004.855 3379.435 1005.135 ;
    END
  END mprj_io_dm[8]
  PIN mprj_io_holdover[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1008.075 3379.435 1008.355 ;
    END
  END mprj_io_holdover[2]
  PIN mprj_io_ib_mode_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1023.255 3379.435 1023.535 ;
    END
  END mprj_io_ib_mode_sel[2]
  PIN mprj_io_inp_dis[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 989.215 3379.435 989.495 ;
    END
  END mprj_io_inp_dis[2]
  PIN mprj_io_oeb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1026.475 3379.435 1026.755 ;
    END
  END mprj_io_oeb[2]
  PIN mprj_io_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1010.835 3379.435 1011.115 ;
    END
  END mprj_io_out[2]
  PIN mprj_io_slow_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 964.835 3379.435 965.115 ;
    END
  END mprj_io_slow_sel[2]
  PIN mprj_io_vtrip_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1020.035 3379.435 1020.315 ;
    END
  END mprj_io_vtrip_sel[2]
  PIN mprj_io_in[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 955.635 3379.435 955.915 ;
    END
  END mprj_io_in[2]
  PIN mprj_io_in_3v3[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1029.235 3379.435 1029.515 ;
    END
  END mprj_io_in_3v3[2]
  PIN mprj_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 1183.200 3555.010 1245.800 ;
    END
  END mprj_io[3]
  PIN mprj_io_analog_en[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1206.015 3379.435 1206.295 ;
    END
  END mprj_io_analog_en[3]
  PIN mprj_io_analog_pol[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1212.455 3379.435 1212.735 ;
    END
  END mprj_io_analog_pol[3]
  PIN mprj_io_analog_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1227.635 3379.435 1227.915 ;
    END
  END mprj_io_analog_sel[3]
  PIN mprj_io_dm[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1200.035 3379.435 1200.315 ;
    END
  END mprj_io_dm[10]
  PIN mprj_io_dm[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1230.855 3379.435 1231.135 ;
    END
  END mprj_io_dm[11]
  PIN mprj_io_dm[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1209.235 3379.435 1209.515 ;
    END
  END mprj_io_dm[9]
  PIN mprj_io_holdover[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1234.075 3379.435 1234.355 ;
    END
  END mprj_io_holdover[3]
  PIN mprj_io_ib_mode_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1249.255 3379.435 1249.535 ;
    END
  END mprj_io_ib_mode_sel[3]
  PIN mprj_io_inp_dis[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1215.215 3379.435 1215.495 ;
    END
  END mprj_io_inp_dis[3]
  PIN mprj_io_oeb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1252.475 3379.435 1252.755 ;
    END
  END mprj_io_oeb[3]
  PIN mprj_io_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1236.835 3379.435 1237.115 ;
    END
  END mprj_io_out[3]
  PIN mprj_io_slow_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1190.835 3379.435 1191.115 ;
    END
  END mprj_io_slow_sel[3]
  PIN mprj_io_vtrip_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1246.035 3379.435 1246.315 ;
    END
  END mprj_io_vtrip_sel[3]
  PIN mprj_io_in[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1181.635 3379.435 1181.915 ;
    END
  END mprj_io_in[3]
  PIN mprj_io_in_3v3[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1255.235 3379.435 1255.515 ;
    END
  END mprj_io_in_3v3[3]
  PIN mprj_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 1408.200 3555.010 1470.800 ;
    END
  END mprj_io[4]
  PIN mprj_io_analog_en[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1431.015 3379.435 1431.295 ;
    END
  END mprj_io_analog_en[4]
  PIN mprj_io_analog_pol[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1437.455 3379.435 1437.735 ;
    END
  END mprj_io_analog_pol[4]
  PIN mprj_io_analog_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1452.635 3379.435 1452.915 ;
    END
  END mprj_io_analog_sel[4]
  PIN mprj_io_dm[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1434.235 3379.435 1434.515 ;
    END
  END mprj_io_dm[12]
  PIN mprj_io_dm[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1425.035 3379.435 1425.315 ;
    END
  END mprj_io_dm[13]
  PIN mprj_io_dm[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1455.855 3379.435 1456.135 ;
    END
  END mprj_io_dm[14]
  PIN mprj_io_holdover[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1459.075 3379.435 1459.355 ;
    END
  END mprj_io_holdover[4]
  PIN mprj_io_ib_mode_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1474.255 3379.435 1474.535 ;
    END
  END mprj_io_ib_mode_sel[4]
  PIN mprj_io_inp_dis[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1440.215 3379.435 1440.495 ;
    END
  END mprj_io_inp_dis[4]
  PIN mprj_io_oeb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1477.475 3379.435 1477.755 ;
    END
  END mprj_io_oeb[4]
  PIN mprj_io_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1461.835 3379.435 1462.115 ;
    END
  END mprj_io_out[4]
  PIN mprj_io_slow_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1415.835 3379.435 1416.115 ;
    END
  END mprj_io_slow_sel[4]
  PIN mprj_io_vtrip_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1471.035 3379.435 1471.315 ;
    END
  END mprj_io_vtrip_sel[4]
  PIN mprj_io_in[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1406.635 3379.435 1406.915 ;
    END
  END mprj_io_in[4]
  PIN mprj_io_in_3v3[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1480.235 3379.435 1480.515 ;
    END
  END mprj_io_in_3v3[4]
  PIN mprj_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 1633.200 3555.010 1695.800 ;
    END
  END mprj_io[5]
  PIN mprj_io_analog_en[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1656.015 3379.435 1656.295 ;
    END
  END mprj_io_analog_en[5]
  PIN mprj_io_analog_pol[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1662.455 3379.435 1662.735 ;
    END
  END mprj_io_analog_pol[5]
  PIN mprj_io_analog_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1677.635 3379.435 1677.915 ;
    END
  END mprj_io_analog_sel[5]
  PIN mprj_io_dm[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1659.235 3379.435 1659.515 ;
    END
  END mprj_io_dm[15]
  PIN mprj_io_dm[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1650.035 3379.435 1650.315 ;
    END
  END mprj_io_dm[16]
  PIN mprj_io_dm[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1680.855 3379.435 1681.135 ;
    END
  END mprj_io_dm[17]
  PIN mprj_io_holdover[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1684.075 3379.435 1684.355 ;
    END
  END mprj_io_holdover[5]
  PIN mprj_io_ib_mode_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1699.255 3379.435 1699.535 ;
    END
  END mprj_io_ib_mode_sel[5]
  PIN mprj_io_inp_dis[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1665.215 3379.435 1665.495 ;
    END
  END mprj_io_inp_dis[5]
  PIN mprj_io_oeb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1702.475 3379.435 1702.755 ;
    END
  END mprj_io_oeb[5]
  PIN mprj_io_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1686.835 3379.435 1687.115 ;
    END
  END mprj_io_out[5]
  PIN mprj_io_slow_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1640.835 3379.435 1641.115 ;
    END
  END mprj_io_slow_sel[5]
  PIN mprj_io_vtrip_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1696.035 3379.435 1696.315 ;
    END
  END mprj_io_vtrip_sel[5]
  PIN mprj_io_in[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1631.635 3379.435 1631.915 ;
    END
  END mprj_io_in[5]
  PIN mprj_io_in_3v3[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1705.235 3379.435 1705.515 ;
    END
  END mprj_io_in_3v3[5]
  PIN mprj_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 1859.200 3555.010 1921.800 ;
    END
  END mprj_io[6]
  PIN mprj_io_analog_en[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1882.015 3379.435 1882.295 ;
    END
  END mprj_io_analog_en[6]
  PIN mprj_io_analog_pol[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1888.455 3379.435 1888.735 ;
    END
  END mprj_io_analog_pol[6]
  PIN mprj_io_analog_sel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1903.635 3379.435 1903.915 ;
    END
  END mprj_io_analog_sel[6]
  PIN mprj_io_dm[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1885.235 3379.435 1885.515 ;
    END
  END mprj_io_dm[18]
  PIN mprj_io_dm[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1876.035 3379.435 1876.315 ;
    END
  END mprj_io_dm[19]
  PIN mprj_io_dm[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1906.855 3379.435 1907.135 ;
    END
  END mprj_io_dm[20]
  PIN mprj_io_holdover[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1910.075 3379.435 1910.355 ;
    END
  END mprj_io_holdover[6]
  PIN mprj_io_ib_mode_sel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1925.255 3379.435 1925.535 ;
    END
  END mprj_io_ib_mode_sel[6]
  PIN mprj_io_inp_dis[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1891.215 3379.435 1891.495 ;
    END
  END mprj_io_inp_dis[6]
  PIN mprj_io_oeb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1928.475 3379.435 1928.755 ;
    END
  END mprj_io_oeb[6]
  PIN mprj_io_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1912.835 3379.435 1913.115 ;
    END
  END mprj_io_out[6]
  PIN mprj_io_slow_sel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1866.835 3379.435 1867.115 ;
    END
  END mprj_io_slow_sel[6]
  PIN mprj_io_vtrip_sel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1922.035 3379.435 1922.315 ;
    END
  END mprj_io_vtrip_sel[6]
  PIN mprj_io_in[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1857.635 3379.435 1857.915 ;
    END
  END mprj_io_in[6]
  PIN mprj_io_in_3v3[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1931.235 3379.435 1931.515 ;
    END
  END mprj_io_in_3v3[6]
  PIN mprj_gpio_analog[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2756.055 3379.435 2756.335 ;
    END
  END mprj_gpio_analog[0]
  PIN mprj_gpio_noesd[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2765.255 3379.435 2765.535 ;
    END
  END mprj_gpio_noesd[0]
  PIN mprj_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 2745.200 3555.010 2807.800 ;
    END
  END mprj_io[7]
  PIN mprj_io_analog_en[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2768.015 3379.435 2768.295 ;
    END
  END mprj_io_analog_en[7]
  PIN mprj_io_analog_pol[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2774.455 3379.435 2774.735 ;
    END
  END mprj_io_analog_pol[7]
  PIN mprj_io_analog_sel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2789.635 3379.435 2789.915 ;
    END
  END mprj_io_analog_sel[7]
  PIN mprj_io_dm[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2771.235 3379.435 2771.515 ;
    END
  END mprj_io_dm[21]
  PIN mprj_io_dm[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2762.035 3379.435 2762.315 ;
    END
  END mprj_io_dm[22]
  PIN mprj_io_dm[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2792.855 3379.435 2793.135 ;
    END
  END mprj_io_dm[23]
  PIN mprj_io_holdover[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2796.075 3379.435 2796.355 ;
    END
  END mprj_io_holdover[7]
  PIN mprj_io_ib_mode_sel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2811.255 3379.435 2811.535 ;
    END
  END mprj_io_ib_mode_sel[7]
  PIN mprj_io_inp_dis[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2777.215 3379.435 2777.495 ;
    END
  END mprj_io_inp_dis[7]
  PIN mprj_io_oeb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2814.475 3379.435 2814.755 ;
    END
  END mprj_io_oeb[7]
  PIN mprj_io_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2798.835 3379.435 2799.115 ;
    END
  END mprj_io_out[7]
  PIN mprj_io_slow_sel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2752.835 3379.435 2753.115 ;
    END
  END mprj_io_slow_sel[7]
  PIN mprj_io_vtrip_sel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2808.035 3379.435 2808.315 ;
    END
  END mprj_io_vtrip_sel[7]
  PIN mprj_io_in[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2743.635 3379.435 2743.915 ;
    END
  END mprj_io_in[7]
  PIN mprj_io_in_3v3[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2817.235 3379.435 2817.515 ;
    END
  END mprj_io_in_3v3[7]
  PIN mprj_gpio_analog[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2982.055 3379.435 2982.335 ;
    END
  END mprj_gpio_analog[1]
  PIN mprj_gpio_noesd[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2991.255 3379.435 2991.535 ;
    END
  END mprj_gpio_noesd[1]
  PIN mprj_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 2971.200 3555.010 3033.800 ;
    END
  END mprj_io[8]
  PIN mprj_io_analog_en[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2994.015 3379.435 2994.295 ;
    END
  END mprj_io_analog_en[8]
  PIN mprj_io_analog_pol[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3000.455 3379.435 3000.735 ;
    END
  END mprj_io_analog_pol[8]
  PIN mprj_io_analog_sel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3015.635 3379.435 3015.915 ;
    END
  END mprj_io_analog_sel[8]
  PIN mprj_io_dm[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2997.235 3379.435 2997.515 ;
    END
  END mprj_io_dm[24]
  PIN mprj_io_dm[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2988.035 3379.435 2988.315 ;
    END
  END mprj_io_dm[25]
  PIN mprj_io_dm[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3018.855 3379.435 3019.135 ;
    END
  END mprj_io_dm[26]
  PIN mprj_io_holdover[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3022.075 3379.435 3022.355 ;
    END
  END mprj_io_holdover[8]
  PIN mprj_io_ib_mode_sel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3037.255 3379.435 3037.535 ;
    END
  END mprj_io_ib_mode_sel[8]
  PIN mprj_io_inp_dis[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3003.215 3379.435 3003.495 ;
    END
  END mprj_io_inp_dis[8]
  PIN mprj_io_oeb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3040.475 3379.435 3040.755 ;
    END
  END mprj_io_oeb[8]
  PIN mprj_io_out[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3024.835 3379.435 3025.115 ;
    END
  END mprj_io_out[8]
  PIN mprj_io_slow_sel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2978.835 3379.435 2979.115 ;
    END
  END mprj_io_slow_sel[8]
  PIN mprj_io_vtrip_sel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3034.035 3379.435 3034.315 ;
    END
  END mprj_io_vtrip_sel[8]
  PIN mprj_io_in[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2969.635 3379.435 2969.915 ;
    END
  END mprj_io_in[8]
  PIN mprj_io_in_3v3[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3043.235 3379.435 3043.515 ;
    END
  END mprj_io_in_3v3[8]
  PIN mprj_gpio_analog[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3207.055 3379.435 3207.335 ;
    END
  END mprj_gpio_analog[2]
  PIN mprj_gpio_noesd[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3216.255 3379.435 3216.535 ;
    END
  END mprj_gpio_noesd[2]
  PIN mprj_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 3196.200 3555.010 3258.800 ;
    END
  END mprj_io[9]
  PIN mprj_io_analog_en[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3219.015 3379.435 3219.295 ;
    END
  END mprj_io_analog_en[9]
  PIN mprj_io_analog_pol[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3225.455 3379.435 3225.735 ;
    END
  END mprj_io_analog_pol[9]
  PIN mprj_io_analog_sel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3240.635 3379.435 3240.915 ;
    END
  END mprj_io_analog_sel[9]
  PIN mprj_io_dm[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3222.235 3379.435 3222.515 ;
    END
  END mprj_io_dm[27]
  PIN mprj_io_dm[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3213.035 3379.435 3213.315 ;
    END
  END mprj_io_dm[28]
  PIN mprj_io_dm[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3243.855 3379.435 3244.135 ;
    END
  END mprj_io_dm[29]
  PIN mprj_io_holdover[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3247.075 3379.435 3247.355 ;
    END
  END mprj_io_holdover[9]
  PIN mprj_io_ib_mode_sel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3262.255 3379.435 3262.535 ;
    END
  END mprj_io_ib_mode_sel[9]
  PIN mprj_io_inp_dis[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3228.215 3379.435 3228.495 ;
    END
  END mprj_io_inp_dis[9]
  PIN mprj_io_oeb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3265.475 3379.435 3265.755 ;
    END
  END mprj_io_oeb[9]
  PIN mprj_io_out[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3249.835 3379.435 3250.115 ;
    END
  END mprj_io_out[9]
  PIN mprj_io_slow_sel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3203.835 3379.435 3204.115 ;
    END
  END mprj_io_slow_sel[9]
  PIN mprj_io_vtrip_sel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3259.035 3379.435 3259.315 ;
    END
  END mprj_io_vtrip_sel[9]
  PIN mprj_io_in[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3194.635 3379.435 3194.915 ;
    END
  END mprj_io_in[9]
  PIN mprj_io_in_3v3[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3268.235 3379.435 3268.515 ;
    END
  END mprj_io_in_3v3[9]
  PIN mprj_gpio_analog[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3984.665 210.965 3984.945 ;
    END
  END mprj_gpio_analog[7]
  PIN mprj_gpio_noesd[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3975.465 210.965 3975.745 ;
    END
  END mprj_gpio_noesd[7]
  PIN mprj_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 3933.200 95.440 3995.800 ;
    END
  END mprj_io[25]
  PIN mprj_io_analog_en[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3972.705 210.965 3972.985 ;
    END
  END mprj_io_analog_en[14]
  PIN mprj_io_analog_pol[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3966.265 210.965 3966.545 ;
    END
  END mprj_io_analog_pol[14]
  PIN mprj_io_analog_sel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3951.085 210.965 3951.365 ;
    END
  END mprj_io_analog_sel[14]
  PIN mprj_io_dm[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3969.485 210.965 3969.765 ;
    END
  END mprj_io_dm[42]
  PIN mprj_io_dm[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3978.685 210.965 3978.965 ;
    END
  END mprj_io_dm[43]
  PIN mprj_io_dm[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3947.865 210.965 3948.145 ;
    END
  END mprj_io_dm[44]
  PIN mprj_io_holdover[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3944.645 210.965 3944.925 ;
    END
  END mprj_io_holdover[14]
  PIN mprj_io_ib_mode_sel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3929.465 210.965 3929.745 ;
    END
  END mprj_io_ib_mode_sel[14]
  PIN mprj_io_inp_dis[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3963.505 210.965 3963.785 ;
    END
  END mprj_io_inp_dis[14]
  PIN mprj_io_oeb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3926.245 210.965 3926.525 ;
    END
  END mprj_io_oeb[14]
  PIN mprj_io_out[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3941.885 210.965 3942.165 ;
    END
  END mprj_io_out[14]
  PIN mprj_io_slow_sel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3987.885 210.965 3988.165 ;
    END
  END mprj_io_slow_sel[14]
  PIN mprj_io_vtrip_sel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3932.685 210.965 3932.965 ;
    END
  END mprj_io_vtrip_sel[14]
  PIN mprj_io_in[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3997.085 210.965 3997.365 ;
    END
  END mprj_io_in[14]
  PIN mprj_io_in_3v3[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3923.485 210.965 3923.765 ;
    END
  END mprj_io_in_3v3[14]
  PIN mprj_gpio_analog[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1402.665 210.965 1402.945 ;
    END
  END mprj_gpio_analog[17]
  PIN mprj_gpio_noesd[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1393.465 210.965 1393.745 ;
    END
  END mprj_gpio_noesd[17]
  PIN mprj_io[35]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 1351.200 95.440 1413.800 ;
    END
  END mprj_io[35]
  PIN mprj_io_analog_en[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1390.705 210.965 1390.985 ;
    END
  END mprj_io_analog_en[24]
  PIN mprj_io_analog_pol[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1384.265 210.965 1384.545 ;
    END
  END mprj_io_analog_pol[24]
  PIN mprj_io_analog_sel[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1369.085 210.965 1369.365 ;
    END
  END mprj_io_analog_sel[24]
  PIN mprj_io_dm[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1387.485 210.965 1387.765 ;
    END
  END mprj_io_dm[72]
  PIN mprj_io_dm[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1396.685 210.965 1396.965 ;
    END
  END mprj_io_dm[73]
  PIN mprj_io_dm[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1365.865 210.965 1366.145 ;
    END
  END mprj_io_dm[74]
  PIN mprj_io_holdover[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1362.645 210.965 1362.925 ;
    END
  END mprj_io_holdover[24]
  PIN mprj_io_ib_mode_sel[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1347.465 210.965 1347.745 ;
    END
  END mprj_io_ib_mode_sel[24]
  PIN mprj_io_inp_dis[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1381.505 210.965 1381.785 ;
    END
  END mprj_io_inp_dis[24]
  PIN mprj_io_oeb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1344.245 210.965 1344.525 ;
    END
  END mprj_io_oeb[24]
  PIN mprj_io_out[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1359.885 210.965 1360.165 ;
    END
  END mprj_io_out[24]
  PIN mprj_io_slow_sel[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1405.885 210.965 1406.165 ;
    END
  END mprj_io_slow_sel[24]
  PIN mprj_io_vtrip_sel[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1350.685 210.965 1350.965 ;
    END
  END mprj_io_vtrip_sel[24]
  PIN mprj_io_in[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1415.085 210.965 1415.365 ;
    END
  END mprj_io_in[24]
  PIN mprj_io_in_3v3[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1341.485 210.965 1341.765 ;
    END
  END mprj_io_in_3v3[24]
  PIN mprj_io[36]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 1135.200 95.440 1197.800 ;
    END
  END mprj_io[36]
  PIN mprj_io_analog_en[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1174.705 210.965 1174.985 ;
    END
  END mprj_io_analog_en[25]
  PIN mprj_io_analog_pol[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1168.265 210.965 1168.545 ;
    END
  END mprj_io_analog_pol[25]
  PIN mprj_io_analog_sel[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1153.085 210.965 1153.365 ;
    END
  END mprj_io_analog_sel[25]
  PIN mprj_io_dm[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1171.485 210.965 1171.765 ;
    END
  END mprj_io_dm[75]
  PIN mprj_io_dm[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1180.685 210.965 1180.965 ;
    END
  END mprj_io_dm[76]
  PIN mprj_io_dm[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1149.865 210.965 1150.145 ;
    END
  END mprj_io_dm[77]
  PIN mprj_io_holdover[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1146.645 210.965 1146.925 ;
    END
  END mprj_io_holdover[25]
  PIN mprj_io_ib_mode_sel[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1131.465 210.965 1131.745 ;
    END
  END mprj_io_ib_mode_sel[25]
  PIN mprj_io_inp_dis[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1165.505 210.965 1165.785 ;
    END
  END mprj_io_inp_dis[25]
  PIN mprj_io_oeb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1128.245 210.965 1128.525 ;
    END
  END mprj_io_oeb[25]
  PIN mprj_io_out[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1143.885 210.965 1144.165 ;
    END
  END mprj_io_out[25]
  PIN mprj_io_slow_sel[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1189.885 210.965 1190.165 ;
    END
  END mprj_io_slow_sel[25]
  PIN mprj_io_vtrip_sel[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1134.685 210.965 1134.965 ;
    END
  END mprj_io_vtrip_sel[25]
  PIN mprj_io_in[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1199.085 210.965 1199.365 ;
    END
  END mprj_io_in[25]
  PIN mprj_io_in_3v3[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1125.485 210.965 1125.765 ;
    END
  END mprj_io_in_3v3[25]
  PIN mprj_io[37]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 919.200 95.440 981.800 ;
    END
  END mprj_io[37]
  PIN mprj_io_analog_en[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 958.705 210.965 958.985 ;
    END
  END mprj_io_analog_en[26]
  PIN mprj_io_analog_pol[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 952.265 210.965 952.545 ;
    END
  END mprj_io_analog_pol[26]
  PIN mprj_io_analog_sel[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 937.085 210.965 937.365 ;
    END
  END mprj_io_analog_sel[26]
  PIN mprj_io_dm[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 955.485 210.965 955.765 ;
    END
  END mprj_io_dm[78]
  PIN mprj_io_dm[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 964.685 210.965 964.965 ;
    END
  END mprj_io_dm[79]
  PIN mprj_io_dm[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 933.865 210.965 934.145 ;
    END
  END mprj_io_dm[80]
  PIN mprj_io_holdover[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 930.645 210.965 930.925 ;
    END
  END mprj_io_holdover[26]
  PIN mprj_io_ib_mode_sel[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 915.465 210.965 915.745 ;
    END
  END mprj_io_ib_mode_sel[26]
  PIN mprj_io_inp_dis[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 949.505 210.965 949.785 ;
    END
  END mprj_io_inp_dis[26]
  PIN mprj_io_oeb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 912.245 210.965 912.525 ;
    END
  END mprj_io_oeb[26]
  PIN mprj_io_out[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 927.885 210.965 928.165 ;
    END
  END mprj_io_out[26]
  PIN mprj_io_slow_sel[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 973.885 210.965 974.165 ;
    END
  END mprj_io_slow_sel[26]
  PIN mprj_io_vtrip_sel[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 918.685 210.965 918.965 ;
    END
  END mprj_io_vtrip_sel[26]
  PIN mprj_io_in[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 983.085 210.965 983.365 ;
    END
  END mprj_io_in[26]
  PIN mprj_io_in_3v3[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 909.485 210.965 909.765 ;
    END
  END mprj_io_in_3v3[26]
  PIN mprj_gpio_analog[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3768.665 210.965 3768.945 ;
    END
  END mprj_gpio_analog[8]
  PIN mprj_gpio_noesd[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3759.465 210.965 3759.745 ;
    END
  END mprj_gpio_noesd[8]
  PIN mprj_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 3717.200 95.440 3779.800 ;
    END
  END mprj_io[26]
  PIN mprj_io_analog_en[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3756.705 210.965 3756.985 ;
    END
  END mprj_io_analog_en[15]
  PIN mprj_io_analog_pol[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3750.265 210.965 3750.545 ;
    END
  END mprj_io_analog_pol[15]
  PIN mprj_io_analog_sel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3735.085 210.965 3735.365 ;
    END
  END mprj_io_analog_sel[15]
  PIN mprj_io_dm[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3753.485 210.965 3753.765 ;
    END
  END mprj_io_dm[45]
  PIN mprj_io_dm[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3762.685 210.965 3762.965 ;
    END
  END mprj_io_dm[46]
  PIN mprj_io_dm[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3731.865 210.965 3732.145 ;
    END
  END mprj_io_dm[47]
  PIN mprj_io_holdover[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3728.645 210.965 3728.925 ;
    END
  END mprj_io_holdover[15]
  PIN mprj_io_ib_mode_sel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3713.465 210.965 3713.745 ;
    END
  END mprj_io_ib_mode_sel[15]
  PIN mprj_io_inp_dis[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3747.505 210.965 3747.785 ;
    END
  END mprj_io_inp_dis[15]
  PIN mprj_io_oeb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3710.245 210.965 3710.525 ;
    END
  END mprj_io_oeb[15]
  PIN mprj_io_out[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3725.885 210.965 3726.165 ;
    END
  END mprj_io_out[15]
  PIN mprj_io_slow_sel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3771.885 210.965 3772.165 ;
    END
  END mprj_io_slow_sel[15]
  PIN mprj_io_vtrip_sel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3716.685 210.965 3716.965 ;
    END
  END mprj_io_vtrip_sel[15]
  PIN mprj_io_in[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3781.085 210.965 3781.365 ;
    END
  END mprj_io_in[15]
  PIN mprj_io_in_3v3[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3707.485 210.965 3707.765 ;
    END
  END mprj_io_in_3v3[15]
  PIN mprj_gpio_analog[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3552.665 210.965 3552.945 ;
    END
  END mprj_gpio_analog[9]
  PIN mprj_gpio_noesd[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3543.465 210.965 3543.745 ;
    END
  END mprj_gpio_noesd[9]
  PIN mprj_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 3501.200 95.440 3563.800 ;
    END
  END mprj_io[27]
  PIN mprj_io_analog_en[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3540.705 210.965 3540.985 ;
    END
  END mprj_io_analog_en[16]
  PIN mprj_io_analog_pol[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3534.265 210.965 3534.545 ;
    END
  END mprj_io_analog_pol[16]
  PIN mprj_io_analog_sel[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3519.085 210.965 3519.365 ;
    END
  END mprj_io_analog_sel[16]
  PIN mprj_io_dm[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3537.485 210.965 3537.765 ;
    END
  END mprj_io_dm[48]
  PIN mprj_io_dm[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3546.685 210.965 3546.965 ;
    END
  END mprj_io_dm[49]
  PIN mprj_io_dm[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3515.865 210.965 3516.145 ;
    END
  END mprj_io_dm[50]
  PIN mprj_io_holdover[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3512.645 210.965 3512.925 ;
    END
  END mprj_io_holdover[16]
  PIN mprj_io_ib_mode_sel[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3497.465 210.965 3497.745 ;
    END
  END mprj_io_ib_mode_sel[16]
  PIN mprj_io_inp_dis[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3531.505 210.965 3531.785 ;
    END
  END mprj_io_inp_dis[16]
  PIN mprj_io_oeb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3494.245 210.965 3494.525 ;
    END
  END mprj_io_oeb[16]
  PIN mprj_io_out[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3509.885 210.965 3510.165 ;
    END
  END mprj_io_out[16]
  PIN mprj_io_slow_sel[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3555.885 210.965 3556.165 ;
    END
  END mprj_io_slow_sel[16]
  PIN mprj_io_vtrip_sel[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3500.685 210.965 3500.965 ;
    END
  END mprj_io_vtrip_sel[16]
  PIN mprj_io_in[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3565.085 210.965 3565.365 ;
    END
  END mprj_io_in[16]
  PIN mprj_io_in_3v3[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3491.485 210.965 3491.765 ;
    END
  END mprj_io_in_3v3[16]
  PIN mprj_gpio_analog[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3336.665 210.965 3336.945 ;
    END
  END mprj_gpio_analog[10]
  PIN mprj_gpio_noesd[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3327.465 210.965 3327.745 ;
    END
  END mprj_gpio_noesd[10]
  PIN mprj_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 3285.200 95.440 3347.800 ;
    END
  END mprj_io[28]
  PIN mprj_io_analog_en[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3324.705 210.965 3324.985 ;
    END
  END mprj_io_analog_en[17]
  PIN mprj_io_analog_pol[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3318.265 210.965 3318.545 ;
    END
  END mprj_io_analog_pol[17]
  PIN mprj_io_analog_sel[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3303.085 210.965 3303.365 ;
    END
  END mprj_io_analog_sel[17]
  PIN mprj_io_dm[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3321.485 210.965 3321.765 ;
    END
  END mprj_io_dm[51]
  PIN mprj_io_dm[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3330.685 210.965 3330.965 ;
    END
  END mprj_io_dm[52]
  PIN mprj_io_dm[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3299.865 210.965 3300.145 ;
    END
  END mprj_io_dm[53]
  PIN mprj_io_holdover[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3296.645 210.965 3296.925 ;
    END
  END mprj_io_holdover[17]
  PIN mprj_io_ib_mode_sel[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3281.465 210.965 3281.745 ;
    END
  END mprj_io_ib_mode_sel[17]
  PIN mprj_io_inp_dis[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3315.505 210.965 3315.785 ;
    END
  END mprj_io_inp_dis[17]
  PIN mprj_io_oeb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3278.245 210.965 3278.525 ;
    END
  END mprj_io_oeb[17]
  PIN mprj_io_out[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3293.885 210.965 3294.165 ;
    END
  END mprj_io_out[17]
  PIN mprj_io_slow_sel[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3339.885 210.965 3340.165 ;
    END
  END mprj_io_slow_sel[17]
  PIN mprj_io_vtrip_sel[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3284.685 210.965 3284.965 ;
    END
  END mprj_io_vtrip_sel[17]
  PIN mprj_io_in[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3349.085 210.965 3349.365 ;
    END
  END mprj_io_in[17]
  PIN mprj_io_in_3v3[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3275.485 210.965 3275.765 ;
    END
  END mprj_io_in_3v3[17]
  PIN mprj_gpio_analog[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3120.665 210.965 3120.945 ;
    END
  END mprj_gpio_analog[11]
  PIN mprj_gpio_noesd[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3111.465 210.965 3111.745 ;
    END
  END mprj_gpio_noesd[11]
  PIN mprj_io[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 3069.200 95.440 3131.800 ;
    END
  END mprj_io[29]
  PIN mprj_io_analog_en[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3108.705 210.965 3108.985 ;
    END
  END mprj_io_analog_en[18]
  PIN mprj_io_analog_pol[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3102.265 210.965 3102.545 ;
    END
  END mprj_io_analog_pol[18]
  PIN mprj_io_analog_sel[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3087.085 210.965 3087.365 ;
    END
  END mprj_io_analog_sel[18]
  PIN mprj_io_dm[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3105.485 210.965 3105.765 ;
    END
  END mprj_io_dm[54]
  PIN mprj_io_dm[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3114.685 210.965 3114.965 ;
    END
  END mprj_io_dm[55]
  PIN mprj_io_dm[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3083.865 210.965 3084.145 ;
    END
  END mprj_io_dm[56]
  PIN mprj_io_holdover[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3080.645 210.965 3080.925 ;
    END
  END mprj_io_holdover[18]
  PIN mprj_io_ib_mode_sel[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3065.465 210.965 3065.745 ;
    END
  END mprj_io_ib_mode_sel[18]
  PIN mprj_io_inp_dis[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3099.505 210.965 3099.785 ;
    END
  END mprj_io_inp_dis[18]
  PIN mprj_io_oeb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3062.245 210.965 3062.525 ;
    END
  END mprj_io_oeb[18]
  PIN mprj_io_out[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3077.885 210.965 3078.165 ;
    END
  END mprj_io_out[18]
  PIN mprj_io_slow_sel[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3123.885 210.965 3124.165 ;
    END
  END mprj_io_slow_sel[18]
  PIN mprj_io_vtrip_sel[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3068.685 210.965 3068.965 ;
    END
  END mprj_io_vtrip_sel[18]
  PIN mprj_io_in[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3133.085 210.965 3133.365 ;
    END
  END mprj_io_in[18]
  PIN mprj_io_in_3v3[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3059.485 210.965 3059.765 ;
    END
  END mprj_io_in_3v3[18]
  PIN mprj_gpio_analog[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2904.665 210.965 2904.945 ;
    END
  END mprj_gpio_analog[12]
  PIN mprj_gpio_noesd[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2895.465 210.965 2895.745 ;
    END
  END mprj_gpio_noesd[12]
  PIN mprj_io[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 2853.200 95.440 2915.800 ;
    END
  END mprj_io[30]
  PIN mprj_io_analog_en[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2892.705 210.965 2892.985 ;
    END
  END mprj_io_analog_en[19]
  PIN mprj_io_analog_pol[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2886.265 210.965 2886.545 ;
    END
  END mprj_io_analog_pol[19]
  PIN mprj_io_analog_sel[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2871.085 210.965 2871.365 ;
    END
  END mprj_io_analog_sel[19]
  PIN mprj_io_dm[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2889.485 210.965 2889.765 ;
    END
  END mprj_io_dm[57]
  PIN mprj_io_dm[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2898.685 210.965 2898.965 ;
    END
  END mprj_io_dm[58]
  PIN mprj_io_dm[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2867.865 210.965 2868.145 ;
    END
  END mprj_io_dm[59]
  PIN mprj_io_holdover[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2864.645 210.965 2864.925 ;
    END
  END mprj_io_holdover[19]
  PIN mprj_io_ib_mode_sel[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2849.465 210.965 2849.745 ;
    END
  END mprj_io_ib_mode_sel[19]
  PIN mprj_io_inp_dis[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2883.505 210.965 2883.785 ;
    END
  END mprj_io_inp_dis[19]
  PIN mprj_io_oeb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2846.245 210.965 2846.525 ;
    END
  END mprj_io_oeb[19]
  PIN mprj_io_out[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2861.885 210.965 2862.165 ;
    END
  END mprj_io_out[19]
  PIN mprj_io_slow_sel[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2907.885 210.965 2908.165 ;
    END
  END mprj_io_slow_sel[19]
  PIN mprj_io_vtrip_sel[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2852.685 210.965 2852.965 ;
    END
  END mprj_io_vtrip_sel[19]
  PIN mprj_io_in[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2917.085 210.965 2917.365 ;
    END
  END mprj_io_in[19]
  PIN mprj_io_in_3v3[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2843.485 210.965 2843.765 ;
    END
  END mprj_io_in_3v3[19]
  PIN mprj_gpio_analog[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2688.665 210.965 2688.945 ;
    END
  END mprj_gpio_analog[13]
  PIN mprj_gpio_noesd[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2679.465 210.965 2679.745 ;
    END
  END mprj_gpio_noesd[13]
  PIN mprj_io[31]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 2637.200 95.440 2699.800 ;
    END
  END mprj_io[31]
  PIN mprj_io_analog_en[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2676.705 210.965 2676.985 ;
    END
  END mprj_io_analog_en[20]
  PIN mprj_io_analog_pol[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2670.265 210.965 2670.545 ;
    END
  END mprj_io_analog_pol[20]
  PIN mprj_io_analog_sel[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2655.085 210.965 2655.365 ;
    END
  END mprj_io_analog_sel[20]
  PIN mprj_io_dm[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2673.485 210.965 2673.765 ;
    END
  END mprj_io_dm[60]
  PIN mprj_io_dm[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2682.685 210.965 2682.965 ;
    END
  END mprj_io_dm[61]
  PIN mprj_io_dm[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2651.865 210.965 2652.145 ;
    END
  END mprj_io_dm[62]
  PIN mprj_io_holdover[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2648.645 210.965 2648.925 ;
    END
  END mprj_io_holdover[20]
  PIN mprj_io_ib_mode_sel[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2633.465 210.965 2633.745 ;
    END
  END mprj_io_ib_mode_sel[20]
  PIN mprj_io_inp_dis[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2667.505 210.965 2667.785 ;
    END
  END mprj_io_inp_dis[20]
  PIN mprj_io_oeb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2630.245 210.965 2630.525 ;
    END
  END mprj_io_oeb[20]
  PIN mprj_io_out[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2645.885 210.965 2646.165 ;
    END
  END mprj_io_out[20]
  PIN mprj_io_slow_sel[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2691.885 210.965 2692.165 ;
    END
  END mprj_io_slow_sel[20]
  PIN mprj_io_vtrip_sel[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2636.685 210.965 2636.965 ;
    END
  END mprj_io_vtrip_sel[20]
  PIN mprj_io_in[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2701.085 210.965 2701.365 ;
    END
  END mprj_io_in[20]
  PIN mprj_io_in_3v3[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2627.485 210.965 2627.765 ;
    END
  END mprj_io_in_3v3[20]
  PIN mprj_gpio_analog[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2050.665 210.965 2050.945 ;
    END
  END mprj_gpio_analog[14]
  PIN mprj_gpio_noesd[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2041.465 210.965 2041.745 ;
    END
  END mprj_gpio_noesd[14]
  PIN mprj_io[32]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 1999.200 95.440 2061.800 ;
    END
  END mprj_io[32]
  PIN mprj_io_analog_en[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2038.705 210.965 2038.985 ;
    END
  END mprj_io_analog_en[21]
  PIN mprj_io_analog_pol[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2032.265 210.965 2032.545 ;
    END
  END mprj_io_analog_pol[21]
  PIN mprj_io_analog_sel[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2017.085 210.965 2017.365 ;
    END
  END mprj_io_analog_sel[21]
  PIN mprj_io_dm[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2035.485 210.965 2035.765 ;
    END
  END mprj_io_dm[63]
  PIN mprj_io_dm[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2044.685 210.965 2044.965 ;
    END
  END mprj_io_dm[64]
  PIN mprj_io_dm[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2013.865 210.965 2014.145 ;
    END
  END mprj_io_dm[65]
  PIN mprj_io_holdover[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2010.645 210.965 2010.925 ;
    END
  END mprj_io_holdover[21]
  PIN mprj_io_ib_mode_sel[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1995.465 210.965 1995.745 ;
    END
  END mprj_io_ib_mode_sel[21]
  PIN mprj_io_inp_dis[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2029.505 210.965 2029.785 ;
    END
  END mprj_io_inp_dis[21]
  PIN mprj_io_oeb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1992.245 210.965 1992.525 ;
    END
  END mprj_io_oeb[21]
  PIN mprj_io_out[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2007.885 210.965 2008.165 ;
    END
  END mprj_io_out[21]
  PIN mprj_io_slow_sel[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2053.885 210.965 2054.165 ;
    END
  END mprj_io_slow_sel[21]
  PIN mprj_io_vtrip_sel[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1998.685 210.965 1998.965 ;
    END
  END mprj_io_vtrip_sel[21]
  PIN mprj_io_in[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2063.085 210.965 2063.365 ;
    END
  END mprj_io_in[21]
  PIN mprj_io_in_3v3[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1989.485 210.965 1989.765 ;
    END
  END mprj_io_in_3v3[21]
  PIN mprj_gpio_analog[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1834.665 210.965 1834.945 ;
    END
  END mprj_gpio_analog[15]
  PIN mprj_gpio_noesd[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1825.465 210.965 1825.745 ;
    END
  END mprj_gpio_noesd[15]
  PIN mprj_io[33]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 1783.200 95.440 1845.800 ;
    END
  END mprj_io[33]
  PIN mprj_io_analog_en[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1822.705 210.965 1822.985 ;
    END
  END mprj_io_analog_en[22]
  PIN mprj_io_analog_pol[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1816.265 210.965 1816.545 ;
    END
  END mprj_io_analog_pol[22]
  PIN mprj_io_analog_sel[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1801.085 210.965 1801.365 ;
    END
  END mprj_io_analog_sel[22]
  PIN mprj_io_dm[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1819.485 210.965 1819.765 ;
    END
  END mprj_io_dm[66]
  PIN mprj_io_dm[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1828.685 210.965 1828.965 ;
    END
  END mprj_io_dm[67]
  PIN mprj_io_dm[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1797.865 210.965 1798.145 ;
    END
  END mprj_io_dm[68]
  PIN mprj_io_holdover[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1794.645 210.965 1794.925 ;
    END
  END mprj_io_holdover[22]
  PIN mprj_io_ib_mode_sel[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1779.465 210.965 1779.745 ;
    END
  END mprj_io_ib_mode_sel[22]
  PIN mprj_io_inp_dis[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1813.505 210.965 1813.785 ;
    END
  END mprj_io_inp_dis[22]
  PIN mprj_io_oeb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1776.245 210.965 1776.525 ;
    END
  END mprj_io_oeb[22]
  PIN mprj_io_out[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1791.885 210.965 1792.165 ;
    END
  END mprj_io_out[22]
  PIN mprj_io_slow_sel[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1837.885 210.965 1838.165 ;
    END
  END mprj_io_slow_sel[22]
  PIN mprj_io_vtrip_sel[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1782.685 210.965 1782.965 ;
    END
  END mprj_io_vtrip_sel[22]
  PIN mprj_io_in[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1847.085 210.965 1847.365 ;
    END
  END mprj_io_in[22]
  PIN mprj_io_in_3v3[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1773.485 210.965 1773.765 ;
    END
  END mprj_io_in_3v3[22]
  PIN mprj_gpio_analog[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1618.665 210.965 1618.945 ;
    END
  END mprj_gpio_analog[16]
  PIN mprj_gpio_noesd[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1609.465 210.965 1609.745 ;
    END
  END mprj_gpio_noesd[16]
  PIN mprj_io[34]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 1567.200 95.440 1629.800 ;
    END
  END mprj_io[34]
  PIN mprj_io_analog_en[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1606.705 210.965 1606.985 ;
    END
  END mprj_io_analog_en[23]
  PIN mprj_io_analog_pol[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1600.265 210.965 1600.545 ;
    END
  END mprj_io_analog_pol[23]
  PIN mprj_io_analog_sel[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1585.085 210.965 1585.365 ;
    END
  END mprj_io_analog_sel[23]
  PIN mprj_io_dm[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1603.485 210.965 1603.765 ;
    END
  END mprj_io_dm[69]
  PIN mprj_io_dm[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1612.685 210.965 1612.965 ;
    END
  END mprj_io_dm[70]
  PIN mprj_io_dm[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1581.865 210.965 1582.145 ;
    END
  END mprj_io_dm[71]
  PIN mprj_io_holdover[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1578.645 210.965 1578.925 ;
    END
  END mprj_io_holdover[23]
  PIN mprj_io_ib_mode_sel[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1563.465 210.965 1563.745 ;
    END
  END mprj_io_ib_mode_sel[23]
  PIN mprj_io_inp_dis[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1597.505 210.965 1597.785 ;
    END
  END mprj_io_inp_dis[23]
  PIN mprj_io_oeb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1560.245 210.965 1560.525 ;
    END
  END mprj_io_oeb[23]
  PIN mprj_io_out[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1575.885 210.965 1576.165 ;
    END
  END mprj_io_out[23]
  PIN mprj_io_slow_sel[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1621.885 210.965 1622.165 ;
    END
  END mprj_io_slow_sel[23]
  PIN mprj_io_vtrip_sel[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1566.685 210.965 1566.965 ;
    END
  END mprj_io_vtrip_sel[23]
  PIN mprj_io_in[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1631.085 210.965 1631.365 ;
    END
  END mprj_io_in[23]
  PIN mprj_io_in_3v3[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1557.485 210.965 1557.765 ;
    END
  END mprj_io_in_3v3[23]
  PIN porb_h
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 3377.130 4378.555 3377.410 4378.585 ;
        RECT 3371.820 4378.275 3377.410 4378.555 ;
        RECT 3377.130 4378.245 3377.410 4378.275 ;
        RECT 3377.355 4356.935 3377.635 4356.965 ;
        RECT 3371.875 4356.655 3377.635 4356.935 ;
        RECT 3377.355 4356.625 3377.635 4356.655 ;
        RECT 210.340 3957.065 213.195 3957.345 ;
        RECT 210.340 3935.435 213.175 3935.715 ;
        RECT 3377.130 3932.555 3377.410 3932.585 ;
        RECT 3371.820 3932.275 3377.410 3932.555 ;
        RECT 3377.130 3932.245 3377.410 3932.275 ;
        RECT 3377.355 3910.935 3377.635 3910.965 ;
        RECT 3371.875 3910.655 3377.635 3910.935 ;
        RECT 3377.355 3910.625 3377.635 3910.655 ;
        RECT 210.340 3741.065 213.195 3741.345 ;
        RECT 210.340 3719.435 213.175 3719.715 ;
        RECT 3377.130 3707.555 3377.410 3707.585 ;
        RECT 3371.820 3707.275 3377.410 3707.555 ;
        RECT 3377.130 3707.245 3377.410 3707.275 ;
        RECT 3377.355 3685.935 3377.635 3685.965 ;
        RECT 3371.875 3685.655 3377.635 3685.935 ;
        RECT 3377.355 3685.625 3377.635 3685.655 ;
        RECT 210.340 3525.065 213.195 3525.345 ;
        RECT 210.340 3503.435 213.175 3503.715 ;
        RECT 3377.130 3482.555 3377.410 3482.585 ;
        RECT 3371.820 3482.275 3377.410 3482.555 ;
        RECT 3377.130 3482.245 3377.410 3482.275 ;
        RECT 3377.355 3460.935 3377.635 3460.965 ;
        RECT 3371.875 3460.655 3377.635 3460.935 ;
        RECT 3377.355 3460.625 3377.635 3460.655 ;
        RECT 210.340 3309.065 213.195 3309.345 ;
        RECT 210.340 3287.435 213.175 3287.715 ;
        RECT 3377.130 3256.555 3377.410 3256.585 ;
        RECT 3371.820 3256.275 3377.410 3256.555 ;
        RECT 3377.130 3256.245 3377.410 3256.275 ;
        RECT 3377.355 3234.935 3377.635 3234.965 ;
        RECT 3371.875 3234.655 3377.635 3234.935 ;
        RECT 3377.355 3234.625 3377.635 3234.655 ;
        RECT 210.340 3093.065 213.195 3093.345 ;
        RECT 210.340 3071.435 213.175 3071.715 ;
        RECT 3377.130 3031.555 3377.410 3031.585 ;
        RECT 3371.820 3031.275 3377.410 3031.555 ;
        RECT 3377.130 3031.245 3377.410 3031.275 ;
        RECT 3377.355 3009.935 3377.635 3009.965 ;
        RECT 3375.665 3009.760 3377.635 3009.935 ;
        RECT 3371.875 3009.655 3377.635 3009.760 ;
        RECT 3371.875 3009.480 3375.945 3009.655 ;
        RECT 3377.355 3009.625 3377.635 3009.655 ;
        RECT 210.340 2877.065 213.195 2877.345 ;
        RECT 210.340 2855.435 213.175 2855.715 ;
        RECT 3377.130 2805.555 3377.410 2805.585 ;
        RECT 3371.820 2805.275 3377.410 2805.555 ;
        RECT 3377.130 2805.245 3377.410 2805.275 ;
        RECT 3377.355 2783.935 3377.635 2783.965 ;
        RECT 3371.875 2783.655 3377.635 2783.935 ;
        RECT 3377.355 2783.625 3377.635 2783.655 ;
        RECT 210.340 2661.065 213.195 2661.345 ;
        RECT 210.340 2639.435 213.175 2639.715 ;
        RECT 210.340 2023.065 213.195 2023.345 ;
        RECT 210.340 2001.435 213.175 2001.715 ;
        RECT 3377.130 1919.555 3377.410 1919.585 ;
        RECT 3371.820 1919.275 3377.410 1919.555 ;
        RECT 3377.130 1919.245 3377.410 1919.275 ;
        RECT 3377.355 1897.935 3377.635 1897.965 ;
        RECT 3371.875 1897.655 3377.635 1897.935 ;
        RECT 3377.355 1897.625 3377.635 1897.655 ;
        RECT 210.340 1807.065 213.195 1807.345 ;
        RECT 210.340 1785.435 213.175 1785.715 ;
        RECT 3377.130 1693.555 3377.410 1693.585 ;
        RECT 3371.820 1693.275 3377.410 1693.555 ;
        RECT 3377.130 1693.245 3377.410 1693.275 ;
        RECT 3377.355 1671.935 3377.635 1671.965 ;
        RECT 3371.875 1671.655 3377.635 1671.935 ;
        RECT 3377.355 1671.625 3377.635 1671.655 ;
        RECT 210.340 1591.065 213.195 1591.345 ;
        RECT 210.340 1569.435 213.175 1569.715 ;
        RECT 3377.130 1468.555 3377.410 1468.585 ;
        RECT 3371.820 1468.275 3377.410 1468.555 ;
        RECT 3377.130 1468.245 3377.410 1468.275 ;
        RECT 3377.355 1446.935 3377.635 1446.965 ;
        RECT 3371.875 1446.655 3377.635 1446.935 ;
        RECT 3377.355 1446.625 3377.635 1446.655 ;
        RECT 210.340 1375.065 213.195 1375.345 ;
        RECT 210.340 1353.435 213.175 1353.715 ;
        RECT 3377.130 1243.555 3377.410 1243.585 ;
        RECT 3371.820 1243.275 3377.410 1243.555 ;
        RECT 3377.130 1243.245 3377.410 1243.275 ;
        RECT 3377.355 1221.935 3377.635 1221.965 ;
        RECT 3371.875 1221.655 3377.635 1221.935 ;
        RECT 3377.355 1221.625 3377.635 1221.655 ;
        RECT 210.340 1159.065 213.195 1159.345 ;
        RECT 210.340 1137.435 213.175 1137.715 ;
        RECT 3377.130 1017.555 3377.410 1017.585 ;
        RECT 3371.820 1017.275 3377.410 1017.555 ;
        RECT 3377.130 1017.245 3377.410 1017.275 ;
        RECT 3377.355 995.935 3377.635 995.965 ;
        RECT 3371.875 995.655 3377.635 995.935 ;
        RECT 3377.355 995.625 3377.635 995.655 ;
        RECT 210.340 943.065 213.195 943.345 ;
        RECT 212.865 906.330 213.185 906.390 ;
        RECT 207.070 906.190 213.185 906.330 ;
        RECT 207.070 887.355 207.210 906.190 ;
        RECT 212.865 906.130 213.185 906.190 ;
        RECT 207.070 887.215 210.210 887.355 ;
        RECT 210.070 209.305 210.210 887.215 ;
        RECT 3377.130 792.555 3377.410 792.585 ;
        RECT 3371.820 792.275 3377.410 792.555 ;
        RECT 3377.130 792.245 3377.410 792.275 ;
        RECT 3377.355 770.935 3377.635 770.965 ;
        RECT 3371.875 770.655 3377.635 770.935 ;
        RECT 3377.355 770.625 3377.635 770.655 ;
        RECT 3377.130 566.555 3377.410 566.585 ;
        RECT 3371.820 566.275 3377.410 566.555 ;
        RECT 3377.130 566.245 3377.410 566.275 ;
        RECT 3377.355 544.935 3377.635 544.965 ;
        RECT 3371.875 544.655 3377.635 544.935 ;
        RECT 3377.355 544.625 3377.635 544.655 ;
        RECT 3371.815 210.475 3372.135 210.535 ;
        RECT 3182.580 210.335 3372.135 210.475 ;
        RECT 976.625 209.305 976.965 209.435 ;
        RECT 998.245 209.305 998.585 209.435 ;
        RECT 1519.625 209.305 1519.965 209.355 ;
        RECT 1541.245 209.305 1541.585 209.365 ;
        RECT 1793.625 209.305 1793.965 209.355 ;
        RECT 1815.245 209.305 1815.585 209.365 ;
        RECT 2067.625 209.305 2067.965 209.355 ;
        RECT 2089.245 209.305 2089.585 209.365 ;
        RECT 2341.625 209.305 2341.965 209.375 ;
        RECT 2363.245 209.305 2363.585 209.380 ;
        RECT 2615.625 209.305 2615.965 209.365 ;
        RECT 2637.245 209.305 2637.585 209.355 ;
        RECT 3182.580 209.305 3182.720 210.335 ;
        RECT 3371.815 210.275 3372.135 210.335 ;
        RECT 210.070 209.165 3182.720 209.305 ;
        RECT 725.425 209.045 725.745 209.165 ;
        RECT 976.625 209.155 976.965 209.165 ;
        RECT 998.245 209.155 998.585 209.165 ;
        RECT 1519.625 209.075 1519.965 209.165 ;
        RECT 1541.245 209.085 1541.585 209.165 ;
        RECT 1793.625 209.075 1793.965 209.165 ;
        RECT 1815.245 209.085 1815.585 209.165 ;
        RECT 2067.625 209.075 2067.965 209.165 ;
        RECT 2089.245 209.085 2089.585 209.165 ;
        RECT 2341.625 209.095 2341.965 209.165 ;
        RECT 2363.245 209.100 2363.585 209.165 ;
        RECT 2615.625 209.085 2615.965 209.165 ;
        RECT 2637.245 209.075 2637.585 209.165 ;
      LAYER via ;
        RECT 3371.850 4378.275 3372.130 4378.555 ;
        RECT 3377.130 4378.275 3377.410 4378.555 ;
        RECT 3371.905 4356.655 3372.185 4356.935 ;
        RECT 3377.355 4356.655 3377.635 4356.935 ;
        RECT 210.370 3957.065 210.650 3957.345 ;
        RECT 212.885 3957.065 213.165 3957.345 ;
        RECT 210.370 3935.435 210.650 3935.715 ;
        RECT 212.865 3935.435 213.145 3935.715 ;
        RECT 3371.850 3932.275 3372.130 3932.555 ;
        RECT 3377.130 3932.275 3377.410 3932.555 ;
        RECT 3371.905 3910.655 3372.185 3910.935 ;
        RECT 3377.355 3910.655 3377.635 3910.935 ;
        RECT 210.370 3741.065 210.650 3741.345 ;
        RECT 212.885 3741.065 213.165 3741.345 ;
        RECT 210.370 3719.435 210.650 3719.715 ;
        RECT 212.865 3719.435 213.145 3719.715 ;
        RECT 3371.850 3707.275 3372.130 3707.555 ;
        RECT 3377.130 3707.275 3377.410 3707.555 ;
        RECT 3371.905 3685.655 3372.185 3685.935 ;
        RECT 3377.355 3685.655 3377.635 3685.935 ;
        RECT 210.370 3525.065 210.650 3525.345 ;
        RECT 212.885 3525.065 213.165 3525.345 ;
        RECT 210.370 3503.435 210.650 3503.715 ;
        RECT 212.865 3503.435 213.145 3503.715 ;
        RECT 3371.850 3482.275 3372.130 3482.555 ;
        RECT 3377.130 3482.275 3377.410 3482.555 ;
        RECT 3371.905 3460.655 3372.185 3460.935 ;
        RECT 3377.355 3460.655 3377.635 3460.935 ;
        RECT 210.370 3309.065 210.650 3309.345 ;
        RECT 212.885 3309.065 213.165 3309.345 ;
        RECT 210.370 3287.435 210.650 3287.715 ;
        RECT 212.865 3287.435 213.145 3287.715 ;
        RECT 3371.850 3256.275 3372.130 3256.555 ;
        RECT 3377.130 3256.275 3377.410 3256.555 ;
        RECT 3371.905 3234.655 3372.185 3234.935 ;
        RECT 3377.355 3234.655 3377.635 3234.935 ;
        RECT 210.370 3093.065 210.650 3093.345 ;
        RECT 212.885 3093.065 213.165 3093.345 ;
        RECT 210.370 3071.435 210.650 3071.715 ;
        RECT 212.865 3071.435 213.145 3071.715 ;
        RECT 3371.850 3031.275 3372.130 3031.555 ;
        RECT 3377.130 3031.275 3377.410 3031.555 ;
        RECT 3371.905 3009.480 3372.185 3009.760 ;
        RECT 3377.355 3009.655 3377.635 3009.935 ;
        RECT 210.370 2877.065 210.650 2877.345 ;
        RECT 212.885 2877.065 213.165 2877.345 ;
        RECT 210.370 2855.435 210.650 2855.715 ;
        RECT 212.865 2855.435 213.145 2855.715 ;
        RECT 3371.850 2805.275 3372.130 2805.555 ;
        RECT 3377.130 2805.275 3377.410 2805.555 ;
        RECT 3371.905 2783.655 3372.185 2783.935 ;
        RECT 3377.355 2783.655 3377.635 2783.935 ;
        RECT 210.370 2661.065 210.650 2661.345 ;
        RECT 212.885 2661.065 213.165 2661.345 ;
        RECT 210.370 2639.435 210.650 2639.715 ;
        RECT 212.865 2639.435 213.145 2639.715 ;
        RECT 210.370 2023.065 210.650 2023.345 ;
        RECT 212.885 2023.065 213.165 2023.345 ;
        RECT 210.370 2001.435 210.650 2001.715 ;
        RECT 212.865 2001.435 213.145 2001.715 ;
        RECT 3371.850 1919.275 3372.130 1919.555 ;
        RECT 3377.130 1919.275 3377.410 1919.555 ;
        RECT 3371.905 1897.655 3372.185 1897.935 ;
        RECT 3377.355 1897.655 3377.635 1897.935 ;
        RECT 210.370 1807.065 210.650 1807.345 ;
        RECT 212.885 1807.065 213.165 1807.345 ;
        RECT 210.370 1785.435 210.650 1785.715 ;
        RECT 212.865 1785.435 213.145 1785.715 ;
        RECT 3371.850 1693.275 3372.130 1693.555 ;
        RECT 3377.130 1693.275 3377.410 1693.555 ;
        RECT 3371.905 1671.655 3372.185 1671.935 ;
        RECT 3377.355 1671.655 3377.635 1671.935 ;
        RECT 210.370 1591.065 210.650 1591.345 ;
        RECT 212.885 1591.065 213.165 1591.345 ;
        RECT 210.370 1569.435 210.650 1569.715 ;
        RECT 212.865 1569.435 213.145 1569.715 ;
        RECT 3371.850 1468.275 3372.130 1468.555 ;
        RECT 3377.130 1468.275 3377.410 1468.555 ;
        RECT 3371.905 1446.655 3372.185 1446.935 ;
        RECT 3377.355 1446.655 3377.635 1446.935 ;
        RECT 210.370 1375.065 210.650 1375.345 ;
        RECT 212.885 1375.065 213.165 1375.345 ;
        RECT 210.370 1353.435 210.650 1353.715 ;
        RECT 212.865 1353.435 213.145 1353.715 ;
        RECT 3371.850 1243.275 3372.130 1243.555 ;
        RECT 3377.130 1243.275 3377.410 1243.555 ;
        RECT 3371.905 1221.655 3372.185 1221.935 ;
        RECT 3377.355 1221.655 3377.635 1221.935 ;
        RECT 210.370 1159.065 210.650 1159.345 ;
        RECT 212.885 1159.065 213.165 1159.345 ;
        RECT 210.370 1137.435 210.650 1137.715 ;
        RECT 212.865 1137.435 213.145 1137.715 ;
        RECT 3371.850 1017.275 3372.130 1017.555 ;
        RECT 3377.130 1017.275 3377.410 1017.555 ;
        RECT 3371.905 995.655 3372.185 995.935 ;
        RECT 3377.355 995.655 3377.635 995.935 ;
        RECT 210.370 943.065 210.650 943.345 ;
        RECT 212.885 943.065 213.165 943.345 ;
        RECT 212.895 906.130 213.155 906.390 ;
        RECT 3371.850 792.275 3372.130 792.555 ;
        RECT 3377.130 792.275 3377.410 792.555 ;
        RECT 3371.905 770.655 3372.185 770.935 ;
        RECT 3377.355 770.655 3377.635 770.935 ;
        RECT 3371.850 566.275 3372.130 566.555 ;
        RECT 3377.130 566.275 3377.410 566.555 ;
        RECT 3371.905 544.655 3372.185 544.935 ;
        RECT 3377.355 544.655 3377.635 544.935 ;
        RECT 725.455 209.045 725.715 209.305 ;
        RECT 976.655 209.155 976.935 209.435 ;
        RECT 998.275 209.155 998.555 209.435 ;
        RECT 1519.655 209.075 1519.935 209.355 ;
        RECT 1541.275 209.085 1541.555 209.365 ;
        RECT 1793.655 209.075 1793.935 209.355 ;
        RECT 1815.275 209.085 1815.555 209.365 ;
        RECT 2067.655 209.075 2067.935 209.355 ;
        RECT 2089.275 209.085 2089.555 209.365 ;
        RECT 2341.655 209.095 2341.935 209.375 ;
        RECT 2363.275 209.100 2363.555 209.380 ;
        RECT 2615.655 209.085 2615.935 209.365 ;
        RECT 2637.275 209.075 2637.555 209.355 ;
        RECT 3371.845 210.275 3372.105 210.535 ;
      LAYER met2 ;
        RECT 3371.880 4378.585 3372.070 4378.735 ;
        RECT 3371.850 4378.245 3372.130 4378.585 ;
        RECT 3377.035 4378.275 3379.435 4378.555 ;
        RECT 3371.880 4356.965 3372.070 4378.245 ;
        RECT 3371.880 4356.625 3372.185 4356.965 ;
        RECT 3377.035 4356.655 3379.435 4356.935 ;
        RECT 212.930 3957.375 213.125 3957.545 ;
        RECT 210.370 3957.345 210.650 3957.375 ;
        RECT 208.565 3957.065 210.965 3957.345 ;
        RECT 210.155 3957.055 210.965 3957.065 ;
        RECT 210.370 3957.035 210.650 3957.055 ;
        RECT 212.885 3957.035 213.165 3957.375 ;
        RECT 212.930 3935.745 213.125 3957.035 ;
        RECT 210.370 3935.725 210.650 3935.745 ;
        RECT 208.565 3935.445 210.965 3935.725 ;
        RECT 210.085 3935.435 210.965 3935.445 ;
        RECT 210.370 3935.405 210.650 3935.435 ;
        RECT 212.865 3935.405 213.145 3935.745 ;
        RECT 212.930 3741.375 213.125 3935.405 ;
        RECT 3371.880 3932.585 3372.070 4356.625 ;
        RECT 3371.850 3932.245 3372.130 3932.585 ;
        RECT 3377.035 3932.275 3379.435 3932.555 ;
        RECT 3371.880 3910.965 3372.070 3932.245 ;
        RECT 3371.880 3910.625 3372.185 3910.965 ;
        RECT 3377.035 3910.655 3379.435 3910.935 ;
        RECT 210.370 3741.345 210.650 3741.375 ;
        RECT 208.565 3741.065 210.965 3741.345 ;
        RECT 210.155 3741.055 210.965 3741.065 ;
        RECT 210.370 3741.035 210.650 3741.055 ;
        RECT 212.885 3741.035 213.165 3741.375 ;
        RECT 212.930 3719.745 213.125 3741.035 ;
        RECT 210.370 3719.725 210.650 3719.745 ;
        RECT 208.565 3719.445 210.965 3719.725 ;
        RECT 210.085 3719.435 210.965 3719.445 ;
        RECT 210.370 3719.405 210.650 3719.435 ;
        RECT 212.865 3719.405 213.145 3719.745 ;
        RECT 212.930 3525.375 213.125 3719.405 ;
        RECT 3371.880 3707.585 3372.070 3910.625 ;
        RECT 3371.850 3707.245 3372.130 3707.585 ;
        RECT 3377.035 3707.275 3379.435 3707.555 ;
        RECT 3371.880 3685.965 3372.070 3707.245 ;
        RECT 3371.880 3685.625 3372.185 3685.965 ;
        RECT 3377.035 3685.655 3379.435 3685.935 ;
        RECT 210.370 3525.345 210.650 3525.375 ;
        RECT 208.565 3525.065 210.965 3525.345 ;
        RECT 210.155 3525.055 210.965 3525.065 ;
        RECT 210.370 3525.035 210.650 3525.055 ;
        RECT 212.885 3525.035 213.165 3525.375 ;
        RECT 212.930 3503.745 213.125 3525.035 ;
        RECT 210.370 3503.725 210.650 3503.745 ;
        RECT 208.565 3503.445 210.965 3503.725 ;
        RECT 210.085 3503.435 210.965 3503.445 ;
        RECT 210.370 3503.405 210.650 3503.435 ;
        RECT 212.865 3503.405 213.145 3503.745 ;
        RECT 212.930 3309.375 213.125 3503.405 ;
        RECT 3371.880 3482.585 3372.070 3685.625 ;
        RECT 3371.850 3482.245 3372.130 3482.585 ;
        RECT 3377.035 3482.275 3379.435 3482.555 ;
        RECT 3371.880 3460.965 3372.070 3482.245 ;
        RECT 3371.880 3460.625 3372.185 3460.965 ;
        RECT 3377.035 3460.655 3379.435 3460.935 ;
        RECT 210.370 3309.345 210.650 3309.375 ;
        RECT 208.565 3309.065 210.965 3309.345 ;
        RECT 210.155 3309.055 210.965 3309.065 ;
        RECT 210.370 3309.035 210.650 3309.055 ;
        RECT 212.885 3309.035 213.165 3309.375 ;
        RECT 212.930 3287.745 213.125 3309.035 ;
        RECT 210.370 3287.725 210.650 3287.745 ;
        RECT 208.565 3287.445 210.965 3287.725 ;
        RECT 210.085 3287.435 210.965 3287.445 ;
        RECT 210.370 3287.405 210.650 3287.435 ;
        RECT 212.865 3287.405 213.145 3287.745 ;
        RECT 212.930 3093.375 213.125 3287.405 ;
        RECT 3371.880 3256.585 3372.070 3460.625 ;
        RECT 3371.850 3256.245 3372.130 3256.585 ;
        RECT 3377.035 3256.275 3379.435 3256.555 ;
        RECT 3371.880 3234.965 3372.070 3256.245 ;
        RECT 3371.880 3234.625 3372.185 3234.965 ;
        RECT 3377.035 3234.655 3379.435 3234.935 ;
        RECT 210.370 3093.345 210.650 3093.375 ;
        RECT 208.565 3093.065 210.965 3093.345 ;
        RECT 210.155 3093.055 210.965 3093.065 ;
        RECT 210.370 3093.035 210.650 3093.055 ;
        RECT 212.885 3093.035 213.165 3093.375 ;
        RECT 212.930 3071.745 213.125 3093.035 ;
        RECT 210.370 3071.725 210.650 3071.745 ;
        RECT 208.565 3071.445 210.965 3071.725 ;
        RECT 210.085 3071.435 210.965 3071.445 ;
        RECT 210.370 3071.405 210.650 3071.435 ;
        RECT 212.865 3071.405 213.145 3071.745 ;
        RECT 212.930 2877.375 213.125 3071.405 ;
        RECT 3371.880 3031.585 3372.070 3234.625 ;
        RECT 3371.850 3031.245 3372.130 3031.585 ;
        RECT 3377.035 3031.275 3379.435 3031.555 ;
        RECT 3371.880 3009.790 3372.070 3031.245 ;
        RECT 3371.880 3009.450 3372.185 3009.790 ;
        RECT 3377.035 3009.655 3379.435 3009.935 ;
        RECT 210.370 2877.345 210.650 2877.375 ;
        RECT 208.565 2877.065 210.965 2877.345 ;
        RECT 210.155 2877.055 210.965 2877.065 ;
        RECT 210.370 2877.035 210.650 2877.055 ;
        RECT 212.885 2877.035 213.165 2877.375 ;
        RECT 212.930 2855.745 213.125 2877.035 ;
        RECT 210.370 2855.725 210.650 2855.745 ;
        RECT 208.565 2855.445 210.965 2855.725 ;
        RECT 210.085 2855.435 210.965 2855.445 ;
        RECT 210.370 2855.405 210.650 2855.435 ;
        RECT 212.865 2855.405 213.145 2855.745 ;
        RECT 212.930 2661.375 213.125 2855.405 ;
        RECT 3371.880 2805.585 3372.070 3009.450 ;
        RECT 3371.850 2805.245 3372.130 2805.585 ;
        RECT 3377.035 2805.275 3379.435 2805.555 ;
        RECT 3371.880 2783.965 3372.070 2805.245 ;
        RECT 3371.880 2783.625 3372.185 2783.965 ;
        RECT 3377.035 2783.655 3379.435 2783.935 ;
        RECT 210.370 2661.345 210.650 2661.375 ;
        RECT 208.565 2661.065 210.965 2661.345 ;
        RECT 210.155 2661.055 210.965 2661.065 ;
        RECT 210.370 2661.035 210.650 2661.055 ;
        RECT 212.885 2661.035 213.165 2661.375 ;
        RECT 212.930 2639.745 213.125 2661.035 ;
        RECT 210.370 2639.725 210.650 2639.745 ;
        RECT 208.565 2639.445 210.965 2639.725 ;
        RECT 210.085 2639.435 210.965 2639.445 ;
        RECT 210.370 2639.405 210.650 2639.435 ;
        RECT 212.865 2639.405 213.145 2639.745 ;
        RECT 212.930 2023.375 213.125 2639.405 ;
        RECT 210.370 2023.345 210.650 2023.375 ;
        RECT 208.565 2023.065 210.965 2023.345 ;
        RECT 210.155 2023.055 210.965 2023.065 ;
        RECT 210.370 2023.035 210.650 2023.055 ;
        RECT 212.885 2023.035 213.165 2023.375 ;
        RECT 212.930 2001.745 213.125 2023.035 ;
        RECT 210.370 2001.725 210.650 2001.745 ;
        RECT 208.565 2001.445 210.965 2001.725 ;
        RECT 210.085 2001.435 210.965 2001.445 ;
        RECT 210.370 2001.405 210.650 2001.435 ;
        RECT 212.865 2001.405 213.145 2001.745 ;
        RECT 212.930 1807.375 213.125 2001.405 ;
        RECT 3371.880 1919.585 3372.070 2783.625 ;
        RECT 3371.850 1919.245 3372.130 1919.585 ;
        RECT 3377.035 1919.275 3379.435 1919.555 ;
        RECT 3371.880 1897.965 3372.070 1919.245 ;
        RECT 3371.880 1897.625 3372.185 1897.965 ;
        RECT 3377.035 1897.655 3379.435 1897.935 ;
        RECT 210.370 1807.345 210.650 1807.375 ;
        RECT 208.565 1807.065 210.965 1807.345 ;
        RECT 210.155 1807.055 210.965 1807.065 ;
        RECT 210.370 1807.035 210.650 1807.055 ;
        RECT 212.885 1807.035 213.165 1807.375 ;
        RECT 212.930 1785.745 213.125 1807.035 ;
        RECT 210.370 1785.725 210.650 1785.745 ;
        RECT 208.565 1785.445 210.965 1785.725 ;
        RECT 210.085 1785.435 210.965 1785.445 ;
        RECT 210.370 1785.405 210.650 1785.435 ;
        RECT 212.865 1785.405 213.145 1785.745 ;
        RECT 212.930 1591.375 213.125 1785.405 ;
        RECT 3371.880 1693.585 3372.070 1897.625 ;
        RECT 3371.850 1693.245 3372.130 1693.585 ;
        RECT 3377.035 1693.275 3379.435 1693.555 ;
        RECT 3371.880 1671.965 3372.070 1693.245 ;
        RECT 3371.880 1671.625 3372.185 1671.965 ;
        RECT 3377.035 1671.655 3379.435 1671.935 ;
        RECT 210.370 1591.345 210.650 1591.375 ;
        RECT 208.565 1591.065 210.965 1591.345 ;
        RECT 210.155 1591.055 210.965 1591.065 ;
        RECT 210.370 1591.035 210.650 1591.055 ;
        RECT 212.885 1591.035 213.165 1591.375 ;
        RECT 212.930 1569.745 213.125 1591.035 ;
        RECT 210.370 1569.725 210.650 1569.745 ;
        RECT 208.565 1569.445 210.965 1569.725 ;
        RECT 210.085 1569.435 210.965 1569.445 ;
        RECT 210.370 1569.405 210.650 1569.435 ;
        RECT 212.865 1569.405 213.145 1569.745 ;
        RECT 212.930 1375.375 213.125 1569.405 ;
        RECT 3371.880 1468.585 3372.070 1671.625 ;
        RECT 3371.850 1468.245 3372.130 1468.585 ;
        RECT 3377.035 1468.275 3379.435 1468.555 ;
        RECT 3371.880 1446.965 3372.070 1468.245 ;
        RECT 3371.880 1446.625 3372.185 1446.965 ;
        RECT 3377.035 1446.655 3379.435 1446.935 ;
        RECT 210.370 1375.345 210.650 1375.375 ;
        RECT 208.565 1375.065 210.965 1375.345 ;
        RECT 210.155 1375.055 210.965 1375.065 ;
        RECT 210.370 1375.035 210.650 1375.055 ;
        RECT 212.885 1375.035 213.165 1375.375 ;
        RECT 212.930 1353.745 213.125 1375.035 ;
        RECT 210.370 1353.725 210.650 1353.745 ;
        RECT 208.565 1353.445 210.965 1353.725 ;
        RECT 210.085 1353.435 210.965 1353.445 ;
        RECT 210.370 1353.405 210.650 1353.435 ;
        RECT 212.865 1353.405 213.145 1353.745 ;
        RECT 212.930 1159.375 213.125 1353.405 ;
        RECT 3371.880 1243.585 3372.070 1446.625 ;
        RECT 3371.850 1243.245 3372.130 1243.585 ;
        RECT 3377.035 1243.275 3379.435 1243.555 ;
        RECT 3371.880 1221.965 3372.070 1243.245 ;
        RECT 3371.880 1221.625 3372.185 1221.965 ;
        RECT 3377.035 1221.655 3379.435 1221.935 ;
        RECT 210.370 1159.345 210.650 1159.375 ;
        RECT 208.565 1159.065 210.965 1159.345 ;
        RECT 210.155 1159.055 210.965 1159.065 ;
        RECT 210.370 1159.035 210.650 1159.055 ;
        RECT 212.885 1159.035 213.165 1159.375 ;
        RECT 212.930 1137.745 213.125 1159.035 ;
        RECT 210.370 1137.725 210.650 1137.745 ;
        RECT 208.565 1137.445 210.965 1137.725 ;
        RECT 210.085 1137.435 210.965 1137.445 ;
        RECT 210.370 1137.405 210.650 1137.435 ;
        RECT 212.865 1137.405 213.145 1137.745 ;
        RECT 212.930 943.375 213.125 1137.405 ;
        RECT 3371.880 1017.585 3372.070 1221.625 ;
        RECT 3371.850 1017.245 3372.130 1017.585 ;
        RECT 3377.035 1017.275 3379.435 1017.555 ;
        RECT 3371.880 995.965 3372.070 1017.245 ;
        RECT 3371.880 995.625 3372.185 995.965 ;
        RECT 3377.035 995.655 3379.435 995.935 ;
        RECT 210.370 943.345 210.650 943.375 ;
        RECT 208.565 943.065 210.965 943.345 ;
        RECT 209.400 943.055 210.965 943.065 ;
        RECT 210.370 943.035 210.650 943.055 ;
        RECT 212.885 943.035 213.165 943.375 ;
        RECT 212.930 921.725 213.125 943.035 ;
        RECT 208.565 921.445 213.125 921.725 ;
        RECT 212.930 906.420 213.125 921.445 ;
        RECT 212.895 906.100 213.155 906.420 ;
        RECT 3371.880 792.585 3372.070 995.625 ;
        RECT 3371.850 792.245 3372.130 792.585 ;
        RECT 3377.035 792.275 3379.435 792.555 ;
        RECT 3371.880 770.965 3372.070 792.245 ;
        RECT 3371.880 770.625 3372.185 770.965 ;
        RECT 3377.035 770.655 3379.435 770.935 ;
        RECT 3371.880 566.585 3372.070 770.625 ;
        RECT 3371.850 566.245 3372.130 566.585 ;
        RECT 3377.035 566.275 3379.435 566.555 ;
        RECT 3371.880 544.965 3372.070 566.245 ;
        RECT 3371.880 544.625 3372.185 544.965 ;
        RECT 3377.035 544.655 3379.435 544.935 ;
        RECT 725.455 198.530 725.715 209.335 ;
        RECT 976.655 208.565 976.935 210.995 ;
        RECT 998.275 208.565 998.555 210.990 ;
        RECT 1519.655 208.565 1519.935 210.965 ;
        RECT 1541.275 208.565 1541.555 210.965 ;
        RECT 1793.655 208.565 1793.935 210.965 ;
        RECT 1815.275 208.565 1815.555 210.965 ;
        RECT 2067.655 208.565 2067.935 210.970 ;
        RECT 2089.275 208.565 2089.555 210.965 ;
        RECT 2341.655 208.565 2341.935 210.995 ;
        RECT 2363.275 208.565 2363.555 210.975 ;
        RECT 2615.655 208.565 2615.935 210.985 ;
        RECT 2637.275 208.565 2637.555 211.005 ;
        RECT 3371.880 210.565 3372.070 544.625 ;
        RECT 3371.845 210.245 3372.105 210.565 ;
    END
  END porb_h
  PIN resetb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 683.565 35.715 720.750 91.545 ;
    END
  END resetb
  PIN resetb_core_h
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.335 199.670 709.065 200.000 ;
    END
  END resetb_core_h
  PIN vdda
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 468.035 181.615 663.965 185.065 ;
    END
  END vdda
  PIN vssa
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 467.730 143.265 964.910 143.595 ;
    END
  END vssa
  PIN vssd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 467.730 158.370 664.270 158.415 ;
        RECT 467.730 153.810 664.345 158.370 ;
        RECT 467.730 153.765 664.270 153.810 ;
    END
  END vssd
  PIN mprj_analog[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3159.720 4988.000 3184.720 5070.350 ;
    END
  END mprj_analog[0]
  PIN mprj_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3142.050 5093.120 3202.890 5153.945 ;
    END
  END mprj_io[15]
  PIN mprj_analog[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2650.720 4988.000 2675.720 5070.350 ;
    END
  END mprj_analog[1]
  PIN mprj_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2633.050 5093.120 2693.890 5153.945 ;
    END
  END mprj_io[16]
  PIN mprj_analog[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2393.720 4988.000 2418.720 5070.350 ;
    END
  END mprj_analog[2]
  PIN mprj_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2376.050 5093.120 2436.890 5153.945 ;
    END
  END mprj_io[17]
  PIN mprj_analog[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3388.000 4783.280 3470.350 4808.280 ;
    END
  END mprj_analog[3]
  PIN mprj_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3493.120 4765.110 3553.945 4825.950 ;
    END
  END mprj_io[14]
  PIN mprj_analog[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1974.390 4988.000 2046.000 5003.685 ;
    END
  END mprj_analog[4]
  PIN mprj_clamp_high[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1974.390 4988.000 1998.290 5013.660 ;
    END
  END mprj_clamp_high[0]
  PIN mprj_clamp_low[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1924.495 4988.000 1948.395 4990.055 ;
    END
  END mprj_clamp_low[0]
  PIN mprj_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1931.050 5093.120 1991.890 5153.945 ;
    END
  END mprj_io[18]
  PIN vccd1_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3489.900 4548.330 3557.160 4602.730 ;
    END
  END vccd1_pad
  PIN vdda1_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3493.120 4099.110 3553.945 4159.950 ;
    END
  END vdda1_pad
  PIN vdda1_pad2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3493.120 2526.110 3553.945 2586.950 ;
    END
  END vdda1_pad2
  PIN vssa1_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2885.050 5093.120 2945.890 5153.945 ;
    END
  END vssa1_pad
  PIN vssa1_pad2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3493.120 2085.110 3553.945 2145.950 ;
    END
  END vssa1_pad2
  PIN vccd1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3353.800 4612.500 3382.205 4612.510 ;
        RECT 3353.800 4588.500 3382.810 4612.500 ;
        RECT 3353.800 4538.300 3382.810 4562.245 ;
        RECT 3353.640 2324.745 3381.780 2348.000 ;
      LAYER via3 ;
        RECT 3354.690 4589.300 3364.720 4611.820 ;
        RECT 3354.760 4538.900 3364.790 4561.420 ;
        RECT 3354.820 2325.480 3364.960 2347.120 ;
      LAYER met4 ;
        RECT 3354.080 4588.570 3367.090 4612.490 ;
        RECT 3354.140 4538.330 3367.060 4562.200 ;
        RECT 3354.130 2324.780 3367.060 2348.010 ;
      LAYER via4 ;
        RECT 3354.690 4589.300 3366.280 4611.820 ;
        RECT 3354.760 4538.900 3366.350 4561.420 ;
        RECT 3354.820 2325.480 3366.520 2347.120 ;
      LAYER met5 ;
        RECT 3354.100 486.470 3367.100 4958.900 ;
    END
  END vccd1
  PIN vdda1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3402.935 2152.035 3406.385 2299.960 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3444.405 2151.730 3444.735 2771.910 ;
    END
  END vssa1
  PIN vssd1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3353.800 4563.740 3382.810 4587.050 ;
        RECT 3353.640 2349.500 3381.780 2373.500 ;
        RECT 3353.640 2299.300 3381.780 2323.245 ;
      LAYER via3 ;
        RECT 3370.800 4564.470 3380.930 4586.350 ;
        RECT 3371.000 2350.360 3380.610 2372.790 ;
        RECT 3371.100 2300.070 3380.710 2322.500 ;
      LAYER met4 ;
        RECT 3370.090 4563.730 3383.080 4587.040 ;
        RECT 3370.130 2349.590 3382.970 2373.630 ;
        RECT 3370.130 2299.270 3382.970 2323.310 ;
      LAYER via4 ;
        RECT 3370.800 4564.470 3382.490 4586.350 ;
        RECT 3371.000 2350.360 3382.170 2372.790 ;
        RECT 3371.100 2300.070 3382.270 2322.500 ;
      LAYER met5 ;
        RECT 3370.100 486.470 3383.100 4958.900 ;
    END
  END vssd1
  PIN vssd1_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3489.900 2309.330 3557.160 2363.730 ;
    END
  END vssd1_pad
  PIN mprj_analog[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 924.720 4988.000 949.720 5070.350 ;
    END
  END mprj_analog[7]
  PIN mprj_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 907.050 5093.120 967.890 5153.945 ;
    END
  END mprj_io[21]
  PIN mprj_analog[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 667.720 4988.000 692.720 5070.350 ;
    END
  END mprj_analog[8]
  PIN mprj_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 650.050 5093.120 710.890 5153.945 ;
    END
  END mprj_io[22]
  PIN mprj_analog[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 410.720 4988.000 435.720 5070.350 ;
    END
  END mprj_analog[9]
  PIN mprj_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 393.050 5093.120 453.890 5153.945 ;
    END
  END mprj_io[23]
  PIN mprj_analog[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 117.650 4800.720 200.000 4825.720 ;
    END
  END mprj_analog[10]
  PIN mprj_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 34.055 4783.050 94.880 4843.890 ;
    END
  END mprj_io[24]
  PIN mprj_analog[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1465.390 4988.000 1537.000 5003.685 ;
    END
  END mprj_analog[5]
  PIN mprj_clamp_high[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1465.390 4988.000 1489.290 5013.660 ;
    END
  END mprj_clamp_high[1]
  PIN mprj_clamp_low[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1415.495 4988.000 1439.395 4990.055 ;
    END
  END mprj_clamp_low[1]
  PIN mprj_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1422.050 5093.120 1482.890 5153.945 ;
    END
  END mprj_io[19]
  PIN mprj_analog[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1202.390 4988.000 1274.000 5003.685 ;
    END
  END mprj_analog[6]
  PIN mprj_clamp_high[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.390 4988.000 1226.290 5013.660 ;
    END
  END mprj_clamp_high[2]
  PIN mprj_clamp_low[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1152.495 4988.000 1176.395 4990.055 ;
    END
  END mprj_clamp_low[2]
  PIN mprj_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1159.050 5093.120 1219.890 5153.945 ;
    END
  END mprj_io[20]
  PIN vccd2_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 30.835 4570.270 98.095 4624.670 ;
    END
  END vccd2_pad
  PIN vdda2_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 34.055 2422.050 94.880 2482.890 ;
    END
  END vdda2_pad
  PIN vssa2_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 34.055 4145.050 94.880 4205.890 ;
    END
  END vssa2_pad
  PIN vccd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 192.515 2277.730 197.965 2416.270 ;
    END
  END vccd
  PIN vccd2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 205.380 4610.755 236.020 4634.700 ;
        RECT 205.380 4560.500 236.020 4584.500 ;
        RECT 206.610 2230.000 236.030 2253.255 ;
      LAYER via3 ;
        RECT 223.390 4611.320 235.280 4634.080 ;
        RECT 223.480 4561.170 235.370 4583.930 ;
        RECT 223.360 2230.520 235.190 2252.670 ;
      LAYER met4 ;
        RECT 222.860 4610.830 235.850 4634.720 ;
        RECT 222.900 4560.590 235.890 4584.480 ;
        RECT 222.860 2230.050 235.890 2253.230 ;
      LAYER via4 ;
        RECT 223.390 4611.320 235.280 4634.080 ;
        RECT 223.480 4561.170 235.370 4583.930 ;
        RECT 223.360 2230.520 235.190 2252.670 ;
      LAYER met5 ;
        RECT 222.890 892.140 235.890 4871.190 ;
    END
  END vccd2
  PIN vdda2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 181.615 2278.035 185.065 2278.995 ;
    END
  END vdda2
  PIN vddio
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 164.665 2277.730 168.115 2416.270 ;
    END
  END vddio
  PIN vssa2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.265 2035.090 143.595 2628.610 ;
    END
  END vssa2
  PIN vssd2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 205.380 4585.950 235.820 4609.260 ;
        RECT 206.610 2254.755 236.030 2278.700 ;
        RECT 206.610 2204.500 236.030 2228.500 ;
      LAYER via3 ;
        RECT 207.420 4586.510 219.270 4608.610 ;
        RECT 207.450 2255.340 219.380 2278.140 ;
        RECT 207.410 2205.070 219.340 2227.870 ;
      LAYER met4 ;
        RECT 206.930 4586.050 219.920 4609.230 ;
        RECT 206.900 2254.740 219.830 2278.620 ;
        RECT 206.870 2204.570 219.800 2228.450 ;
      LAYER via4 ;
        RECT 207.420 4586.510 219.270 4608.610 ;
        RECT 207.450 2255.340 219.380 2278.140 ;
        RECT 207.410 2205.070 219.340 2227.870 ;
      LAYER met5 ;
        RECT 206.890 892.140 219.890 4871.190 ;
    END
  END vssd2
  PIN vssd2_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 30.835 2214.270 98.095 2268.670 ;
    END
  END vssd2_pad
  PIN vssio
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.035 2278.225 24.215 2280.465 ;
    END
  END vssio
  PIN flash_csb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1534.835 208.565 1535.115 210.965 ;
    END
  END flash_csb_core
  PIN flash_clk_ieb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.215 208.565 1787.495 210.965 ;
    END
  END flash_clk_ieb_core
  PIN flash_clk_oeb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1824.475 208.565 1824.755 210.965 ;
    END
  END flash_clk_oeb_core
  PIN flash_clk_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1808.835 208.565 1809.115 210.965 ;
    END
  END flash_clk_core
  PIN flash_csb_oeb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1550.475 208.565 1550.755 210.965 ;
    END
  END flash_csb_oeb_core
  PIN flash_csb_ieb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1513.215 208.565 1513.495 210.965 ;
    END
  END flash_csb_ieb_core
  OBS
      LAYER pwell ;
        RECT 1155.495 4988.935 1163.285 5011.790 ;
      LAYER nwell ;
        RECT 1163.860 4988.685 1222.965 4990.205 ;
      LAYER pwell ;
        RECT 1418.495 4988.935 1426.285 5011.790 ;
      LAYER nwell ;
        RECT 1426.860 4988.685 1485.965 4990.205 ;
        RECT 1678.860 4988.685 1737.965 4990.205 ;
      LAYER pwell ;
        RECT 1927.495 4988.935 1935.285 5011.790 ;
      LAYER nwell ;
        RECT 1935.860 4988.685 1994.965 4990.205 ;
        RECT 2889.860 4988.685 2948.965 4990.205 ;
        RECT 197.795 4360.860 199.315 4419.965 ;
      LAYER pwell ;
        RECT 176.210 4352.495 199.065 4360.285 ;
      LAYER nwell ;
        RECT 197.795 4149.860 199.315 4208.965 ;
      LAYER pwell ;
        RECT 3388.935 4155.715 3411.790 4163.505 ;
      LAYER nwell ;
        RECT 3388.685 4096.035 3390.205 4155.140 ;
      LAYER pwell ;
        RECT 3388.935 2582.715 3411.790 2590.505 ;
      LAYER nwell ;
        RECT 3388.685 2523.035 3390.205 2582.140 ;
        RECT 197.795 2426.860 199.315 2485.965 ;
      LAYER pwell ;
        RECT 176.210 2418.495 199.065 2426.285 ;
      LAYER nwell ;
        RECT 3388.685 2082.035 3390.205 2141.140 ;
        RECT 197.795 562.860 199.315 621.965 ;
      LAYER pwell ;
        RECT 176.210 554.495 199.065 562.285 ;
      LAYER nwell ;
        RECT 398.035 197.795 457.140 199.315 ;
        RECT 2849.035 197.795 2908.140 199.315 ;
        RECT 3118.035 197.795 3177.140 199.315 ;
      LAYER pwell ;
        RECT 3177.715 176.210 3185.505 199.065 ;
        RECT 679.530 103.265 738.130 103.270 ;
        RECT 662.870 102.005 738.130 103.265 ;
        RECT 662.870 100.770 666.070 102.005 ;
        RECT 679.530 100.770 738.130 102.005 ;
        RECT 662.870 97.475 738.130 100.770 ;
        RECT 662.870 75.865 664.440 97.475 ;
        RECT 736.565 75.865 738.130 97.475 ;
        RECT 662.870 70.685 738.130 75.865 ;
        RECT 662.870 69.645 676.090 70.685 ;
        RECT 696.250 69.645 738.130 70.685 ;
      LAYER nwell ;
        RECT 662.670 59.620 738.330 69.335 ;
      LAYER pwell ;
        RECT 662.710 55.435 738.290 59.315 ;
      LAYER nwell ;
        RECT 662.380 53.310 738.515 55.120 ;
        RECT 662.380 31.485 664.905 53.310 ;
        RECT 736.325 31.485 738.515 53.310 ;
        RECT 662.380 29.790 738.515 31.485 ;
      LAYER li1 ;
        RECT 388.905 5036.265 458.045 5169.100 ;
        RECT 645.905 5036.265 715.045 5169.100 ;
        RECT 902.905 5036.265 972.045 5169.100 ;
        RECT 1152.610 4990.035 1224.855 5187.695 ;
        RECT 1415.610 4990.035 1487.855 5187.695 ;
        RECT 1668.070 4990.035 1739.775 5187.695 ;
        RECT 1924.610 4990.035 1996.855 5187.695 ;
        RECT 2371.905 5036.265 2441.045 5169.100 ;
        RECT 2628.905 5036.265 2698.045 5169.100 ;
        RECT 2879.070 4990.035 2950.775 5187.695 ;
        RECT 3137.905 5036.265 3207.045 5169.100 ;
        RECT 1152.610 4989.065 1163.155 4990.035 ;
        RECT 1164.035 4989.920 1165.045 4990.035 ;
        RECT 1221.730 4989.920 1222.680 4990.035 ;
        RECT 1164.035 4988.970 1222.680 4989.920 ;
        RECT 1415.610 4989.065 1426.155 4990.035 ;
        RECT 1427.035 4989.920 1428.045 4990.035 ;
        RECT 1484.730 4989.920 1485.680 4990.035 ;
        RECT 1427.035 4988.970 1485.680 4989.920 ;
        RECT 1679.065 4989.890 1680.045 4990.035 ;
        RECT 1736.760 4989.890 1737.650 4990.035 ;
        RECT 1679.065 4989.000 1737.650 4989.890 ;
        RECT 1924.610 4989.065 1935.155 4990.035 ;
        RECT 1936.035 4989.920 1937.045 4990.035 ;
        RECT 1993.730 4989.920 1994.680 4990.035 ;
        RECT 1936.035 4988.970 1994.680 4989.920 ;
        RECT 2890.065 4989.890 2891.045 4990.035 ;
        RECT 2947.760 4989.890 2948.650 4990.035 ;
        RECT 2890.065 4989.000 2948.650 4989.890 ;
        RECT 18.900 4778.905 151.735 4848.045 ;
        RECT 3436.265 4760.955 3569.100 4830.095 ;
        RECT 0.305 4419.680 197.965 4421.855 ;
        RECT 0.305 4418.730 199.030 4419.680 ;
        RECT 0.305 4362.045 197.965 4418.730 ;
        RECT 198.080 4362.045 199.030 4418.730 ;
        RECT 0.305 4361.035 199.030 4362.045 ;
        RECT 0.305 4360.155 197.965 4361.035 ;
        RECT 0.305 4349.610 198.935 4360.155 ;
        RECT 3388.230 4311.840 3587.705 4392.160 ;
        RECT 0.305 4208.650 197.965 4210.775 ;
        RECT 0.305 4207.760 199.000 4208.650 ;
        RECT 0.305 4151.045 197.965 4207.760 ;
        RECT 198.110 4151.045 199.000 4207.760 ;
        RECT 3389.065 4155.845 3587.695 4166.390 ;
        RECT 3390.035 4154.965 3587.695 4155.845 ;
        RECT 0.305 4150.065 199.000 4151.045 ;
        RECT 3388.970 4153.955 3587.695 4154.965 ;
        RECT 0.305 4139.070 197.965 4150.065 ;
        RECT 3388.970 4097.270 3389.920 4153.955 ;
        RECT 3390.035 4097.270 3587.695 4153.955 ;
        RECT 3388.970 4096.320 3587.695 4097.270 ;
        RECT 3390.035 4094.145 3587.695 4096.320 ;
        RECT 0.295 3921.840 199.770 4002.160 ;
        RECT 3388.230 3865.840 3587.705 3946.160 ;
        RECT 0.295 3705.840 199.770 3786.160 ;
        RECT 3388.230 3640.840 3587.705 3721.160 ;
        RECT 0.295 3489.840 199.770 3570.160 ;
        RECT 3388.230 3415.840 3587.705 3496.160 ;
        RECT 0.295 3273.840 199.770 3354.160 ;
        RECT 3388.230 3189.840 3587.705 3270.160 ;
        RECT 0.295 3057.840 199.770 3138.160 ;
        RECT 3388.230 2964.840 3587.705 3045.160 ;
        RECT 0.295 2841.840 199.770 2922.160 ;
        RECT 3388.230 2738.840 3587.705 2819.160 ;
        RECT 0.295 2625.840 199.770 2706.160 ;
        RECT 3389.065 2582.845 3587.695 2593.390 ;
        RECT 3390.035 2581.965 3587.695 2582.845 ;
        RECT 3388.970 2580.955 3587.695 2581.965 ;
        RECT 3388.970 2524.270 3389.920 2580.955 ;
        RECT 3390.035 2524.270 3587.695 2580.955 ;
        RECT 3388.970 2523.320 3587.695 2524.270 ;
        RECT 3390.035 2521.145 3587.695 2523.320 ;
        RECT 0.305 2485.680 197.965 2487.855 ;
        RECT 0.305 2484.730 199.030 2485.680 ;
        RECT 0.305 2428.045 197.965 2484.730 ;
        RECT 198.080 2428.045 199.030 2484.730 ;
        RECT 0.305 2427.035 199.030 2428.045 ;
        RECT 0.305 2426.155 197.965 2427.035 ;
        RECT 0.305 2415.610 198.935 2426.155 ;
        RECT 3390.035 2140.935 3587.695 2151.930 ;
        RECT 3389.000 2139.955 3587.695 2140.935 ;
        RECT 3389.000 2083.240 3389.890 2139.955 ;
        RECT 3390.035 2083.240 3587.695 2139.955 ;
        RECT 3389.000 2082.350 3587.695 2083.240 ;
        RECT 3390.035 2080.225 3587.695 2082.350 ;
        RECT 0.295 1987.840 199.770 2068.160 ;
        RECT 3388.230 1852.840 3587.705 1933.160 ;
        RECT 0.295 1771.840 199.770 1852.160 ;
        RECT 0.295 1555.840 199.770 1636.160 ;
        RECT 3388.230 1626.840 3587.705 1707.160 ;
        RECT 0.295 1339.840 199.770 1420.160 ;
        RECT 3388.230 1401.840 3587.705 1482.160 ;
        RECT 0.295 1123.840 199.770 1204.160 ;
        RECT 3388.230 1176.840 3587.705 1257.160 ;
        RECT 0.295 907.840 199.770 988.160 ;
        RECT 3388.230 950.840 3587.705 1031.160 ;
        RECT 3388.230 725.840 3587.705 806.160 ;
        RECT 0.305 621.680 197.965 623.855 ;
        RECT 0.305 620.730 199.030 621.680 ;
        RECT 0.305 564.045 197.965 620.730 ;
        RECT 198.080 564.045 199.030 620.730 ;
        RECT 0.305 563.035 199.030 564.045 ;
        RECT 0.305 562.155 197.965 563.035 ;
        RECT 0.305 551.610 198.935 562.155 ;
        RECT 3388.230 499.840 3587.705 580.160 ;
        RECT 0.220 340.240 196.980 414.755 ;
        RECT 398.350 198.110 456.935 199.000 ;
        RECT 398.350 197.965 399.240 198.110 ;
        RECT 455.955 197.965 456.935 198.110 ;
        RECT 396.225 0.305 467.930 197.965 ;
        RECT 663.000 98.605 738.000 199.815 ;
        RECT 663.000 69.775 738.265 98.605 ;
        RECT 663.000 59.185 738.000 69.775 ;
        RECT 662.840 55.565 738.160 59.185 ;
        RECT 663.000 0.780 738.000 55.565 ;
        RECT 931.840 0.295 1012.160 199.770 ;
        RECT 1206.245 0.220 1280.760 196.980 ;
        RECT 1474.840 0.295 1555.160 199.770 ;
        RECT 1748.840 0.295 1829.160 199.770 ;
        RECT 2022.840 0.295 2103.160 199.770 ;
        RECT 2296.840 0.295 2377.160 199.770 ;
        RECT 2570.840 0.295 2651.160 199.770 ;
        RECT 2849.350 198.110 2907.935 199.000 ;
        RECT 2849.350 197.965 2850.240 198.110 ;
        RECT 2906.955 197.965 2907.935 198.110 ;
        RECT 3118.320 198.080 3176.965 199.030 ;
        RECT 3118.320 197.965 3119.270 198.080 ;
        RECT 3175.955 197.965 3176.965 198.080 ;
        RECT 3177.845 197.965 3188.390 198.935 ;
        RECT 2847.225 0.305 2918.930 197.965 ;
        RECT 3116.145 0.305 3188.390 197.965 ;
      LAYER met1 ;
        RECT 390.250 5034.255 456.440 5036.855 ;
        RECT 647.250 5034.255 713.440 5036.855 ;
        RECT 904.250 5034.255 970.440 5036.855 ;
        RECT 1152.185 4990.035 1224.915 5187.725 ;
        RECT 1415.185 4990.035 1487.915 5187.725 ;
        RECT 1667.185 4990.035 1740.620 5187.725 ;
        RECT 1924.185 4990.035 1996.915 5187.725 ;
        RECT 2373.250 5034.255 2439.440 5036.855 ;
        RECT 2630.250 5034.255 2696.440 5036.855 ;
        RECT 2878.185 4990.035 2951.620 5187.725 ;
        RECT 3139.250 5034.255 3205.440 5036.855 ;
        RECT 1155.625 4989.130 1160.855 4990.035 ;
        RECT 1164.035 4989.920 1165.350 4990.035 ;
        POLYGON 1165.350 4990.035 1165.465 4989.920 1165.350 4989.920 ;
        POLYGON 1221.540 4990.035 1221.540 4989.920 1221.425 4989.920 ;
        RECT 1221.540 4989.920 1222.680 4990.035 ;
        RECT 1164.035 4988.970 1222.680 4989.920 ;
        RECT 1418.625 4989.130 1423.855 4990.035 ;
        RECT 1427.035 4989.920 1428.350 4990.035 ;
        POLYGON 1428.350 4990.035 1428.465 4989.920 1428.350 4989.920 ;
        POLYGON 1484.540 4990.035 1484.540 4989.920 1484.425 4989.920 ;
        RECT 1484.540 4989.920 1485.680 4990.035 ;
        RECT 1427.035 4988.970 1485.680 4989.920 ;
        RECT 1679.035 4989.920 1680.350 4990.035 ;
        POLYGON 1680.350 4990.035 1680.465 4989.920 1680.350 4989.920 ;
        POLYGON 1736.540 4990.035 1736.540 4989.920 1736.425 4989.920 ;
        RECT 1736.540 4989.920 1737.680 4990.035 ;
        RECT 1679.035 4988.970 1737.680 4989.920 ;
        RECT 1927.625 4989.130 1932.855 4990.035 ;
        RECT 1936.035 4989.920 1937.350 4990.035 ;
        POLYGON 1937.350 4990.035 1937.465 4989.920 1937.350 4989.920 ;
        POLYGON 1993.540 4990.035 1993.540 4989.920 1993.425 4989.920 ;
        RECT 1993.540 4989.920 1994.680 4990.035 ;
        RECT 1936.035 4988.970 1994.680 4989.920 ;
        RECT 2890.035 4989.920 2891.350 4990.035 ;
        POLYGON 2891.350 4990.035 2891.465 4989.920 2891.350 4989.920 ;
        POLYGON 2947.540 4990.035 2947.540 4989.920 2947.425 4989.920 ;
        RECT 2947.540 4989.920 2948.680 4990.035 ;
        RECT 2890.035 4988.970 2948.680 4989.920 ;
        RECT 151.145 4780.250 153.745 4846.440 ;
        RECT 3434.255 4762.560 3436.855 4828.750 ;
        RECT 0.275 4419.680 197.965 4421.915 ;
        RECT 0.275 4418.540 199.030 4419.680 ;
        RECT 0.275 4362.350 197.965 4418.540 ;
        POLYGON 197.965 4418.540 198.080 4418.540 198.080 4418.425 ;
        POLYGON 198.080 4362.465 198.080 4362.350 197.965 4362.350 ;
        RECT 198.080 4362.350 199.030 4418.540 ;
      LAYER met1 ;
        RECT 3377.325 4375.335 3377.605 4375.365 ;
        RECT 3370.330 4375.055 3377.605 4375.335 ;
        RECT 3377.325 4375.025 3377.605 4375.055 ;
      LAYER met1 ;
        RECT 0.275 4361.035 199.030 4362.350 ;
        RECT 0.275 4357.855 197.965 4361.035 ;
      LAYER met1 ;
        RECT 3377.185 4360.155 3377.465 4360.185 ;
        RECT 3369.795 4359.875 3377.465 4360.155 ;
        RECT 3377.185 4359.845 3377.465 4359.875 ;
      LAYER met1 ;
        RECT 0.275 4352.625 198.870 4357.855 ;
      LAYER met1 ;
        RECT 3377.095 4353.715 3377.375 4353.745 ;
        RECT 3374.225 4353.435 3377.375 4353.715 ;
        RECT 3377.095 4353.405 3377.375 4353.435 ;
      LAYER met1 ;
        RECT 0.275 4349.185 197.965 4352.625 ;
      LAYER met1 ;
        RECT 3377.170 4322.895 3377.450 4322.925 ;
        RECT 3370.820 4322.615 3377.450 4322.895 ;
        RECT 3377.170 4322.585 3377.450 4322.615 ;
        RECT 3374.260 4313.415 3377.815 4313.675 ;
      LAYER met1 ;
        RECT 3381.155 4311.855 3588.000 4392.145 ;
        RECT 0.275 4208.680 197.965 4211.620 ;
        RECT 0.275 4207.540 199.030 4208.680 ;
        RECT 0.275 4151.350 197.965 4207.540 ;
        POLYGON 197.965 4207.540 198.080 4207.540 198.080 4207.425 ;
        POLYGON 198.080 4151.465 198.080 4151.350 197.965 4151.350 ;
        RECT 198.080 4151.350 199.030 4207.540 ;
        RECT 3390.035 4163.375 3587.725 4166.815 ;
        RECT 3389.130 4158.145 3587.725 4163.375 ;
        RECT 3390.035 4154.965 3587.725 4158.145 ;
        RECT 0.275 4150.035 199.030 4151.350 ;
        RECT 3388.970 4153.650 3587.725 4154.965 ;
        RECT 0.275 4138.185 197.965 4150.035 ;
        RECT 3388.970 4097.460 3389.920 4153.650 ;
        POLYGON 3389.920 4153.650 3390.035 4153.650 3389.920 4153.535 ;
        POLYGON 3389.920 4097.575 3390.035 4097.460 3389.920 4097.460 ;
        RECT 3390.035 4097.460 3587.725 4153.650 ;
        RECT 3388.970 4096.320 3587.725 4097.460 ;
        RECT 3390.035 4094.085 3587.725 4096.320 ;
        RECT 0.000 3921.855 206.845 4002.145 ;
      LAYER met1 ;
        RECT 210.340 4000.335 212.695 4000.615 ;
        RECT 210.340 3991.115 214.230 3991.395 ;
        RECT 210.340 3960.275 212.680 3960.555 ;
        RECT 210.340 3953.855 215.265 3954.135 ;
        RECT 210.340 3938.665 214.740 3938.945 ;
        RECT 3377.325 3929.335 3377.605 3929.365 ;
        RECT 3370.330 3929.055 3377.605 3929.335 ;
        RECT 3377.325 3929.025 3377.605 3929.055 ;
        RECT 3377.185 3914.155 3377.465 3914.185 ;
        RECT 3369.795 3913.875 3377.465 3914.155 ;
        RECT 3377.185 3913.845 3377.465 3913.875 ;
        RECT 3377.095 3907.715 3377.375 3907.745 ;
        RECT 3374.225 3907.435 3377.375 3907.715 ;
        RECT 3377.095 3907.405 3377.375 3907.435 ;
        RECT 3377.170 3876.895 3377.450 3876.925 ;
        RECT 3370.820 3876.615 3377.450 3876.895 ;
        RECT 3377.170 3876.585 3377.450 3876.615 ;
        RECT 3374.260 3867.415 3377.815 3867.675 ;
      LAYER met1 ;
        RECT 3381.155 3865.855 3588.000 3946.145 ;
        RECT 0.000 3705.855 206.845 3786.145 ;
      LAYER met1 ;
        RECT 209.725 3782.335 212.695 3782.615 ;
        RECT 210.340 3775.115 214.230 3775.395 ;
        RECT 210.340 3744.275 212.680 3744.555 ;
        RECT 210.340 3737.855 215.265 3738.135 ;
        RECT 210.340 3722.665 214.740 3722.945 ;
        RECT 3377.325 3704.335 3377.605 3704.365 ;
        RECT 3370.330 3704.055 3377.605 3704.335 ;
        RECT 3377.325 3704.025 3377.605 3704.055 ;
        RECT 3377.185 3689.155 3377.465 3689.185 ;
        RECT 3369.795 3688.875 3377.465 3689.155 ;
        RECT 3377.185 3688.845 3377.465 3688.875 ;
        RECT 3377.095 3682.715 3377.375 3682.745 ;
        RECT 3375.225 3682.435 3377.375 3682.715 ;
        RECT 3377.095 3682.405 3377.375 3682.435 ;
        RECT 3377.170 3651.895 3377.450 3651.925 ;
        RECT 3370.820 3651.615 3377.450 3651.895 ;
        RECT 3377.170 3651.585 3377.450 3651.615 ;
        RECT 3375.260 3642.415 3377.815 3642.675 ;
      LAYER met1 ;
        RECT 3381.155 3640.855 3588.000 3721.145 ;
      LAYER met1 ;
        RECT 210.655 3570.225 215.825 3570.505 ;
      LAYER met1 ;
        RECT 0.000 3489.855 206.845 3570.145 ;
      LAYER met1 ;
        RECT 210.340 3559.115 214.230 3559.395 ;
        RECT 210.340 3528.275 215.850 3528.555 ;
        RECT 210.340 3521.855 215.265 3522.135 ;
        RECT 210.340 3506.665 214.740 3506.945 ;
        RECT 3377.325 3479.335 3377.605 3479.365 ;
        RECT 3370.330 3479.055 3377.605 3479.335 ;
        RECT 3377.325 3479.025 3377.605 3479.055 ;
        RECT 3377.185 3464.155 3377.465 3464.185 ;
        RECT 3369.795 3463.875 3377.465 3464.155 ;
        RECT 3377.185 3463.845 3377.465 3463.875 ;
        RECT 3377.095 3457.715 3377.375 3457.745 ;
        RECT 3374.225 3457.435 3377.375 3457.715 ;
        RECT 3377.095 3457.405 3377.375 3457.435 ;
        RECT 3377.170 3426.895 3377.450 3426.925 ;
        RECT 3370.820 3426.615 3377.450 3426.895 ;
        RECT 3377.170 3426.585 3377.450 3426.615 ;
        RECT 3374.260 3417.415 3377.815 3417.675 ;
      LAYER met1 ;
        RECT 3381.155 3415.855 3588.000 3496.145 ;
        RECT 0.000 3273.855 206.845 3354.145 ;
      LAYER met1 ;
        RECT 209.815 3350.335 212.695 3350.615 ;
        RECT 210.340 3343.115 214.230 3343.395 ;
        RECT 210.340 3312.275 212.680 3312.555 ;
        RECT 210.340 3305.855 215.265 3306.135 ;
        RECT 210.340 3290.665 214.740 3290.945 ;
        RECT 3377.325 3253.335 3377.605 3253.365 ;
        RECT 3370.330 3253.055 3377.605 3253.335 ;
        RECT 3377.325 3253.025 3377.605 3253.055 ;
        RECT 3377.185 3238.155 3377.465 3238.185 ;
        RECT 3369.795 3237.875 3377.465 3238.155 ;
        RECT 3377.185 3237.845 3377.465 3237.875 ;
        RECT 3377.095 3231.715 3377.375 3231.745 ;
        RECT 3374.225 3231.435 3377.375 3231.715 ;
        RECT 3377.095 3231.405 3377.375 3231.435 ;
        RECT 3377.170 3200.895 3377.450 3200.925 ;
        RECT 3370.820 3200.615 3377.450 3200.895 ;
        RECT 3377.170 3200.585 3377.450 3200.615 ;
        RECT 3374.260 3191.415 3377.815 3191.675 ;
      LAYER met1 ;
        RECT 3381.155 3189.855 3588.000 3270.145 ;
        RECT 0.000 3057.855 206.845 3138.145 ;
      LAYER met1 ;
        RECT 210.340 3136.335 212.695 3136.615 ;
        RECT 210.340 3128.115 214.230 3128.395 ;
        RECT 210.340 3096.275 212.680 3096.555 ;
        RECT 210.340 3089.855 215.265 3090.135 ;
        RECT 210.340 3074.665 214.740 3074.945 ;
        RECT 3377.325 3028.335 3377.605 3028.365 ;
        RECT 3370.330 3028.055 3377.605 3028.335 ;
        RECT 3377.325 3028.025 3377.605 3028.055 ;
        RECT 3377.185 3013.155 3377.465 3013.185 ;
        RECT 3369.795 3012.875 3377.465 3013.155 ;
        RECT 3377.185 3012.845 3377.465 3012.875 ;
        RECT 3377.095 3006.715 3377.375 3006.745 ;
        RECT 3374.075 3006.435 3377.375 3006.715 ;
        RECT 3377.095 3006.405 3377.375 3006.435 ;
        RECT 3377.170 2975.895 3377.450 2975.925 ;
        RECT 3370.820 2975.615 3377.450 2975.895 ;
        RECT 3377.170 2975.585 3377.450 2975.615 ;
        RECT 3374.110 2966.415 3377.815 2966.675 ;
      LAYER met1 ;
        RECT 3381.155 2964.855 3588.000 3045.145 ;
        RECT 0.000 2841.855 206.845 2922.145 ;
      LAYER met1 ;
        RECT 210.340 2920.335 212.395 2920.615 ;
        RECT 210.495 2912.395 210.835 2912.410 ;
        RECT 210.490 2912.115 214.230 2912.395 ;
        RECT 210.340 2880.275 212.380 2880.555 ;
        RECT 210.340 2873.855 215.265 2874.135 ;
        RECT 210.340 2858.665 214.740 2858.945 ;
        RECT 3377.325 2802.335 3377.605 2802.365 ;
        RECT 3370.330 2802.055 3377.605 2802.335 ;
        RECT 3377.325 2802.025 3377.605 2802.055 ;
        RECT 3377.185 2787.155 3377.465 2787.185 ;
        RECT 3369.795 2786.875 3377.465 2787.155 ;
        RECT 3377.185 2786.845 3377.465 2786.875 ;
        RECT 3377.095 2780.715 3377.375 2780.745 ;
        RECT 3374.225 2780.435 3377.375 2780.715 ;
        RECT 3377.095 2780.405 3377.375 2780.435 ;
        RECT 3377.170 2749.895 3377.450 2749.925 ;
        RECT 3370.820 2749.615 3377.450 2749.895 ;
        RECT 3377.170 2749.585 3377.450 2749.615 ;
        RECT 3374.260 2740.415 3377.815 2740.675 ;
      LAYER met1 ;
        RECT 3381.155 2738.855 3588.000 2819.145 ;
        RECT 0.000 2625.855 206.845 2706.145 ;
      LAYER met1 ;
        RECT 210.340 2704.335 212.295 2704.615 ;
        RECT 210.340 2695.115 214.230 2695.395 ;
        RECT 210.340 2664.275 212.280 2664.555 ;
        RECT 210.340 2657.855 215.265 2658.135 ;
        RECT 210.340 2642.665 214.740 2642.945 ;
      LAYER met1 ;
        RECT 3390.035 2590.375 3587.725 2593.815 ;
        RECT 3389.130 2585.145 3587.725 2590.375 ;
        RECT 3390.035 2581.965 3587.725 2585.145 ;
        RECT 3388.970 2580.650 3587.725 2581.965 ;
        RECT 3388.970 2524.460 3389.920 2580.650 ;
        POLYGON 3389.920 2580.650 3390.035 2580.650 3389.920 2580.535 ;
        POLYGON 3389.920 2524.575 3390.035 2524.460 3389.920 2524.460 ;
        RECT 3390.035 2524.460 3587.725 2580.650 ;
        RECT 3388.970 2523.320 3587.725 2524.460 ;
        RECT 3390.035 2521.085 3587.725 2523.320 ;
        RECT 0.275 2485.680 197.965 2487.915 ;
        RECT 0.275 2484.540 199.030 2485.680 ;
        RECT 0.275 2428.350 197.965 2484.540 ;
        POLYGON 197.965 2484.540 198.080 2484.540 198.080 2484.425 ;
        POLYGON 198.080 2428.465 198.080 2428.350 197.965 2428.350 ;
        RECT 198.080 2428.350 199.030 2484.540 ;
        RECT 0.275 2427.035 199.030 2428.350 ;
        RECT 0.275 2423.855 197.965 2427.035 ;
        RECT 0.275 2418.625 198.870 2423.855 ;
        RECT 0.275 2415.185 197.965 2418.625 ;
        RECT 3390.035 2140.965 3587.725 2152.815 ;
        RECT 3388.970 2139.650 3587.725 2140.965 ;
        RECT 3388.970 2083.460 3389.920 2139.650 ;
        POLYGON 3389.920 2139.650 3390.035 2139.650 3389.920 2139.535 ;
        POLYGON 3389.920 2083.575 3390.035 2083.460 3389.920 2083.460 ;
        RECT 3390.035 2083.460 3587.725 2139.650 ;
        RECT 3388.970 2082.320 3587.725 2083.460 ;
        RECT 3390.035 2079.380 3587.725 2082.320 ;
        RECT 0.000 1987.855 206.845 2068.145 ;
      LAYER met1 ;
        RECT 210.340 2066.335 212.695 2066.615 ;
        RECT 210.340 2057.115 214.230 2057.395 ;
        RECT 210.340 2026.275 212.680 2026.555 ;
        RECT 210.340 2019.855 215.265 2020.135 ;
        RECT 210.340 2004.665 214.740 2004.945 ;
        RECT 3377.325 1916.335 3377.605 1916.365 ;
        RECT 3370.330 1916.055 3377.605 1916.335 ;
        RECT 3377.325 1916.025 3377.605 1916.055 ;
        RECT 3377.185 1901.155 3377.465 1901.185 ;
        RECT 3369.795 1900.875 3377.465 1901.155 ;
        RECT 3377.185 1900.845 3377.465 1900.875 ;
        RECT 3377.095 1894.715 3377.375 1894.745 ;
        RECT 3374.225 1894.435 3377.375 1894.715 ;
        RECT 3377.095 1894.405 3377.375 1894.435 ;
        RECT 3377.170 1863.895 3377.450 1863.925 ;
        RECT 3370.820 1863.615 3377.450 1863.895 ;
        RECT 3377.170 1863.585 3377.450 1863.615 ;
        RECT 3374.260 1854.415 3377.815 1854.675 ;
      LAYER met1 ;
        RECT 3381.155 1852.855 3588.000 1933.145 ;
        RECT 0.000 1771.855 206.845 1852.145 ;
      LAYER met1 ;
        RECT 210.340 1850.335 212.695 1850.615 ;
        RECT 210.340 1841.115 214.230 1841.395 ;
        RECT 210.340 1810.275 212.680 1810.555 ;
        RECT 210.340 1803.855 215.265 1804.135 ;
        RECT 210.340 1788.665 214.740 1788.945 ;
        RECT 3377.325 1690.335 3377.605 1690.365 ;
        RECT 3370.330 1690.055 3377.605 1690.335 ;
        RECT 3377.325 1690.025 3377.605 1690.055 ;
        RECT 3377.185 1675.155 3377.465 1675.185 ;
        RECT 3369.795 1674.875 3377.465 1675.155 ;
        RECT 3377.185 1674.845 3377.465 1674.875 ;
        RECT 3377.095 1668.715 3377.375 1668.745 ;
        RECT 3373.225 1668.435 3377.375 1668.715 ;
        RECT 3377.095 1668.405 3377.375 1668.435 ;
        RECT 3377.170 1637.895 3377.450 1637.925 ;
        RECT 3370.820 1637.615 3377.450 1637.895 ;
        RECT 3377.170 1637.585 3377.450 1637.615 ;
      LAYER met1 ;
        RECT 0.000 1555.855 206.845 1636.145 ;
      LAYER met1 ;
        RECT 210.340 1634.335 212.695 1634.615 ;
        RECT 3373.260 1628.415 3377.815 1628.675 ;
      LAYER met1 ;
        RECT 3381.155 1626.855 3588.000 1707.145 ;
      LAYER met1 ;
        RECT 210.340 1625.115 214.230 1625.395 ;
        RECT 210.340 1594.275 212.680 1594.555 ;
        RECT 210.340 1587.855 215.265 1588.135 ;
        RECT 210.340 1572.665 214.740 1572.945 ;
        RECT 3377.325 1465.335 3377.605 1465.365 ;
        RECT 3370.330 1465.055 3377.605 1465.335 ;
        RECT 3377.325 1465.025 3377.605 1465.055 ;
        RECT 3377.185 1450.155 3377.465 1450.185 ;
        RECT 3369.795 1449.875 3377.465 1450.155 ;
        RECT 3377.185 1449.845 3377.465 1449.875 ;
        RECT 3377.095 1443.715 3377.375 1443.745 ;
        RECT 3373.225 1443.435 3377.375 1443.715 ;
        RECT 3377.095 1443.405 3377.375 1443.435 ;
      LAYER met1 ;
        RECT 0.000 1339.855 206.845 1420.145 ;
      LAYER met1 ;
        RECT 210.340 1418.335 212.695 1418.615 ;
        RECT 3377.170 1412.895 3377.450 1412.925 ;
        RECT 3370.820 1412.615 3377.450 1412.895 ;
        RECT 3377.170 1412.585 3377.450 1412.615 ;
        RECT 210.340 1409.115 214.230 1409.395 ;
        RECT 3373.260 1403.415 3377.815 1403.675 ;
      LAYER met1 ;
        RECT 3381.155 1401.855 3588.000 1482.145 ;
      LAYER met1 ;
        RECT 210.340 1378.275 212.680 1378.555 ;
        RECT 210.340 1371.855 215.265 1372.135 ;
        RECT 210.340 1356.665 214.740 1356.945 ;
        RECT 3377.325 1240.335 3377.605 1240.365 ;
        RECT 3370.330 1240.055 3377.605 1240.335 ;
        RECT 3377.325 1240.025 3377.605 1240.055 ;
        RECT 3377.185 1225.155 3377.465 1225.185 ;
        RECT 3369.795 1224.875 3377.465 1225.155 ;
        RECT 3377.185 1224.845 3377.465 1224.875 ;
        RECT 3377.095 1218.715 3377.375 1218.745 ;
        RECT 3373.225 1218.435 3377.375 1218.715 ;
        RECT 3377.095 1218.405 3377.375 1218.435 ;
      LAYER met1 ;
        RECT 0.000 1123.855 206.845 1204.145 ;
      LAYER met1 ;
        RECT 210.340 1202.335 212.695 1202.615 ;
        RECT 210.340 1193.115 214.230 1193.395 ;
        RECT 3377.170 1187.895 3377.450 1187.925 ;
        RECT 3370.820 1187.615 3377.450 1187.895 ;
        RECT 3377.170 1187.585 3377.450 1187.615 ;
        RECT 3373.260 1178.415 3377.815 1178.675 ;
      LAYER met1 ;
        RECT 3381.155 1176.855 3588.000 1257.145 ;
      LAYER met1 ;
        RECT 210.340 1162.275 212.680 1162.555 ;
        RECT 210.340 1155.855 215.265 1156.135 ;
        RECT 210.340 1140.665 214.740 1140.945 ;
        RECT 3377.325 1014.335 3377.605 1014.365 ;
        RECT 3370.330 1014.055 3377.605 1014.335 ;
        RECT 3377.325 1014.025 3377.605 1014.055 ;
        RECT 3377.185 999.155 3377.465 999.185 ;
        RECT 3369.795 998.875 3377.465 999.155 ;
        RECT 3377.185 998.845 3377.465 998.875 ;
        RECT 3377.095 992.715 3377.375 992.745 ;
        RECT 3373.225 992.435 3377.375 992.715 ;
        RECT 3377.095 992.405 3377.375 992.435 ;
      LAYER met1 ;
        RECT 0.000 907.855 206.845 988.145 ;
      LAYER met1 ;
        RECT 210.340 986.335 212.695 986.615 ;
        RECT 210.340 977.115 214.230 977.395 ;
        RECT 3377.170 961.895 3377.450 961.925 ;
        RECT 3370.820 961.615 3377.450 961.895 ;
        RECT 3377.170 961.585 3377.450 961.615 ;
        RECT 3373.260 952.415 3377.815 952.675 ;
      LAYER met1 ;
        RECT 3381.155 950.855 3588.000 1031.145 ;
      LAYER met1 ;
        RECT 210.340 946.275 212.680 946.555 ;
        RECT 210.340 939.855 215.265 940.135 ;
        RECT 210.340 924.665 214.740 924.945 ;
        RECT 213.920 905.395 214.240 905.400 ;
        RECT 208.120 905.145 214.285 905.395 ;
        RECT 208.120 888.515 208.370 905.145 ;
        RECT 213.920 905.140 214.240 905.145 ;
        RECT 214.430 904.895 214.750 904.900 ;
        RECT 208.620 904.645 214.830 904.895 ;
        RECT 208.620 889.015 208.870 904.645 ;
        RECT 214.430 904.640 214.750 904.645 ;
        RECT 214.920 904.395 215.240 904.400 ;
        RECT 209.120 904.145 215.315 904.395 ;
        RECT 209.120 889.515 209.370 904.145 ;
        RECT 214.920 904.140 215.240 904.145 ;
        RECT 209.120 889.265 212.370 889.515 ;
        RECT 208.620 888.765 211.870 889.015 ;
        RECT 208.120 888.265 211.370 888.515 ;
      LAYER met1 ;
        RECT 0.275 621.680 197.965 623.915 ;
        RECT 0.275 620.540 199.030 621.680 ;
        RECT 0.275 564.350 197.965 620.540 ;
        POLYGON 197.965 620.540 198.080 620.540 198.080 620.425 ;
        POLYGON 198.080 564.465 198.080 564.350 197.965 564.350 ;
        RECT 198.080 564.350 199.030 620.540 ;
        RECT 0.275 563.035 199.030 564.350 ;
        RECT 0.275 559.855 197.965 563.035 ;
        RECT 0.275 554.625 198.870 559.855 ;
        RECT 0.275 551.185 197.965 554.625 ;
        RECT 159.640 425.935 163.510 426.195 ;
        RECT 159.640 421.935 204.500 425.935 ;
        POLYGON 204.500 425.935 208.500 421.935 204.500 421.935 ;
        RECT 159.640 416.200 208.500 421.935 ;
        RECT 159.640 415.245 163.510 416.200 ;
        RECT 0.160 396.565 197.965 415.000 ;
        RECT 198.780 396.565 208.500 416.200 ;
        RECT 0.160 360.495 208.500 396.565 ;
        RECT 0.160 356.655 198.000 360.495 ;
        RECT 198.980 358.655 208.500 360.495 ;
        POLYGON 198.980 358.655 200.980 358.655 200.980 356.655 ;
        RECT 200.980 356.655 206.500 358.655 ;
        POLYGON 206.500 358.655 208.500 358.655 206.500 356.655 ;
        RECT 0.160 340.120 197.965 356.655 ;
      LAYER met1 ;
        RECT 211.120 349.935 211.370 888.265 ;
        RECT 211.050 347.125 211.480 349.935 ;
        RECT 211.120 210.670 211.370 347.125 ;
        RECT 211.620 212.750 211.870 888.765 ;
        RECT 212.120 563.775 212.370 889.265 ;
        RECT 3377.325 789.335 3377.605 789.365 ;
        RECT 3370.330 789.055 3377.605 789.335 ;
        RECT 3377.325 789.025 3377.605 789.055 ;
        RECT 3377.185 774.155 3377.465 774.185 ;
        RECT 3369.795 773.875 3377.465 774.155 ;
        RECT 3377.185 773.845 3377.465 773.875 ;
        RECT 3377.095 767.715 3377.375 767.745 ;
        RECT 3373.225 767.435 3377.375 767.715 ;
        RECT 3377.095 767.405 3377.375 767.435 ;
        RECT 3377.170 736.895 3377.450 736.925 ;
        RECT 3370.820 736.615 3377.450 736.895 ;
        RECT 3377.170 736.585 3377.450 736.615 ;
        RECT 3373.260 727.415 3377.815 727.675 ;
      LAYER met1 ;
        RECT 3381.155 725.855 3588.000 806.145 ;
      LAYER met1 ;
        RECT 212.070 561.770 212.595 563.775 ;
        RECT 3377.325 563.335 3377.605 563.365 ;
        RECT 3370.330 563.055 3377.605 563.335 ;
        RECT 3377.325 563.025 3377.605 563.055 ;
        RECT 211.605 212.030 211.870 212.750 ;
        RECT 211.620 211.975 211.870 212.030 ;
        RECT 212.120 211.670 212.370 561.770 ;
        RECT 3377.185 548.155 3377.465 548.185 ;
        RECT 3369.795 547.875 3377.465 548.155 ;
        RECT 3377.185 547.845 3377.465 547.875 ;
        RECT 3377.095 541.715 3377.375 541.745 ;
        RECT 3373.225 541.435 3377.375 541.715 ;
        RECT 3377.095 541.405 3377.375 541.435 ;
        RECT 3377.170 510.895 3377.450 510.925 ;
        RECT 3370.820 510.615 3377.450 510.895 ;
        RECT 3377.170 510.585 3377.450 510.615 ;
        RECT 3373.260 501.415 3377.815 501.675 ;
      LAYER met1 ;
        RECT 3381.155 499.855 3588.000 580.145 ;
      LAYER met1 ;
        RECT 2856.605 213.185 2858.820 214.920 ;
        RECT 2529.510 212.925 3370.645 213.185 ;
        RECT 1476.400 212.750 1476.720 212.775 ;
        RECT 1516.420 212.750 1516.740 212.775 ;
        RECT 1750.400 212.750 1750.720 212.775 ;
        RECT 1790.420 212.750 1790.740 212.775 ;
        RECT 2024.400 212.750 2024.720 212.775 ;
        RECT 2064.420 212.750 2064.740 212.775 ;
        RECT 1476.380 212.540 1516.740 212.750 ;
        RECT 1750.380 212.540 1790.740 212.750 ;
        RECT 2024.380 212.540 2064.740 212.750 ;
        RECT 1476.400 212.515 1476.720 212.540 ;
        RECT 1516.420 212.515 1516.740 212.540 ;
        RECT 1750.400 212.515 1750.720 212.540 ;
        RECT 1790.420 212.515 1790.740 212.540 ;
        RECT 2024.400 212.515 2024.720 212.540 ;
        RECT 2064.420 212.515 2064.740 212.540 ;
        RECT 2529.510 212.320 2529.770 212.925 ;
        RECT 2856.605 212.915 2858.820 212.925 ;
        RECT 2618.880 212.540 2619.200 212.545 ;
        RECT 3369.800 212.540 3370.120 212.545 ;
        RECT 212.635 212.060 2529.770 212.320 ;
        RECT 2530.420 212.290 3370.180 212.540 ;
        RECT 979.880 211.670 980.200 211.675 ;
        RECT 1522.880 211.670 1523.200 211.675 ;
        RECT 1796.880 211.670 1797.200 211.675 ;
        RECT 2070.880 211.670 2071.200 211.675 ;
        RECT 2344.880 211.670 2345.200 211.675 ;
        RECT 2530.420 211.670 2530.670 212.290 ;
        RECT 2618.880 212.285 2619.200 212.290 ;
        RECT 3369.800 212.285 3370.120 212.290 ;
        RECT 2634.050 212.040 2634.370 212.045 ;
        RECT 212.120 211.420 2530.670 211.670 ;
        RECT 2530.920 211.790 2634.440 212.040 ;
        RECT 979.880 211.415 980.200 211.420 ;
        RECT 1522.880 211.415 1523.200 211.420 ;
        RECT 1796.880 211.415 1797.200 211.420 ;
        RECT 2070.880 211.415 2071.200 211.420 ;
        RECT 2344.880 211.415 2345.200 211.420 ;
        RECT 454.315 211.170 455.470 211.225 ;
        RECT 995.080 211.170 995.400 211.175 ;
        RECT 1538.050 211.170 1538.370 211.175 ;
        RECT 1812.050 211.170 1812.370 211.175 ;
        RECT 2086.050 211.170 2086.370 211.175 ;
        RECT 2360.050 211.170 2360.370 211.175 ;
        RECT 2530.920 211.170 2531.170 211.790 ;
        RECT 2634.050 211.785 2634.370 211.790 ;
        RECT 2581.600 211.540 2581.920 211.545 ;
        RECT 3370.800 211.540 3371.120 211.545 ;
        RECT 454.230 210.920 2531.170 211.170 ;
        RECT 2531.420 211.290 3371.160 211.540 ;
        RECT 454.315 210.870 455.470 210.920 ;
        RECT 995.080 210.915 995.400 210.920 ;
        RECT 1538.050 210.915 1538.370 210.920 ;
        RECT 1812.050 210.915 1812.370 210.920 ;
        RECT 2086.050 210.915 2086.370 210.920 ;
        RECT 2360.050 210.915 2360.370 210.920 ;
        RECT 729.235 210.670 729.565 210.680 ;
        RECT 942.600 210.670 942.920 210.675 ;
        RECT 964.200 210.670 964.520 210.675 ;
        RECT 1007.430 210.670 1007.750 210.675 ;
        RECT 1485.600 210.670 1485.920 210.675 ;
        RECT 1759.600 210.670 1759.920 210.675 ;
        RECT 1802.825 210.670 1803.165 210.695 ;
        RECT 2033.600 210.670 2033.920 210.675 ;
        RECT 2307.600 210.670 2307.920 210.675 ;
        RECT 2531.420 210.670 2531.670 211.290 ;
        RECT 2581.600 211.285 2581.920 211.290 ;
        RECT 3370.800 211.285 3371.120 211.290 ;
        RECT 2584.810 211.040 2585.130 211.045 ;
        RECT 2599.970 211.040 2600.290 211.045 ;
        RECT 2606.470 211.040 2606.790 211.045 ;
        RECT 2621.590 211.040 2621.910 211.045 ;
        RECT 2628.050 211.040 2628.370 211.045 ;
        RECT 2640.040 211.040 2640.360 211.045 ;
        RECT 2643.230 211.040 2643.550 211.045 ;
        RECT 211.120 210.420 2531.670 210.670 ;
        RECT 2531.920 210.790 2643.680 211.040 ;
        RECT 729.235 210.410 729.565 210.420 ;
        RECT 942.600 210.415 942.920 210.420 ;
        RECT 964.200 210.415 964.520 210.420 ;
        RECT 1007.430 210.415 1007.750 210.420 ;
        RECT 1485.600 210.415 1485.920 210.420 ;
        RECT 1498.005 210.380 1498.345 210.420 ;
        RECT 1528.825 210.370 1529.165 210.420 ;
        RECT 1759.600 210.415 1759.920 210.420 ;
        RECT 1772.005 210.390 1772.345 210.420 ;
        RECT 1802.825 210.415 1803.165 210.420 ;
        RECT 2033.600 210.415 2033.920 210.420 ;
        RECT 2307.600 210.415 2307.920 210.420 ;
        RECT 945.810 210.170 946.130 210.175 ;
        RECT 955.020 210.170 955.340 210.175 ;
        RECT 960.970 210.170 961.290 210.175 ;
        RECT 967.470 210.170 967.790 210.175 ;
        RECT 982.590 210.170 982.910 210.175 ;
        RECT 985.850 210.170 986.170 210.175 ;
        RECT 989.050 210.170 989.370 210.175 ;
        RECT 991.840 210.170 992.160 210.175 ;
        RECT 1001.040 210.170 1001.360 210.175 ;
        RECT 1004.230 210.170 1004.550 210.175 ;
        RECT 1268.065 210.170 1269.135 210.215 ;
        RECT 1488.810 210.170 1489.130 210.175 ;
        RECT 1503.970 210.170 1504.290 210.175 ;
        RECT 1510.470 210.170 1510.790 210.175 ;
        RECT 1525.590 210.170 1525.910 210.175 ;
        RECT 1532.050 210.170 1532.370 210.175 ;
        RECT 1544.040 210.170 1544.360 210.175 ;
        RECT 1547.230 210.170 1547.550 210.175 ;
        RECT 1762.810 210.170 1763.130 210.175 ;
        RECT 1777.970 210.170 1778.290 210.175 ;
        RECT 1784.470 210.170 1784.790 210.175 ;
        RECT 1799.590 210.170 1799.910 210.175 ;
        RECT 1806.050 210.170 1806.370 210.175 ;
        RECT 1818.040 210.170 1818.360 210.175 ;
        RECT 1821.230 210.170 1821.550 210.175 ;
        RECT 2036.810 210.170 2037.130 210.175 ;
        RECT 2051.970 210.170 2052.290 210.175 ;
        RECT 2058.470 210.170 2058.790 210.175 ;
        RECT 2073.590 210.170 2073.910 210.175 ;
        RECT 2080.050 210.170 2080.370 210.175 ;
        RECT 2092.040 210.170 2092.360 210.175 ;
        RECT 2095.230 210.170 2095.550 210.175 ;
        RECT 2310.810 210.170 2311.130 210.175 ;
        RECT 2325.970 210.170 2326.290 210.175 ;
        RECT 2332.470 210.170 2332.790 210.175 ;
        RECT 2347.590 210.170 2347.910 210.175 ;
        RECT 2354.050 210.170 2354.370 210.175 ;
        RECT 2366.040 210.170 2366.360 210.175 ;
        RECT 2369.230 210.170 2369.550 210.175 ;
        RECT 2531.920 210.170 2532.170 210.790 ;
        RECT 2584.810 210.785 2585.130 210.790 ;
        RECT 2599.970 210.785 2600.290 210.790 ;
        RECT 2606.470 210.785 2606.790 210.790 ;
        RECT 2621.590 210.785 2621.910 210.790 ;
        RECT 2628.050 210.785 2628.370 210.790 ;
        RECT 2640.040 210.785 2640.360 210.790 ;
        RECT 2643.230 210.785 2643.550 210.790 ;
        RECT 2572.400 210.570 2572.720 210.595 ;
        RECT 2612.420 210.570 2612.740 210.595 ;
        RECT 2572.380 210.360 2612.740 210.570 ;
        RECT 2572.400 210.335 2572.720 210.360 ;
        RECT 2612.420 210.335 2612.740 210.360 ;
        RECT 945.800 209.920 2532.170 210.170 ;
        RECT 945.810 209.915 946.130 209.920 ;
        RECT 955.020 209.915 955.340 209.920 ;
        RECT 960.970 209.915 961.290 209.920 ;
        RECT 967.470 209.915 967.790 209.920 ;
        RECT 982.590 209.915 982.910 209.920 ;
        RECT 985.850 209.915 986.170 209.920 ;
        RECT 989.050 209.915 989.370 209.920 ;
        RECT 991.840 209.915 992.160 209.920 ;
        RECT 1001.040 209.915 1001.360 209.920 ;
        RECT 1004.230 209.915 1004.550 209.920 ;
        RECT 1268.065 209.755 1269.135 209.920 ;
        RECT 1488.810 209.915 1489.130 209.920 ;
        RECT 1503.970 209.915 1504.290 209.920 ;
        RECT 1507.205 209.885 1507.545 209.920 ;
        RECT 1510.470 209.915 1510.790 209.920 ;
        RECT 1525.590 209.915 1525.910 209.920 ;
        RECT 1532.050 209.915 1532.370 209.920 ;
        RECT 1544.040 209.915 1544.360 209.920 ;
        RECT 1547.230 209.915 1547.550 209.920 ;
        RECT 1762.810 209.915 1763.130 209.920 ;
        RECT 1777.970 209.915 1778.290 209.920 ;
        RECT 1781.205 209.870 1781.545 209.920 ;
        RECT 1784.470 209.915 1784.790 209.920 ;
        RECT 1799.590 209.915 1799.910 209.920 ;
        RECT 1806.050 209.915 1806.370 209.920 ;
        RECT 1818.040 209.915 1818.360 209.920 ;
        RECT 1821.230 209.915 1821.550 209.920 ;
        RECT 2036.810 209.915 2037.130 209.920 ;
        RECT 2051.970 209.915 2052.290 209.920 ;
        RECT 2058.470 209.915 2058.790 209.920 ;
        RECT 2073.590 209.915 2073.910 209.920 ;
        RECT 2080.050 209.915 2080.370 209.920 ;
        RECT 2092.040 209.915 2092.360 209.920 ;
        RECT 2095.230 209.915 2095.550 209.920 ;
        RECT 2310.810 209.915 2311.130 209.920 ;
        RECT 2325.970 209.915 2326.290 209.920 ;
        RECT 2332.470 209.915 2332.790 209.920 ;
        RECT 2347.590 209.915 2347.910 209.920 ;
        RECT 2354.050 209.915 2354.370 209.920 ;
        RECT 2366.040 209.915 2366.360 209.920 ;
        RECT 2369.230 209.915 2369.550 209.920 ;
        RECT 933.400 209.700 933.720 209.725 ;
        RECT 973.420 209.700 973.740 209.725 ;
        RECT 2298.400 209.700 2298.720 209.725 ;
        RECT 2338.420 209.700 2338.740 209.725 ;
        RECT 933.380 209.490 973.740 209.700 ;
        RECT 2298.380 209.490 2338.740 209.700 ;
        RECT 933.400 209.465 933.720 209.490 ;
        RECT 973.420 209.465 973.740 209.490 ;
        RECT 2298.400 209.465 2298.720 209.490 ;
        RECT 2338.420 209.465 2338.740 209.490 ;
      LAYER met1 ;
        POLYGON 1199.065 208.500 1199.065 206.845 1197.410 206.845 ;
        RECT 1199.065 206.845 1262.345 208.500 ;
      LAYER met1 ;
        RECT 664.960 201.105 665.280 201.140 ;
        RECT 719.595 201.105 719.915 201.140 ;
        RECT 664.960 200.915 719.915 201.105 ;
        RECT 664.960 200.880 665.280 200.915 ;
        RECT 719.595 200.880 719.915 200.915 ;
        RECT 712.850 200.320 713.110 200.640 ;
      LAYER met1 ;
        RECT 663.000 199.390 704.700 199.815 ;
      LAYER met1 ;
        RECT 704.980 199.670 705.240 200.000 ;
      LAYER met1 ;
        RECT 705.520 199.390 706.565 199.815 ;
      LAYER met1 ;
        RECT 706.845 199.670 707.495 200.000 ;
      LAYER met1 ;
        RECT 707.775 199.390 709.490 199.815 ;
      LAYER met1 ;
        RECT 709.770 199.670 710.420 200.000 ;
      LAYER met1 ;
        RECT 710.700 199.390 712.585 199.815 ;
        RECT 398.320 198.080 456.965 199.030 ;
        RECT 398.320 197.965 399.460 198.080 ;
        POLYGON 399.460 198.080 399.575 198.080 399.460 197.965 ;
        POLYGON 455.535 198.080 455.650 198.080 455.650 197.965 ;
        RECT 455.650 197.965 456.965 198.080 ;
        RECT 395.380 0.275 468.815 197.965 ;
        RECT 663.000 189.745 712.585 199.390 ;
      LAYER met1 ;
        RECT 712.865 190.025 713.095 200.320 ;
      LAYER met1 ;
        RECT 713.375 199.390 715.060 199.815 ;
      LAYER met1 ;
        RECT 715.340 199.670 715.640 200.000 ;
      LAYER met1 ;
        RECT 715.920 199.390 722.585 199.815 ;
      LAYER met1 ;
        RECT 722.865 199.670 723.445 200.000 ;
      LAYER met1 ;
        RECT 723.725 199.390 725.175 199.815 ;
      LAYER met1 ;
        RECT 725.455 199.670 725.715 200.000 ;
      LAYER met1 ;
        RECT 725.995 199.390 738.000 199.815 ;
        RECT 713.375 189.745 738.000 199.390 ;
        RECT 663.000 104.105 738.000 189.745 ;
        RECT 662.855 69.780 738.145 104.105 ;
        RECT 663.000 68.725 738.000 69.780 ;
        RECT 662.855 29.910 738.145 68.725 ;
        RECT 663.000 0.790 738.000 29.910 ;
        RECT 931.855 0.000 1012.145 206.845 ;
        POLYGON 1197.410 206.845 1197.410 204.500 1195.065 204.500 ;
        RECT 1197.410 206.500 1262.345 206.845 ;
        POLYGON 1262.345 208.500 1264.345 206.500 1262.345 206.500 ;
        RECT 1197.410 204.500 1264.345 206.500 ;
        RECT 1195.065 200.980 1264.345 204.500 ;
        RECT 1195.065 198.980 1262.345 200.980 ;
        POLYGON 1262.345 200.980 1264.345 200.980 1262.345 198.980 ;
        RECT 1195.065 198.780 1260.505 198.980 ;
        RECT 1195.065 163.510 1204.800 198.780 ;
        RECT 1224.435 198.000 1260.505 198.780 ;
        RECT 1224.435 197.965 1264.345 198.000 ;
        RECT 1194.805 159.640 1205.755 163.510 ;
        RECT 1206.000 0.160 1280.880 197.965 ;
        RECT 1474.855 0.000 1555.145 206.845 ;
        RECT 1748.855 0.000 1829.145 206.845 ;
        RECT 2022.855 0.000 2103.145 206.845 ;
        RECT 2296.855 0.000 2377.145 206.845 ;
        RECT 2570.855 0.000 2651.145 206.845 ;
        RECT 2849.320 198.080 2907.965 199.030 ;
        RECT 2849.320 197.965 2850.460 198.080 ;
        POLYGON 2850.460 198.080 2850.575 198.080 2850.460 197.965 ;
        POLYGON 2906.535 198.080 2906.650 198.080 2906.650 197.965 ;
        RECT 2906.650 197.965 2907.965 198.080 ;
        RECT 3118.320 198.080 3176.965 199.030 ;
        RECT 3118.320 197.965 3119.460 198.080 ;
        POLYGON 3119.460 198.080 3119.575 198.080 3119.460 197.965 ;
        POLYGON 3175.535 198.080 3175.650 198.080 3175.650 197.965 ;
        RECT 3175.650 197.965 3176.965 198.080 ;
        RECT 3180.145 197.965 3185.375 198.870 ;
        RECT 2846.380 0.275 2919.815 197.965 ;
        RECT 3116.085 0.275 3188.815 197.965 ;
      LAYER via ;
        RECT 3370.360 4375.055 3370.640 4375.335 ;
        RECT 3377.325 4375.055 3377.605 4375.335 ;
        RECT 3369.825 4359.875 3370.105 4360.155 ;
        RECT 3377.185 4359.875 3377.465 4360.155 ;
        RECT 3374.255 4353.435 3374.535 4353.715 ;
        RECT 3377.095 4353.435 3377.375 4353.715 ;
        RECT 3370.850 4322.615 3371.130 4322.895 ;
        RECT 3377.170 4322.615 3377.450 4322.895 ;
        RECT 3374.290 4313.415 3374.550 4313.675 ;
        RECT 3377.525 4313.415 3377.785 4313.675 ;
        RECT 210.370 4000.335 210.650 4000.615 ;
        RECT 212.385 4000.335 212.665 4000.615 ;
        RECT 210.370 3991.115 210.650 3991.395 ;
        RECT 213.920 3991.115 214.200 3991.395 ;
        RECT 210.370 3960.275 210.650 3960.555 ;
        RECT 212.370 3960.275 212.650 3960.555 ;
        RECT 210.370 3953.855 210.650 3954.135 ;
        RECT 214.955 3953.855 215.235 3954.135 ;
        RECT 210.370 3938.665 210.650 3938.945 ;
        RECT 214.430 3938.665 214.710 3938.945 ;
        RECT 3370.360 3929.055 3370.640 3929.335 ;
        RECT 3377.325 3929.055 3377.605 3929.335 ;
        RECT 3369.825 3913.875 3370.105 3914.155 ;
        RECT 3377.185 3913.875 3377.465 3914.155 ;
        RECT 3374.255 3907.435 3374.535 3907.715 ;
        RECT 3377.095 3907.435 3377.375 3907.715 ;
        RECT 3370.850 3876.615 3371.130 3876.895 ;
        RECT 3377.170 3876.615 3377.450 3876.895 ;
        RECT 3374.290 3867.415 3374.550 3867.675 ;
        RECT 3377.525 3867.415 3377.785 3867.675 ;
        RECT 209.755 3782.335 210.035 3782.615 ;
        RECT 212.385 3782.335 212.665 3782.615 ;
        RECT 210.370 3775.115 210.650 3775.395 ;
        RECT 213.920 3775.115 214.200 3775.395 ;
        RECT 210.370 3744.275 210.650 3744.555 ;
        RECT 212.370 3744.275 212.650 3744.555 ;
        RECT 210.370 3737.855 210.650 3738.135 ;
        RECT 214.955 3737.855 215.235 3738.135 ;
        RECT 210.370 3722.665 210.650 3722.945 ;
        RECT 214.430 3722.665 214.710 3722.945 ;
        RECT 3370.360 3704.055 3370.640 3704.335 ;
        RECT 3377.325 3704.055 3377.605 3704.335 ;
        RECT 3369.825 3688.875 3370.105 3689.155 ;
        RECT 3377.185 3688.875 3377.465 3689.155 ;
        RECT 3375.255 3682.435 3375.535 3682.715 ;
        RECT 3377.095 3682.435 3377.375 3682.715 ;
        RECT 3370.850 3651.615 3371.130 3651.895 ;
        RECT 3377.170 3651.615 3377.450 3651.895 ;
        RECT 3375.290 3642.415 3375.550 3642.675 ;
        RECT 3377.525 3642.415 3377.785 3642.675 ;
        RECT 210.685 3570.225 210.965 3570.505 ;
        RECT 215.515 3570.225 215.795 3570.505 ;
        RECT 210.370 3559.115 210.650 3559.395 ;
        RECT 213.920 3559.115 214.200 3559.395 ;
        RECT 210.370 3528.275 210.650 3528.555 ;
        RECT 215.540 3528.275 215.820 3528.555 ;
        RECT 210.370 3521.855 210.650 3522.135 ;
        RECT 214.955 3521.855 215.235 3522.135 ;
        RECT 210.370 3506.665 210.650 3506.945 ;
        RECT 214.430 3506.665 214.710 3506.945 ;
        RECT 3370.360 3479.055 3370.640 3479.335 ;
        RECT 3377.325 3479.055 3377.605 3479.335 ;
        RECT 3369.825 3463.875 3370.105 3464.155 ;
        RECT 3377.185 3463.875 3377.465 3464.155 ;
        RECT 3374.255 3457.435 3374.535 3457.715 ;
        RECT 3377.095 3457.435 3377.375 3457.715 ;
        RECT 3370.850 3426.615 3371.130 3426.895 ;
        RECT 3377.170 3426.615 3377.450 3426.895 ;
        RECT 3374.290 3417.415 3374.550 3417.675 ;
        RECT 3377.525 3417.415 3377.785 3417.675 ;
        RECT 209.845 3350.335 210.125 3350.615 ;
        RECT 212.385 3350.335 212.665 3350.615 ;
        RECT 210.370 3343.115 210.650 3343.395 ;
        RECT 213.920 3343.115 214.200 3343.395 ;
        RECT 210.370 3312.275 210.650 3312.555 ;
        RECT 212.370 3312.275 212.650 3312.555 ;
        RECT 210.370 3305.855 210.650 3306.135 ;
        RECT 214.955 3305.855 215.235 3306.135 ;
        RECT 210.370 3290.665 210.650 3290.945 ;
        RECT 214.430 3290.665 214.710 3290.945 ;
        RECT 3370.360 3253.055 3370.640 3253.335 ;
        RECT 3377.325 3253.055 3377.605 3253.335 ;
        RECT 3369.825 3237.875 3370.105 3238.155 ;
        RECT 3377.185 3237.875 3377.465 3238.155 ;
        RECT 3374.255 3231.435 3374.535 3231.715 ;
        RECT 3377.095 3231.435 3377.375 3231.715 ;
        RECT 3370.850 3200.615 3371.130 3200.895 ;
        RECT 3377.170 3200.615 3377.450 3200.895 ;
        RECT 3374.290 3191.415 3374.550 3191.675 ;
        RECT 3377.525 3191.415 3377.785 3191.675 ;
        RECT 210.370 3136.335 210.650 3136.615 ;
        RECT 212.385 3136.335 212.665 3136.615 ;
        RECT 210.370 3128.115 210.650 3128.395 ;
        RECT 213.920 3128.115 214.200 3128.395 ;
        RECT 210.370 3096.275 210.650 3096.555 ;
        RECT 212.370 3096.275 212.650 3096.555 ;
        RECT 210.370 3089.855 210.650 3090.135 ;
        RECT 214.955 3089.855 215.235 3090.135 ;
        RECT 210.370 3074.665 210.650 3074.945 ;
        RECT 214.430 3074.665 214.710 3074.945 ;
        RECT 3370.360 3028.055 3370.640 3028.335 ;
        RECT 3377.325 3028.055 3377.605 3028.335 ;
        RECT 3369.825 3012.875 3370.105 3013.155 ;
        RECT 3377.185 3012.875 3377.465 3013.155 ;
        RECT 3374.105 3006.435 3374.385 3006.715 ;
        RECT 3377.095 3006.435 3377.375 3006.715 ;
        RECT 3370.850 2975.615 3371.130 2975.895 ;
        RECT 3377.170 2975.615 3377.450 2975.895 ;
        RECT 3374.140 2966.415 3374.400 2966.675 ;
        RECT 3377.525 2966.415 3377.785 2966.675 ;
        RECT 210.370 2920.335 210.650 2920.615 ;
        RECT 212.085 2920.335 212.365 2920.615 ;
        RECT 210.525 2912.130 210.805 2912.410 ;
        RECT 213.920 2912.115 214.200 2912.395 ;
        RECT 210.370 2880.275 210.650 2880.555 ;
        RECT 212.070 2880.275 212.350 2880.555 ;
        RECT 210.370 2873.855 210.650 2874.135 ;
        RECT 214.955 2873.855 215.235 2874.135 ;
        RECT 210.370 2858.665 210.650 2858.945 ;
        RECT 214.430 2858.665 214.710 2858.945 ;
        RECT 3370.360 2802.055 3370.640 2802.335 ;
        RECT 3377.325 2802.055 3377.605 2802.335 ;
        RECT 3369.825 2786.875 3370.105 2787.155 ;
        RECT 3377.185 2786.875 3377.465 2787.155 ;
        RECT 3374.255 2780.435 3374.535 2780.715 ;
        RECT 3377.095 2780.435 3377.375 2780.715 ;
        RECT 3370.850 2749.615 3371.130 2749.895 ;
        RECT 3377.170 2749.615 3377.450 2749.895 ;
        RECT 3374.290 2740.415 3374.550 2740.675 ;
        RECT 3377.525 2740.415 3377.785 2740.675 ;
        RECT 210.370 2704.335 210.650 2704.615 ;
        RECT 211.985 2704.335 212.265 2704.615 ;
        RECT 210.370 2695.115 210.650 2695.395 ;
        RECT 213.920 2695.115 214.200 2695.395 ;
        RECT 210.370 2664.275 210.650 2664.555 ;
        RECT 211.970 2664.275 212.250 2664.555 ;
        RECT 210.370 2657.855 210.650 2658.135 ;
        RECT 214.955 2657.855 215.235 2658.135 ;
        RECT 210.370 2642.665 210.650 2642.945 ;
        RECT 214.430 2642.665 214.710 2642.945 ;
        RECT 210.370 2066.335 210.650 2066.615 ;
        RECT 212.385 2066.335 212.665 2066.615 ;
        RECT 210.370 2057.115 210.650 2057.395 ;
        RECT 213.920 2057.115 214.200 2057.395 ;
        RECT 210.370 2026.275 210.650 2026.555 ;
        RECT 212.370 2026.275 212.650 2026.555 ;
        RECT 210.370 2019.855 210.650 2020.135 ;
        RECT 214.955 2019.855 215.235 2020.135 ;
        RECT 210.370 2004.665 210.650 2004.945 ;
        RECT 214.430 2004.665 214.710 2004.945 ;
        RECT 3370.360 1916.055 3370.640 1916.335 ;
        RECT 3377.325 1916.055 3377.605 1916.335 ;
        RECT 3369.825 1900.875 3370.105 1901.155 ;
        RECT 3377.185 1900.875 3377.465 1901.155 ;
        RECT 3374.255 1894.435 3374.535 1894.715 ;
        RECT 3377.095 1894.435 3377.375 1894.715 ;
        RECT 3370.850 1863.615 3371.130 1863.895 ;
        RECT 3377.170 1863.615 3377.450 1863.895 ;
        RECT 3374.290 1854.415 3374.550 1854.675 ;
        RECT 3377.525 1854.415 3377.785 1854.675 ;
        RECT 210.370 1850.335 210.650 1850.615 ;
        RECT 212.385 1850.335 212.665 1850.615 ;
        RECT 210.370 1841.115 210.650 1841.395 ;
        RECT 213.920 1841.115 214.200 1841.395 ;
        RECT 210.370 1810.275 210.650 1810.555 ;
        RECT 212.370 1810.275 212.650 1810.555 ;
        RECT 210.370 1803.855 210.650 1804.135 ;
        RECT 214.955 1803.855 215.235 1804.135 ;
        RECT 210.370 1788.665 210.650 1788.945 ;
        RECT 214.430 1788.665 214.710 1788.945 ;
        RECT 3370.360 1690.055 3370.640 1690.335 ;
        RECT 3377.325 1690.055 3377.605 1690.335 ;
        RECT 3369.825 1674.875 3370.105 1675.155 ;
        RECT 3377.185 1674.875 3377.465 1675.155 ;
        RECT 3373.255 1668.435 3373.535 1668.715 ;
        RECT 3377.095 1668.435 3377.375 1668.715 ;
        RECT 3370.850 1637.615 3371.130 1637.895 ;
        RECT 3377.170 1637.615 3377.450 1637.895 ;
        RECT 210.370 1634.335 210.650 1634.615 ;
        RECT 212.385 1634.335 212.665 1634.615 ;
        RECT 3373.290 1628.415 3373.550 1628.675 ;
        RECT 3377.525 1628.415 3377.785 1628.675 ;
        RECT 210.370 1625.115 210.650 1625.395 ;
        RECT 213.920 1625.115 214.200 1625.395 ;
        RECT 210.370 1594.275 210.650 1594.555 ;
        RECT 212.370 1594.275 212.650 1594.555 ;
        RECT 210.370 1587.855 210.650 1588.135 ;
        RECT 214.955 1587.855 215.235 1588.135 ;
        RECT 210.370 1572.665 210.650 1572.945 ;
        RECT 214.430 1572.665 214.710 1572.945 ;
        RECT 3370.360 1465.055 3370.640 1465.335 ;
        RECT 3377.325 1465.055 3377.605 1465.335 ;
        RECT 3369.825 1449.875 3370.105 1450.155 ;
        RECT 3377.185 1449.875 3377.465 1450.155 ;
        RECT 3373.255 1443.435 3373.535 1443.715 ;
        RECT 3377.095 1443.435 3377.375 1443.715 ;
        RECT 210.370 1418.335 210.650 1418.615 ;
        RECT 212.385 1418.335 212.665 1418.615 ;
        RECT 3370.850 1412.615 3371.130 1412.895 ;
        RECT 3377.170 1412.615 3377.450 1412.895 ;
        RECT 210.370 1409.115 210.650 1409.395 ;
        RECT 213.920 1409.115 214.200 1409.395 ;
        RECT 3373.290 1403.415 3373.550 1403.675 ;
        RECT 3377.525 1403.415 3377.785 1403.675 ;
        RECT 210.370 1378.275 210.650 1378.555 ;
        RECT 212.370 1378.275 212.650 1378.555 ;
        RECT 210.370 1371.855 210.650 1372.135 ;
        RECT 214.955 1371.855 215.235 1372.135 ;
        RECT 210.370 1356.665 210.650 1356.945 ;
        RECT 214.430 1356.665 214.710 1356.945 ;
        RECT 3370.360 1240.055 3370.640 1240.335 ;
        RECT 3377.325 1240.055 3377.605 1240.335 ;
        RECT 3369.825 1224.875 3370.105 1225.155 ;
        RECT 3377.185 1224.875 3377.465 1225.155 ;
        RECT 3373.255 1218.435 3373.535 1218.715 ;
        RECT 3377.095 1218.435 3377.375 1218.715 ;
        RECT 210.370 1202.335 210.650 1202.615 ;
        RECT 212.385 1202.335 212.665 1202.615 ;
        RECT 210.370 1193.115 210.650 1193.395 ;
        RECT 213.920 1193.115 214.200 1193.395 ;
        RECT 3370.850 1187.615 3371.130 1187.895 ;
        RECT 3377.170 1187.615 3377.450 1187.895 ;
        RECT 3373.290 1178.415 3373.550 1178.675 ;
        RECT 3377.525 1178.415 3377.785 1178.675 ;
        RECT 210.370 1162.275 210.650 1162.555 ;
        RECT 212.370 1162.275 212.650 1162.555 ;
        RECT 210.370 1155.855 210.650 1156.135 ;
        RECT 214.955 1155.855 215.235 1156.135 ;
        RECT 210.370 1140.665 210.650 1140.945 ;
        RECT 214.430 1140.665 214.710 1140.945 ;
        RECT 3370.360 1014.055 3370.640 1014.335 ;
        RECT 3377.325 1014.055 3377.605 1014.335 ;
        RECT 3369.825 998.875 3370.105 999.155 ;
        RECT 3377.185 998.875 3377.465 999.155 ;
        RECT 3373.255 992.435 3373.535 992.715 ;
        RECT 3377.095 992.435 3377.375 992.715 ;
        RECT 210.370 986.335 210.650 986.615 ;
        RECT 212.385 986.335 212.665 986.615 ;
        RECT 210.370 977.115 210.650 977.395 ;
        RECT 213.920 977.115 214.200 977.395 ;
        RECT 3370.850 961.615 3371.130 961.895 ;
        RECT 3377.170 961.615 3377.450 961.895 ;
        RECT 3373.290 952.415 3373.550 952.675 ;
        RECT 3377.525 952.415 3377.785 952.675 ;
        RECT 210.370 946.275 210.650 946.555 ;
        RECT 212.370 946.275 212.650 946.555 ;
        RECT 210.370 939.855 210.650 940.135 ;
        RECT 214.955 939.855 215.235 940.135 ;
        RECT 210.370 924.665 210.650 924.945 ;
        RECT 214.430 924.665 214.710 924.945 ;
        RECT 213.950 905.140 214.210 905.400 ;
        RECT 214.460 904.640 214.720 904.900 ;
        RECT 214.950 904.140 215.210 904.400 ;
        RECT 211.080 347.205 211.445 349.835 ;
        RECT 3370.360 789.055 3370.640 789.335 ;
        RECT 3377.325 789.055 3377.605 789.335 ;
        RECT 3369.825 773.875 3370.105 774.155 ;
        RECT 3377.185 773.875 3377.465 774.155 ;
        RECT 3373.255 767.435 3373.535 767.715 ;
        RECT 3377.095 767.435 3377.375 767.715 ;
        RECT 3370.850 736.615 3371.130 736.895 ;
        RECT 3377.170 736.615 3377.450 736.895 ;
        RECT 3373.290 727.415 3373.550 727.675 ;
        RECT 3377.525 727.415 3377.785 727.675 ;
        RECT 212.140 561.855 212.550 563.670 ;
        RECT 3370.360 563.055 3370.640 563.335 ;
        RECT 3377.325 563.055 3377.605 563.335 ;
        RECT 211.605 212.060 211.870 212.720 ;
        RECT 3369.825 547.875 3370.105 548.155 ;
        RECT 3377.185 547.875 3377.465 548.155 ;
        RECT 3373.255 541.435 3373.535 541.715 ;
        RECT 3377.095 541.435 3377.375 541.715 ;
        RECT 3370.850 510.615 3371.130 510.895 ;
        RECT 3377.170 510.615 3377.450 510.895 ;
        RECT 3373.290 501.415 3373.550 501.675 ;
        RECT 3377.525 501.415 3377.785 501.675 ;
        RECT 2856.730 213.005 2858.685 214.805 ;
        RECT 3370.355 212.925 3370.615 213.185 ;
        RECT 1476.430 212.515 1476.690 212.775 ;
        RECT 1516.450 212.515 1516.710 212.775 ;
        RECT 1750.430 212.515 1750.690 212.775 ;
        RECT 1790.450 212.515 1790.710 212.775 ;
        RECT 2024.430 212.515 2024.690 212.775 ;
        RECT 2064.450 212.515 2064.710 212.775 ;
        RECT 212.910 212.060 213.670 212.320 ;
        RECT 704.980 212.060 705.240 212.320 ;
        RECT 712.850 212.060 713.110 212.320 ;
        RECT 715.375 212.060 715.635 212.320 ;
        RECT 717.160 212.060 717.420 212.320 ;
        RECT 723.010 212.060 723.270 212.320 ;
        RECT 979.910 211.415 980.170 211.675 ;
        RECT 1522.910 211.415 1523.170 211.675 ;
        RECT 1796.910 211.415 1797.170 211.675 ;
        RECT 2070.910 211.415 2071.170 211.675 ;
        RECT 2344.910 211.415 2345.170 211.675 ;
        RECT 2618.910 212.285 2619.170 212.545 ;
        RECT 3369.830 212.285 3370.090 212.545 ;
        RECT 454.360 210.915 455.425 211.195 ;
        RECT 995.110 210.915 995.370 211.175 ;
        RECT 1538.080 210.915 1538.340 211.175 ;
        RECT 1812.080 210.915 1812.340 211.175 ;
        RECT 2086.080 210.915 2086.340 211.175 ;
        RECT 2360.080 210.915 2360.340 211.175 ;
        RECT 2634.080 211.785 2634.340 212.045 ;
        RECT 729.265 210.410 729.535 210.680 ;
        RECT 942.630 210.415 942.890 210.675 ;
        RECT 964.230 210.415 964.490 210.675 ;
        RECT 1007.460 210.415 1007.720 210.675 ;
        RECT 1485.630 210.415 1485.890 210.675 ;
        RECT 1498.035 210.380 1498.315 210.660 ;
        RECT 1528.855 210.370 1529.135 210.650 ;
        RECT 1759.630 210.415 1759.890 210.675 ;
        RECT 1772.035 210.390 1772.315 210.670 ;
        RECT 1802.855 210.415 1803.135 210.695 ;
        RECT 2033.630 210.415 2033.890 210.675 ;
        RECT 2307.630 210.415 2307.890 210.675 ;
        RECT 2581.630 211.285 2581.890 211.545 ;
        RECT 3370.830 211.285 3371.090 211.545 ;
        RECT 945.840 209.915 946.100 210.175 ;
        RECT 955.050 209.915 955.310 210.175 ;
        RECT 961.000 209.915 961.260 210.175 ;
        RECT 967.500 209.915 967.760 210.175 ;
        RECT 982.620 209.915 982.880 210.175 ;
        RECT 985.880 209.915 986.140 210.175 ;
        RECT 989.080 209.915 989.340 210.175 ;
        RECT 991.870 209.915 992.130 210.175 ;
        RECT 1001.070 209.915 1001.330 210.175 ;
        RECT 1004.260 209.915 1004.520 210.175 ;
        RECT 1268.110 209.810 1269.075 210.170 ;
        RECT 1488.840 209.915 1489.100 210.175 ;
        RECT 1504.000 209.915 1504.260 210.175 ;
        RECT 1507.235 209.885 1507.515 210.165 ;
        RECT 1510.500 209.915 1510.760 210.175 ;
        RECT 1525.620 209.915 1525.880 210.175 ;
        RECT 1532.080 209.915 1532.340 210.175 ;
        RECT 1544.070 209.915 1544.330 210.175 ;
        RECT 1547.260 209.915 1547.520 210.175 ;
        RECT 1762.840 209.915 1763.100 210.175 ;
        RECT 1778.000 209.915 1778.260 210.175 ;
        RECT 1781.235 209.870 1781.515 210.150 ;
        RECT 1784.500 209.915 1784.760 210.175 ;
        RECT 1799.620 209.915 1799.880 210.175 ;
        RECT 1806.080 209.915 1806.340 210.175 ;
        RECT 1818.070 209.915 1818.330 210.175 ;
        RECT 1821.260 209.915 1821.520 210.175 ;
        RECT 2036.840 209.915 2037.100 210.175 ;
        RECT 2052.000 209.915 2052.260 210.175 ;
        RECT 2058.500 209.915 2058.760 210.175 ;
        RECT 2073.620 209.915 2073.880 210.175 ;
        RECT 2080.080 209.915 2080.340 210.175 ;
        RECT 2092.070 209.915 2092.330 210.175 ;
        RECT 2095.260 209.915 2095.520 210.175 ;
        RECT 2310.840 209.915 2311.100 210.175 ;
        RECT 2326.000 209.915 2326.260 210.175 ;
        RECT 2332.500 209.915 2332.760 210.175 ;
        RECT 2347.620 209.915 2347.880 210.175 ;
        RECT 2354.080 209.915 2354.340 210.175 ;
        RECT 2366.070 209.915 2366.330 210.175 ;
        RECT 2369.260 209.915 2369.520 210.175 ;
        RECT 2584.840 210.785 2585.100 211.045 ;
        RECT 2600.000 210.785 2600.260 211.045 ;
        RECT 2606.500 210.785 2606.760 211.045 ;
        RECT 2621.620 210.785 2621.880 211.045 ;
        RECT 2628.080 210.785 2628.340 211.045 ;
        RECT 2640.070 210.785 2640.330 211.045 ;
        RECT 2643.260 210.785 2643.520 211.045 ;
        RECT 2572.430 210.335 2572.690 210.595 ;
        RECT 2612.450 210.335 2612.710 210.595 ;
        RECT 933.430 209.465 933.690 209.725 ;
        RECT 973.450 209.465 973.710 209.725 ;
        RECT 2298.430 209.465 2298.690 209.725 ;
        RECT 2338.450 209.465 2338.710 209.725 ;
        RECT 664.990 200.880 665.250 201.140 ;
        RECT 719.625 200.880 719.885 201.140 ;
        RECT 712.850 200.350 713.110 200.610 ;
      LAYER met2 ;
        RECT 390.250 5034.255 456.440 5036.855 ;
        RECT 647.250 5034.255 713.440 5036.855 ;
        RECT 904.250 5034.255 970.440 5036.855 ;
        RECT 1152.265 5013.940 1226.290 5183.075 ;
        RECT 1415.265 5013.940 1489.290 5183.075 ;
        RECT 1152.265 4990.335 1202.110 5013.940 ;
        RECT 1415.265 4990.335 1465.110 5013.940 ;
        RECT 1176.675 4990.035 1202.110 4990.335 ;
        RECT 1439.675 4990.035 1465.110 4990.335 ;
        RECT 1667.265 4990.035 1741.290 5183.075 ;
        RECT 1924.265 5013.940 1998.290 5183.075 ;
        RECT 2373.250 5034.255 2439.440 5036.855 ;
        RECT 2630.250 5034.255 2696.440 5036.855 ;
        RECT 1924.265 4990.335 1974.110 5013.940 ;
        RECT 1948.675 4990.035 1974.110 4990.335 ;
        RECT 2878.265 4990.035 2952.290 5183.075 ;
        RECT 3139.250 5034.255 3205.440 5036.855 ;
        RECT 1177.895 4988.000 1179.895 4989.920 ;
        RECT 1440.895 4988.000 1442.895 4989.920 ;
        RECT 1667.495 4988.000 1691.395 4990.035 ;
        RECT 1692.895 4988.000 1694.895 4989.920 ;
        RECT 1717.390 4988.000 1741.290 4990.035 ;
        RECT 1949.895 4988.000 1951.895 4989.920 ;
        RECT 2878.495 4988.000 2902.395 4990.035 ;
        RECT 2903.895 4988.000 2905.895 4989.920 ;
        RECT 2928.390 4988.000 2952.290 4990.035 ;
        RECT 151.145 4780.250 153.745 4846.440 ;
        RECT 3434.255 4762.560 3436.855 4828.750 ;
        RECT 4.925 4399.390 200.000 4423.290 ;
        RECT 4.925 4373.395 197.965 4399.390 ;
        RECT 3379.435 4390.795 3588.000 4391.790 ;
        RECT 3379.715 4389.955 3588.000 4390.795 ;
        RECT 3379.435 4388.035 3588.000 4389.955 ;
        RECT 3379.715 4387.195 3588.000 4388.035 ;
        RECT 3379.435 4384.815 3588.000 4387.195 ;
        RECT 3379.715 4383.975 3588.000 4384.815 ;
        RECT 3379.435 4381.595 3588.000 4383.975 ;
        RECT 3379.715 4380.755 3588.000 4381.595 ;
        RECT 3379.435 4378.835 3588.000 4380.755 ;
        RECT 3379.715 4377.995 3588.000 4378.835 ;
        RECT 198.080 4374.895 200.000 4376.895 ;
        RECT 3379.435 4375.615 3588.000 4377.995 ;
      LAYER met2 ;
        RECT 3370.330 4375.365 3370.580 4375.510 ;
        RECT 3370.330 4375.025 3370.640 4375.365 ;
        RECT 3377.035 4375.055 3379.435 4375.335 ;
      LAYER met2 ;
        RECT 4.925 4349.495 200.000 4373.395 ;
      LAYER met2 ;
        RECT 3369.830 4360.185 3370.080 4360.275 ;
        RECT 3369.805 4359.845 3370.105 4360.185 ;
      LAYER met2 ;
        RECT 4.925 4349.265 197.965 4349.495 ;
        RECT 4.925 4188.390 200.000 4212.290 ;
        RECT 4.925 4162.395 197.965 4188.390 ;
        RECT 198.080 4163.895 200.000 4165.895 ;
        RECT 4.925 4138.495 200.000 4162.395 ;
        RECT 4.925 4138.265 197.965 4138.495 ;
        RECT 0.000 4000.865 208.565 4001.915 ;
        RECT 0.000 4000.025 208.285 4000.865 ;
      LAYER met2 ;
        RECT 212.370 4000.645 212.650 4000.720 ;
        RECT 210.370 4000.625 210.650 4000.645 ;
        RECT 209.945 4000.605 210.965 4000.625 ;
        RECT 209.910 4000.585 210.965 4000.605 ;
        RECT 208.565 4000.305 210.965 4000.585 ;
        RECT 212.370 4000.305 212.665 4000.645 ;
      LAYER met2 ;
        RECT 0.000 3997.645 208.565 4000.025 ;
        RECT 0.000 3996.805 208.285 3997.645 ;
        RECT 0.000 3994.425 208.565 3996.805 ;
        RECT 0.000 3993.585 208.285 3994.425 ;
      LAYER met2 ;
        RECT 208.565 3993.865 210.965 3994.145 ;
      LAYER met2 ;
        RECT 0.000 3991.665 208.565 3993.585 ;
        RECT 0.000 3990.825 208.285 3991.665 ;
      LAYER met2 ;
        RECT 210.370 3991.405 210.650 3991.425 ;
        RECT 209.945 3991.385 210.965 3991.405 ;
        RECT 208.565 3991.105 210.965 3991.385 ;
        RECT 210.370 3991.085 210.650 3991.105 ;
      LAYER met2 ;
        RECT 0.000 3988.445 208.565 3990.825 ;
        RECT 0.000 3987.605 208.285 3988.445 ;
        RECT 0.000 3985.225 208.565 3987.605 ;
        RECT 0.000 3984.385 208.285 3985.225 ;
        RECT 0.000 3982.465 208.565 3984.385 ;
        RECT 0.000 3981.625 208.285 3982.465 ;
      LAYER met2 ;
        RECT 208.565 3981.905 210.965 3982.185 ;
      LAYER met2 ;
        RECT 0.000 3979.245 208.565 3981.625 ;
        RECT 0.000 3978.405 208.285 3979.245 ;
        RECT 0.000 3976.025 208.565 3978.405 ;
        RECT 0.000 3975.185 208.285 3976.025 ;
        RECT 0.000 3973.265 208.565 3975.185 ;
        RECT 0.000 3972.425 208.285 3973.265 ;
        RECT 0.000 3970.045 208.565 3972.425 ;
        RECT 0.000 3969.205 208.285 3970.045 ;
        RECT 0.000 3966.825 208.565 3969.205 ;
        RECT 0.000 3965.985 208.285 3966.825 ;
        RECT 0.000 3964.065 208.565 3965.985 ;
        RECT 0.000 3963.225 208.285 3964.065 ;
        RECT 0.000 3960.845 208.565 3963.225 ;
        RECT 0.000 3960.005 208.285 3960.845 ;
      LAYER met2 ;
        RECT 210.370 3960.565 210.650 3960.585 ;
        RECT 208.565 3960.285 210.965 3960.565 ;
        RECT 209.400 3960.265 210.965 3960.285 ;
        RECT 210.370 3960.245 210.650 3960.265 ;
        RECT 212.370 3960.245 212.650 4000.305 ;
        RECT 213.960 3991.425 214.210 3991.775 ;
        RECT 213.920 3991.085 214.210 3991.425 ;
      LAYER met2 ;
        RECT 0.000 3957.625 208.565 3960.005 ;
        RECT 0.000 3956.785 208.285 3957.625 ;
        RECT 0.000 3954.405 208.565 3956.785 ;
        RECT 0.000 3953.565 208.285 3954.405 ;
      LAYER met2 ;
        RECT 210.370 3954.135 210.650 3954.165 ;
        RECT 210.145 3954.125 210.965 3954.135 ;
        RECT 208.565 3953.845 210.965 3954.125 ;
        RECT 210.370 3953.825 210.650 3953.845 ;
      LAYER met2 ;
        RECT 0.000 3951.645 208.565 3953.565 ;
        RECT 0.000 3950.805 208.285 3951.645 ;
        RECT 0.000 3948.425 208.565 3950.805 ;
        RECT 0.000 3947.585 208.285 3948.425 ;
        RECT 0.000 3945.205 208.565 3947.585 ;
        RECT 0.000 3944.365 208.285 3945.205 ;
        RECT 0.000 3942.445 208.565 3944.365 ;
        RECT 0.000 3941.605 208.285 3942.445 ;
        RECT 0.000 3939.225 208.565 3941.605 ;
        RECT 0.000 3938.385 208.285 3939.225 ;
      LAYER met2 ;
        RECT 210.370 3938.945 210.650 3938.975 ;
        RECT 208.565 3938.665 210.965 3938.945 ;
        RECT 210.370 3938.635 210.650 3938.665 ;
      LAYER met2 ;
        RECT 0.000 3936.005 208.565 3938.385 ;
        RECT 0.000 3935.165 208.285 3936.005 ;
        RECT 0.000 3933.245 208.565 3935.165 ;
        RECT 0.000 3932.405 208.285 3933.245 ;
        RECT 0.000 3930.025 208.565 3932.405 ;
        RECT 0.000 3929.185 208.285 3930.025 ;
        RECT 0.000 3926.805 208.565 3929.185 ;
        RECT 0.000 3925.965 208.285 3926.805 ;
        RECT 0.000 3924.045 208.565 3925.965 ;
        RECT 0.000 3923.205 208.285 3924.045 ;
        RECT 0.000 3922.210 208.565 3923.205 ;
        RECT 0.000 3784.865 208.565 3785.915 ;
        RECT 0.000 3784.025 208.285 3784.865 ;
      LAYER met2 ;
        RECT 208.565 3784.305 210.965 3784.585 ;
      LAYER met2 ;
        RECT 0.000 3781.645 208.565 3784.025 ;
      LAYER met2 ;
        RECT 209.755 3782.305 210.035 3784.305 ;
        RECT 212.370 3782.645 212.650 3782.720 ;
        RECT 212.370 3782.305 212.665 3782.645 ;
      LAYER met2 ;
        RECT 0.000 3780.805 208.285 3781.645 ;
        RECT 0.000 3778.425 208.565 3780.805 ;
        RECT 0.000 3777.585 208.285 3778.425 ;
      LAYER met2 ;
        RECT 208.565 3777.865 210.965 3778.145 ;
      LAYER met2 ;
        RECT 0.000 3775.665 208.565 3777.585 ;
        RECT 0.000 3774.825 208.285 3775.665 ;
      LAYER met2 ;
        RECT 210.370 3775.405 210.650 3775.425 ;
        RECT 209.945 3775.385 210.965 3775.405 ;
        RECT 208.565 3775.105 210.965 3775.385 ;
        RECT 210.370 3775.085 210.650 3775.105 ;
      LAYER met2 ;
        RECT 0.000 3772.445 208.565 3774.825 ;
        RECT 0.000 3771.605 208.285 3772.445 ;
        RECT 0.000 3769.225 208.565 3771.605 ;
        RECT 0.000 3768.385 208.285 3769.225 ;
        RECT 0.000 3766.465 208.565 3768.385 ;
        RECT 0.000 3765.625 208.285 3766.465 ;
      LAYER met2 ;
        RECT 208.565 3765.905 210.965 3766.185 ;
      LAYER met2 ;
        RECT 0.000 3763.245 208.565 3765.625 ;
        RECT 0.000 3762.405 208.285 3763.245 ;
        RECT 0.000 3760.025 208.565 3762.405 ;
        RECT 0.000 3759.185 208.285 3760.025 ;
        RECT 0.000 3757.265 208.565 3759.185 ;
        RECT 0.000 3756.425 208.285 3757.265 ;
        RECT 0.000 3754.045 208.565 3756.425 ;
        RECT 0.000 3753.205 208.285 3754.045 ;
        RECT 0.000 3750.825 208.565 3753.205 ;
        RECT 0.000 3749.985 208.285 3750.825 ;
        RECT 0.000 3748.065 208.565 3749.985 ;
        RECT 0.000 3747.225 208.285 3748.065 ;
        RECT 0.000 3744.845 208.565 3747.225 ;
        RECT 0.000 3744.005 208.285 3744.845 ;
      LAYER met2 ;
        RECT 210.370 3744.565 210.650 3744.585 ;
        RECT 208.565 3744.285 210.965 3744.565 ;
        RECT 209.400 3744.265 210.965 3744.285 ;
        RECT 210.370 3744.245 210.650 3744.265 ;
        RECT 212.370 3744.245 212.650 3782.305 ;
        RECT 213.960 3775.425 214.210 3991.085 ;
        RECT 214.960 3954.165 215.210 3954.425 ;
        RECT 214.955 3953.825 215.235 3954.165 ;
        RECT 214.460 3938.975 214.710 3939.100 ;
        RECT 214.430 3938.635 214.710 3938.975 ;
        RECT 213.920 3775.085 214.210 3775.425 ;
      LAYER met2 ;
        RECT 0.000 3741.625 208.565 3744.005 ;
        RECT 0.000 3740.785 208.285 3741.625 ;
        RECT 0.000 3738.405 208.565 3740.785 ;
        RECT 0.000 3737.565 208.285 3738.405 ;
      LAYER met2 ;
        RECT 210.370 3738.135 210.650 3738.165 ;
        RECT 210.145 3738.125 210.965 3738.135 ;
        RECT 208.565 3737.845 210.965 3738.125 ;
        RECT 210.370 3737.825 210.650 3737.845 ;
      LAYER met2 ;
        RECT 0.000 3735.645 208.565 3737.565 ;
        RECT 0.000 3734.805 208.285 3735.645 ;
        RECT 0.000 3732.425 208.565 3734.805 ;
        RECT 0.000 3731.585 208.285 3732.425 ;
        RECT 0.000 3729.205 208.565 3731.585 ;
        RECT 0.000 3728.365 208.285 3729.205 ;
        RECT 0.000 3726.445 208.565 3728.365 ;
        RECT 0.000 3725.605 208.285 3726.445 ;
        RECT 0.000 3723.225 208.565 3725.605 ;
        RECT 0.000 3722.385 208.285 3723.225 ;
      LAYER met2 ;
        RECT 210.370 3722.945 210.650 3722.975 ;
        RECT 208.565 3722.665 210.965 3722.945 ;
        RECT 210.370 3722.635 210.650 3722.665 ;
      LAYER met2 ;
        RECT 0.000 3720.005 208.565 3722.385 ;
        RECT 0.000 3719.165 208.285 3720.005 ;
        RECT 0.000 3717.245 208.565 3719.165 ;
        RECT 0.000 3716.405 208.285 3717.245 ;
        RECT 0.000 3714.025 208.565 3716.405 ;
        RECT 0.000 3713.185 208.285 3714.025 ;
        RECT 0.000 3710.805 208.565 3713.185 ;
        RECT 0.000 3709.965 208.285 3710.805 ;
        RECT 0.000 3708.045 208.565 3709.965 ;
        RECT 0.000 3707.205 208.285 3708.045 ;
        RECT 0.000 3706.210 208.565 3707.205 ;
        RECT 0.000 3568.865 208.565 3569.915 ;
        RECT 0.000 3568.025 208.285 3568.865 ;
      LAYER met2 ;
        RECT 210.685 3568.585 210.965 3570.535 ;
        RECT 208.565 3568.305 210.965 3568.585 ;
      LAYER met2 ;
        RECT 0.000 3565.645 208.565 3568.025 ;
        RECT 0.000 3564.805 208.285 3565.645 ;
        RECT 0.000 3562.425 208.565 3564.805 ;
        RECT 0.000 3561.585 208.285 3562.425 ;
      LAYER met2 ;
        RECT 208.565 3561.865 210.965 3562.145 ;
      LAYER met2 ;
        RECT 0.000 3559.665 208.565 3561.585 ;
        RECT 0.000 3558.825 208.285 3559.665 ;
      LAYER met2 ;
        RECT 213.960 3559.425 214.210 3775.085 ;
        RECT 214.460 3722.975 214.710 3938.635 ;
        RECT 214.960 3738.165 215.210 3953.825 ;
        RECT 3369.830 3914.185 3370.080 4359.845 ;
        RECT 3370.330 3929.365 3370.580 4375.025 ;
      LAYER met2 ;
        RECT 3379.715 4374.775 3588.000 4375.615 ;
        RECT 3379.435 4372.395 3588.000 4374.775 ;
        RECT 3379.715 4371.555 3588.000 4372.395 ;
        RECT 3379.435 4369.635 3588.000 4371.555 ;
        RECT 3379.715 4368.795 3588.000 4369.635 ;
        RECT 3379.435 4366.415 3588.000 4368.795 ;
        RECT 3379.715 4365.575 3588.000 4366.415 ;
        RECT 3379.435 4363.195 3588.000 4365.575 ;
        RECT 3379.715 4362.355 3588.000 4363.195 ;
        RECT 3379.435 4360.435 3588.000 4362.355 ;
      LAYER met2 ;
        RECT 3377.035 4359.875 3379.435 4360.155 ;
      LAYER met2 ;
        RECT 3379.715 4359.595 3588.000 4360.435 ;
        RECT 3379.435 4357.215 3588.000 4359.595 ;
        RECT 3379.715 4356.375 3588.000 4357.215 ;
        RECT 3379.435 4353.995 3588.000 4356.375 ;
      LAYER met2 ;
        RECT 3374.290 4353.745 3374.570 4353.840 ;
        RECT 3374.255 4353.405 3374.570 4353.745 ;
        RECT 3377.035 4353.435 3379.435 4353.715 ;
        RECT 3370.830 4322.925 3371.080 4323.010 ;
        RECT 3370.830 4322.585 3371.130 4322.925 ;
        RECT 3370.330 3929.025 3370.640 3929.365 ;
        RECT 3369.805 3913.845 3370.105 3914.185 ;
        RECT 214.955 3737.825 215.235 3738.165 ;
        RECT 214.430 3722.635 214.710 3722.975 ;
        RECT 210.370 3559.405 210.650 3559.425 ;
        RECT 209.945 3559.385 210.965 3559.405 ;
        RECT 208.565 3559.105 210.965 3559.385 ;
        RECT 210.370 3559.085 210.650 3559.105 ;
        RECT 213.920 3559.085 214.210 3559.425 ;
      LAYER met2 ;
        RECT 0.000 3556.445 208.565 3558.825 ;
        RECT 0.000 3555.605 208.285 3556.445 ;
        RECT 0.000 3553.225 208.565 3555.605 ;
        RECT 0.000 3552.385 208.285 3553.225 ;
        RECT 0.000 3550.465 208.565 3552.385 ;
        RECT 0.000 3549.625 208.285 3550.465 ;
      LAYER met2 ;
        RECT 208.565 3549.905 210.965 3550.185 ;
      LAYER met2 ;
        RECT 0.000 3547.245 208.565 3549.625 ;
        RECT 0.000 3546.405 208.285 3547.245 ;
        RECT 0.000 3544.025 208.565 3546.405 ;
        RECT 0.000 3543.185 208.285 3544.025 ;
        RECT 0.000 3541.265 208.565 3543.185 ;
        RECT 0.000 3540.425 208.285 3541.265 ;
        RECT 0.000 3538.045 208.565 3540.425 ;
        RECT 0.000 3537.205 208.285 3538.045 ;
        RECT 0.000 3534.825 208.565 3537.205 ;
        RECT 0.000 3533.985 208.285 3534.825 ;
        RECT 0.000 3532.065 208.565 3533.985 ;
        RECT 0.000 3531.225 208.285 3532.065 ;
        RECT 0.000 3528.845 208.565 3531.225 ;
        RECT 0.000 3528.005 208.285 3528.845 ;
      LAYER met2 ;
        RECT 210.370 3528.565 210.650 3528.585 ;
        RECT 208.565 3528.285 210.965 3528.565 ;
        RECT 209.400 3528.265 210.965 3528.285 ;
        RECT 210.370 3528.245 210.650 3528.265 ;
      LAYER met2 ;
        RECT 0.000 3525.625 208.565 3528.005 ;
        RECT 0.000 3524.785 208.285 3525.625 ;
        RECT 0.000 3522.405 208.565 3524.785 ;
        RECT 0.000 3521.565 208.285 3522.405 ;
      LAYER met2 ;
        RECT 210.370 3522.135 210.650 3522.165 ;
        RECT 210.145 3522.125 210.965 3522.135 ;
        RECT 208.565 3521.845 210.965 3522.125 ;
        RECT 210.370 3521.825 210.650 3521.845 ;
      LAYER met2 ;
        RECT 0.000 3519.645 208.565 3521.565 ;
        RECT 0.000 3518.805 208.285 3519.645 ;
        RECT 0.000 3516.425 208.565 3518.805 ;
        RECT 0.000 3515.585 208.285 3516.425 ;
        RECT 0.000 3513.205 208.565 3515.585 ;
        RECT 0.000 3512.365 208.285 3513.205 ;
        RECT 0.000 3510.445 208.565 3512.365 ;
        RECT 0.000 3509.605 208.285 3510.445 ;
        RECT 0.000 3507.225 208.565 3509.605 ;
        RECT 0.000 3506.385 208.285 3507.225 ;
      LAYER met2 ;
        RECT 210.370 3506.945 210.650 3506.975 ;
        RECT 208.565 3506.665 210.965 3506.945 ;
        RECT 210.370 3506.635 210.650 3506.665 ;
      LAYER met2 ;
        RECT 0.000 3504.005 208.565 3506.385 ;
        RECT 0.000 3503.165 208.285 3504.005 ;
        RECT 0.000 3501.245 208.565 3503.165 ;
        RECT 0.000 3500.405 208.285 3501.245 ;
        RECT 0.000 3498.025 208.565 3500.405 ;
        RECT 0.000 3497.185 208.285 3498.025 ;
        RECT 0.000 3494.805 208.565 3497.185 ;
        RECT 0.000 3493.965 208.285 3494.805 ;
        RECT 0.000 3492.045 208.565 3493.965 ;
        RECT 0.000 3491.205 208.285 3492.045 ;
        RECT 0.000 3490.210 208.565 3491.205 ;
        RECT 0.000 3352.865 208.565 3353.915 ;
        RECT 0.000 3352.025 208.285 3352.865 ;
      LAYER met2 ;
        RECT 208.565 3352.305 210.965 3352.585 ;
      LAYER met2 ;
        RECT 0.000 3349.645 208.565 3352.025 ;
      LAYER met2 ;
        RECT 209.845 3350.305 210.125 3352.305 ;
        RECT 212.370 3350.645 212.650 3350.720 ;
        RECT 212.370 3350.305 212.665 3350.645 ;
      LAYER met2 ;
        RECT 0.000 3348.805 208.285 3349.645 ;
        RECT 0.000 3346.425 208.565 3348.805 ;
        RECT 0.000 3345.585 208.285 3346.425 ;
      LAYER met2 ;
        RECT 208.565 3345.865 210.965 3346.145 ;
      LAYER met2 ;
        RECT 0.000 3343.665 208.565 3345.585 ;
        RECT 0.000 3342.825 208.285 3343.665 ;
      LAYER met2 ;
        RECT 210.370 3343.405 210.650 3343.425 ;
        RECT 209.945 3343.385 210.965 3343.405 ;
        RECT 208.565 3343.105 210.965 3343.385 ;
        RECT 210.370 3343.085 210.650 3343.105 ;
      LAYER met2 ;
        RECT 0.000 3340.445 208.565 3342.825 ;
        RECT 0.000 3339.605 208.285 3340.445 ;
        RECT 0.000 3337.225 208.565 3339.605 ;
        RECT 0.000 3336.385 208.285 3337.225 ;
        RECT 0.000 3334.465 208.565 3336.385 ;
        RECT 0.000 3333.625 208.285 3334.465 ;
      LAYER met2 ;
        RECT 208.565 3333.905 210.965 3334.185 ;
      LAYER met2 ;
        RECT 0.000 3331.245 208.565 3333.625 ;
        RECT 0.000 3330.405 208.285 3331.245 ;
        RECT 0.000 3328.025 208.565 3330.405 ;
        RECT 0.000 3327.185 208.285 3328.025 ;
        RECT 0.000 3325.265 208.565 3327.185 ;
        RECT 0.000 3324.425 208.285 3325.265 ;
        RECT 0.000 3322.045 208.565 3324.425 ;
        RECT 0.000 3321.205 208.285 3322.045 ;
        RECT 0.000 3318.825 208.565 3321.205 ;
        RECT 0.000 3317.985 208.285 3318.825 ;
        RECT 0.000 3316.065 208.565 3317.985 ;
        RECT 0.000 3315.225 208.285 3316.065 ;
        RECT 0.000 3312.845 208.565 3315.225 ;
        RECT 0.000 3312.005 208.285 3312.845 ;
      LAYER met2 ;
        RECT 210.370 3312.565 210.650 3312.585 ;
        RECT 208.565 3312.285 210.965 3312.565 ;
        RECT 209.400 3312.265 210.965 3312.285 ;
        RECT 210.370 3312.245 210.650 3312.265 ;
        RECT 212.370 3312.245 212.650 3350.305 ;
        RECT 213.960 3343.425 214.210 3559.085 ;
        RECT 214.460 3506.975 214.710 3722.635 ;
        RECT 214.960 3522.165 215.210 3737.825 ;
        RECT 3369.830 3689.185 3370.080 3913.845 ;
        RECT 3370.330 3704.365 3370.580 3929.025 ;
        RECT 3370.830 3876.925 3371.080 4322.585 ;
        RECT 3374.290 4313.385 3374.570 4353.405 ;
      LAYER met2 ;
        RECT 3379.715 4353.155 3588.000 4353.995 ;
        RECT 3379.435 4350.775 3588.000 4353.155 ;
        RECT 3379.715 4349.935 3588.000 4350.775 ;
        RECT 3379.435 4348.015 3588.000 4349.935 ;
        RECT 3379.715 4347.175 3588.000 4348.015 ;
        RECT 3379.435 4344.795 3588.000 4347.175 ;
        RECT 3379.715 4343.955 3588.000 4344.795 ;
        RECT 3379.435 4341.575 3588.000 4343.955 ;
        RECT 3379.715 4340.735 3588.000 4341.575 ;
        RECT 3379.435 4338.815 3588.000 4340.735 ;
        RECT 3379.715 4337.975 3588.000 4338.815 ;
        RECT 3379.435 4335.595 3588.000 4337.975 ;
        RECT 3379.715 4334.755 3588.000 4335.595 ;
        RECT 3379.435 4332.375 3588.000 4334.755 ;
      LAYER met2 ;
        RECT 3377.035 4331.815 3379.435 4332.095 ;
      LAYER met2 ;
        RECT 3379.715 4331.535 3588.000 4332.375 ;
        RECT 3379.435 4329.615 3588.000 4331.535 ;
        RECT 3379.715 4328.775 3588.000 4329.615 ;
        RECT 3379.435 4326.395 3588.000 4328.775 ;
        RECT 3379.715 4325.555 3588.000 4326.395 ;
        RECT 3379.435 4323.175 3588.000 4325.555 ;
      LAYER met2 ;
        RECT 3377.035 4322.615 3379.435 4322.895 ;
      LAYER met2 ;
        RECT 3379.715 4322.335 3588.000 4323.175 ;
        RECT 3379.435 4320.415 3588.000 4322.335 ;
      LAYER met2 ;
        RECT 3377.035 4319.855 3379.435 4320.135 ;
      LAYER met2 ;
        RECT 3379.715 4319.575 3588.000 4320.415 ;
        RECT 3379.435 4317.195 3588.000 4319.575 ;
        RECT 3379.715 4316.355 3588.000 4317.195 ;
        RECT 3379.435 4313.975 3588.000 4316.355 ;
      LAYER met2 ;
        RECT 3377.525 4313.695 3377.785 4313.705 ;
        RECT 3377.035 4313.415 3379.435 4313.695 ;
        RECT 3377.525 4313.385 3377.785 4313.415 ;
      LAYER met2 ;
        RECT 3379.715 4313.135 3588.000 4313.975 ;
        RECT 3379.435 4312.085 3588.000 4313.135 ;
        RECT 3390.035 4166.505 3583.075 4166.735 ;
        RECT 3388.000 4142.605 3583.075 4166.505 ;
        RECT 3388.000 4139.105 3389.920 4141.105 ;
        RECT 3390.035 4116.610 3583.075 4142.605 ;
        RECT 3388.000 4092.710 3583.075 4116.610 ;
        RECT 3379.435 3944.795 3588.000 3945.790 ;
        RECT 3379.715 3943.955 3588.000 3944.795 ;
        RECT 3379.435 3942.035 3588.000 3943.955 ;
        RECT 3379.715 3941.195 3588.000 3942.035 ;
        RECT 3379.435 3938.815 3588.000 3941.195 ;
        RECT 3379.715 3937.975 3588.000 3938.815 ;
        RECT 3379.435 3935.595 3588.000 3937.975 ;
        RECT 3379.715 3934.755 3588.000 3935.595 ;
        RECT 3379.435 3932.835 3588.000 3934.755 ;
        RECT 3379.715 3931.995 3588.000 3932.835 ;
        RECT 3379.435 3929.615 3588.000 3931.995 ;
      LAYER met2 ;
        RECT 3377.035 3929.055 3379.435 3929.335 ;
      LAYER met2 ;
        RECT 3379.715 3928.775 3588.000 3929.615 ;
        RECT 3379.435 3926.395 3588.000 3928.775 ;
        RECT 3379.715 3925.555 3588.000 3926.395 ;
        RECT 3379.435 3923.635 3588.000 3925.555 ;
        RECT 3379.715 3922.795 3588.000 3923.635 ;
        RECT 3379.435 3920.415 3588.000 3922.795 ;
        RECT 3379.715 3919.575 3588.000 3920.415 ;
        RECT 3379.435 3917.195 3588.000 3919.575 ;
        RECT 3379.715 3916.355 3588.000 3917.195 ;
        RECT 3379.435 3914.435 3588.000 3916.355 ;
      LAYER met2 ;
        RECT 3377.035 3913.875 3379.435 3914.155 ;
      LAYER met2 ;
        RECT 3379.715 3913.595 3588.000 3914.435 ;
        RECT 3379.435 3911.215 3588.000 3913.595 ;
        RECT 3379.715 3910.375 3588.000 3911.215 ;
        RECT 3379.435 3907.995 3588.000 3910.375 ;
      LAYER met2 ;
        RECT 3374.290 3907.745 3374.570 3907.840 ;
        RECT 3374.255 3907.405 3374.570 3907.745 ;
        RECT 3377.035 3907.435 3379.435 3907.715 ;
        RECT 3370.830 3876.585 3371.130 3876.925 ;
        RECT 3370.330 3704.025 3370.640 3704.365 ;
        RECT 3369.805 3688.845 3370.105 3689.185 ;
        RECT 215.515 3528.585 215.795 3570.535 ;
        RECT 215.515 3528.245 215.820 3528.585 ;
        RECT 215.515 3528.240 215.795 3528.245 ;
        RECT 214.955 3521.825 215.235 3522.165 ;
        RECT 214.430 3506.635 214.710 3506.975 ;
        RECT 213.920 3343.085 214.210 3343.425 ;
      LAYER met2 ;
        RECT 0.000 3309.625 208.565 3312.005 ;
        RECT 0.000 3308.785 208.285 3309.625 ;
        RECT 0.000 3306.405 208.565 3308.785 ;
        RECT 0.000 3305.565 208.285 3306.405 ;
      LAYER met2 ;
        RECT 210.370 3306.135 210.650 3306.165 ;
        RECT 210.145 3306.125 210.965 3306.135 ;
        RECT 208.565 3305.845 210.965 3306.125 ;
        RECT 210.370 3305.825 210.650 3305.845 ;
      LAYER met2 ;
        RECT 0.000 3303.645 208.565 3305.565 ;
        RECT 0.000 3302.805 208.285 3303.645 ;
        RECT 0.000 3300.425 208.565 3302.805 ;
        RECT 0.000 3299.585 208.285 3300.425 ;
        RECT 0.000 3297.205 208.565 3299.585 ;
        RECT 0.000 3296.365 208.285 3297.205 ;
        RECT 0.000 3294.445 208.565 3296.365 ;
        RECT 0.000 3293.605 208.285 3294.445 ;
        RECT 0.000 3291.225 208.565 3293.605 ;
        RECT 0.000 3290.385 208.285 3291.225 ;
      LAYER met2 ;
        RECT 210.370 3290.945 210.650 3290.975 ;
        RECT 208.565 3290.665 210.965 3290.945 ;
        RECT 210.370 3290.635 210.650 3290.665 ;
      LAYER met2 ;
        RECT 0.000 3288.005 208.565 3290.385 ;
        RECT 0.000 3287.165 208.285 3288.005 ;
        RECT 0.000 3285.245 208.565 3287.165 ;
        RECT 0.000 3284.405 208.285 3285.245 ;
        RECT 0.000 3282.025 208.565 3284.405 ;
        RECT 0.000 3281.185 208.285 3282.025 ;
        RECT 0.000 3278.805 208.565 3281.185 ;
        RECT 0.000 3277.965 208.285 3278.805 ;
        RECT 0.000 3276.045 208.565 3277.965 ;
        RECT 0.000 3275.205 208.285 3276.045 ;
        RECT 0.000 3274.210 208.565 3275.205 ;
        RECT 0.000 3136.865 208.565 3137.915 ;
        RECT 0.000 3136.025 208.285 3136.865 ;
      LAYER met2 ;
        RECT 212.370 3136.645 212.650 3136.720 ;
        RECT 210.370 3136.625 210.650 3136.645 ;
        RECT 209.945 3136.605 210.965 3136.625 ;
        RECT 209.910 3136.585 210.965 3136.605 ;
        RECT 208.565 3136.305 210.965 3136.585 ;
        RECT 212.370 3136.305 212.665 3136.645 ;
      LAYER met2 ;
        RECT 0.000 3133.645 208.565 3136.025 ;
        RECT 0.000 3132.805 208.285 3133.645 ;
        RECT 0.000 3130.425 208.565 3132.805 ;
        RECT 0.000 3129.585 208.285 3130.425 ;
      LAYER met2 ;
        RECT 208.565 3129.865 210.965 3130.145 ;
      LAYER met2 ;
        RECT 0.000 3127.665 208.565 3129.585 ;
      LAYER met2 ;
        RECT 210.345 3128.425 210.625 3128.455 ;
        RECT 210.345 3128.405 210.650 3128.425 ;
        RECT 210.290 3128.105 210.715 3128.405 ;
        RECT 210.345 3128.085 210.650 3128.105 ;
      LAYER met2 ;
        RECT 0.000 3126.825 208.285 3127.665 ;
      LAYER met2 ;
        RECT 210.345 3127.385 210.625 3128.085 ;
        RECT 208.565 3127.105 210.965 3127.385 ;
      LAYER met2 ;
        RECT 0.000 3124.445 208.565 3126.825 ;
        RECT 0.000 3123.605 208.285 3124.445 ;
        RECT 0.000 3121.225 208.565 3123.605 ;
        RECT 0.000 3120.385 208.285 3121.225 ;
        RECT 0.000 3118.465 208.565 3120.385 ;
        RECT 0.000 3117.625 208.285 3118.465 ;
      LAYER met2 ;
        RECT 208.565 3117.905 210.965 3118.185 ;
      LAYER met2 ;
        RECT 0.000 3115.245 208.565 3117.625 ;
        RECT 0.000 3114.405 208.285 3115.245 ;
        RECT 0.000 3112.025 208.565 3114.405 ;
        RECT 0.000 3111.185 208.285 3112.025 ;
        RECT 0.000 3109.265 208.565 3111.185 ;
        RECT 0.000 3108.425 208.285 3109.265 ;
        RECT 0.000 3106.045 208.565 3108.425 ;
        RECT 0.000 3105.205 208.285 3106.045 ;
        RECT 0.000 3102.825 208.565 3105.205 ;
        RECT 0.000 3101.985 208.285 3102.825 ;
        RECT 0.000 3100.065 208.565 3101.985 ;
        RECT 0.000 3099.225 208.285 3100.065 ;
        RECT 0.000 3096.845 208.565 3099.225 ;
        RECT 0.000 3096.005 208.285 3096.845 ;
      LAYER met2 ;
        RECT 210.370 3096.565 210.650 3096.585 ;
        RECT 208.565 3096.285 210.965 3096.565 ;
        RECT 209.400 3096.265 210.965 3096.285 ;
        RECT 210.370 3096.245 210.650 3096.265 ;
        RECT 212.370 3096.245 212.650 3136.305 ;
        RECT 213.960 3128.425 214.210 3343.085 ;
        RECT 214.460 3290.975 214.710 3506.635 ;
        RECT 214.960 3306.165 215.210 3521.825 ;
        RECT 3369.830 3464.185 3370.080 3688.845 ;
        RECT 3370.330 3479.365 3370.580 3704.025 ;
        RECT 3370.830 3651.925 3371.080 3876.585 ;
        RECT 3374.290 3867.385 3374.570 3907.405 ;
      LAYER met2 ;
        RECT 3379.715 3907.155 3588.000 3907.995 ;
        RECT 3379.435 3904.775 3588.000 3907.155 ;
        RECT 3379.715 3903.935 3588.000 3904.775 ;
        RECT 3379.435 3902.015 3588.000 3903.935 ;
        RECT 3379.715 3901.175 3588.000 3902.015 ;
        RECT 3379.435 3898.795 3588.000 3901.175 ;
        RECT 3379.715 3897.955 3588.000 3898.795 ;
        RECT 3379.435 3895.575 3588.000 3897.955 ;
        RECT 3379.715 3894.735 3588.000 3895.575 ;
        RECT 3379.435 3892.815 3588.000 3894.735 ;
        RECT 3379.715 3891.975 3588.000 3892.815 ;
        RECT 3379.435 3889.595 3588.000 3891.975 ;
        RECT 3379.715 3888.755 3588.000 3889.595 ;
        RECT 3379.435 3886.375 3588.000 3888.755 ;
      LAYER met2 ;
        RECT 3377.035 3885.815 3379.435 3886.095 ;
      LAYER met2 ;
        RECT 3379.715 3885.535 3588.000 3886.375 ;
        RECT 3379.435 3883.615 3588.000 3885.535 ;
        RECT 3379.715 3882.775 3588.000 3883.615 ;
        RECT 3379.435 3880.395 3588.000 3882.775 ;
        RECT 3379.715 3879.555 3588.000 3880.395 ;
        RECT 3379.435 3877.175 3588.000 3879.555 ;
      LAYER met2 ;
        RECT 3377.035 3876.615 3379.435 3876.895 ;
      LAYER met2 ;
        RECT 3379.715 3876.335 3588.000 3877.175 ;
        RECT 3379.435 3874.415 3588.000 3876.335 ;
      LAYER met2 ;
        RECT 3377.035 3873.855 3379.435 3874.135 ;
      LAYER met2 ;
        RECT 3379.715 3873.575 3588.000 3874.415 ;
        RECT 3379.435 3871.195 3588.000 3873.575 ;
        RECT 3379.715 3870.355 3588.000 3871.195 ;
        RECT 3379.435 3867.975 3588.000 3870.355 ;
      LAYER met2 ;
        RECT 3377.525 3867.695 3377.785 3867.705 ;
        RECT 3377.035 3867.415 3379.435 3867.695 ;
        RECT 3377.525 3867.385 3377.785 3867.415 ;
      LAYER met2 ;
        RECT 3379.715 3867.135 3588.000 3867.975 ;
        RECT 3379.435 3866.085 3588.000 3867.135 ;
        RECT 3379.435 3719.795 3588.000 3720.790 ;
        RECT 3379.715 3718.955 3588.000 3719.795 ;
        RECT 3379.435 3717.035 3588.000 3718.955 ;
        RECT 3379.715 3716.195 3588.000 3717.035 ;
        RECT 3379.435 3713.815 3588.000 3716.195 ;
        RECT 3379.715 3712.975 3588.000 3713.815 ;
        RECT 3379.435 3710.595 3588.000 3712.975 ;
        RECT 3379.715 3709.755 3588.000 3710.595 ;
        RECT 3379.435 3707.835 3588.000 3709.755 ;
        RECT 3379.715 3706.995 3588.000 3707.835 ;
        RECT 3379.435 3704.615 3588.000 3706.995 ;
      LAYER met2 ;
        RECT 3377.035 3704.055 3379.435 3704.335 ;
      LAYER met2 ;
        RECT 3379.715 3703.775 3588.000 3704.615 ;
        RECT 3379.435 3701.395 3588.000 3703.775 ;
        RECT 3379.715 3700.555 3588.000 3701.395 ;
        RECT 3379.435 3698.635 3588.000 3700.555 ;
        RECT 3379.715 3697.795 3588.000 3698.635 ;
        RECT 3379.435 3695.415 3588.000 3697.795 ;
        RECT 3379.715 3694.575 3588.000 3695.415 ;
        RECT 3379.435 3692.195 3588.000 3694.575 ;
        RECT 3379.715 3691.355 3588.000 3692.195 ;
        RECT 3379.435 3689.435 3588.000 3691.355 ;
      LAYER met2 ;
        RECT 3377.035 3688.875 3379.435 3689.155 ;
      LAYER met2 ;
        RECT 3379.715 3688.595 3588.000 3689.435 ;
        RECT 3379.435 3686.215 3588.000 3688.595 ;
        RECT 3379.715 3685.375 3588.000 3686.215 ;
        RECT 3379.435 3682.995 3588.000 3685.375 ;
      LAYER met2 ;
        RECT 3375.290 3682.745 3375.570 3682.840 ;
        RECT 3375.255 3682.405 3375.570 3682.745 ;
        RECT 3377.035 3682.435 3379.435 3682.715 ;
        RECT 3370.830 3651.585 3371.130 3651.925 ;
        RECT 3370.330 3479.025 3370.640 3479.365 ;
        RECT 3369.805 3463.845 3370.105 3464.185 ;
        RECT 214.955 3305.825 215.235 3306.165 ;
        RECT 214.430 3290.635 214.710 3290.975 ;
        RECT 213.920 3128.085 214.210 3128.425 ;
      LAYER met2 ;
        RECT 0.000 3093.625 208.565 3096.005 ;
        RECT 0.000 3092.785 208.285 3093.625 ;
        RECT 0.000 3090.405 208.565 3092.785 ;
        RECT 0.000 3089.565 208.285 3090.405 ;
      LAYER met2 ;
        RECT 210.370 3090.135 210.650 3090.165 ;
        RECT 210.145 3090.125 210.965 3090.135 ;
        RECT 208.565 3089.845 210.965 3090.125 ;
        RECT 210.370 3089.825 210.650 3089.845 ;
      LAYER met2 ;
        RECT 0.000 3087.645 208.565 3089.565 ;
        RECT 0.000 3086.805 208.285 3087.645 ;
        RECT 0.000 3084.425 208.565 3086.805 ;
        RECT 0.000 3083.585 208.285 3084.425 ;
        RECT 0.000 3081.205 208.565 3083.585 ;
        RECT 0.000 3080.365 208.285 3081.205 ;
        RECT 0.000 3078.445 208.565 3080.365 ;
        RECT 0.000 3077.605 208.285 3078.445 ;
        RECT 0.000 3075.225 208.565 3077.605 ;
        RECT 0.000 3074.385 208.285 3075.225 ;
      LAYER met2 ;
        RECT 210.370 3074.945 210.650 3074.975 ;
        RECT 208.565 3074.665 210.965 3074.945 ;
        RECT 210.370 3074.635 210.650 3074.665 ;
      LAYER met2 ;
        RECT 0.000 3072.005 208.565 3074.385 ;
        RECT 0.000 3071.165 208.285 3072.005 ;
        RECT 0.000 3069.245 208.565 3071.165 ;
        RECT 0.000 3068.405 208.285 3069.245 ;
        RECT 0.000 3066.025 208.565 3068.405 ;
        RECT 0.000 3065.185 208.285 3066.025 ;
        RECT 0.000 3062.805 208.565 3065.185 ;
        RECT 0.000 3061.965 208.285 3062.805 ;
        RECT 0.000 3060.045 208.565 3061.965 ;
        RECT 0.000 3059.205 208.285 3060.045 ;
        RECT 0.000 3058.210 208.565 3059.205 ;
        RECT 0.000 2920.865 208.565 2921.915 ;
        RECT 0.000 2920.025 208.285 2920.865 ;
      LAYER met2 ;
        RECT 212.070 2920.645 212.350 2920.720 ;
        RECT 210.370 2920.625 210.650 2920.645 ;
        RECT 209.945 2920.605 210.965 2920.625 ;
        RECT 209.910 2920.585 210.965 2920.605 ;
        RECT 208.565 2920.305 210.965 2920.585 ;
        RECT 212.070 2920.305 212.365 2920.645 ;
      LAYER met2 ;
        RECT 0.000 2917.645 208.565 2920.025 ;
        RECT 0.000 2916.805 208.285 2917.645 ;
        RECT 0.000 2914.425 208.565 2916.805 ;
        RECT 0.000 2913.585 208.285 2914.425 ;
      LAYER met2 ;
        RECT 208.565 2913.865 210.965 2914.145 ;
      LAYER met2 ;
        RECT 0.000 2911.665 208.565 2913.585 ;
        RECT 0.000 2910.825 208.285 2911.665 ;
      LAYER met2 ;
        RECT 210.525 2911.385 210.805 2912.440 ;
        RECT 208.565 2911.105 210.965 2911.385 ;
      LAYER met2 ;
        RECT 0.000 2908.445 208.565 2910.825 ;
        RECT 0.000 2907.605 208.285 2908.445 ;
        RECT 0.000 2905.225 208.565 2907.605 ;
        RECT 0.000 2904.385 208.285 2905.225 ;
        RECT 0.000 2902.465 208.565 2904.385 ;
        RECT 0.000 2901.625 208.285 2902.465 ;
      LAYER met2 ;
        RECT 208.565 2901.905 210.965 2902.185 ;
      LAYER met2 ;
        RECT 0.000 2899.245 208.565 2901.625 ;
        RECT 0.000 2898.405 208.285 2899.245 ;
        RECT 0.000 2896.025 208.565 2898.405 ;
        RECT 0.000 2895.185 208.285 2896.025 ;
        RECT 0.000 2893.265 208.565 2895.185 ;
        RECT 0.000 2892.425 208.285 2893.265 ;
        RECT 0.000 2890.045 208.565 2892.425 ;
        RECT 0.000 2889.205 208.285 2890.045 ;
        RECT 0.000 2886.825 208.565 2889.205 ;
        RECT 0.000 2885.985 208.285 2886.825 ;
        RECT 0.000 2884.065 208.565 2885.985 ;
        RECT 0.000 2883.225 208.285 2884.065 ;
        RECT 0.000 2880.845 208.565 2883.225 ;
        RECT 0.000 2880.005 208.285 2880.845 ;
      LAYER met2 ;
        RECT 210.370 2880.565 210.650 2880.585 ;
        RECT 208.565 2880.285 210.965 2880.565 ;
        RECT 209.400 2880.265 210.965 2880.285 ;
        RECT 210.370 2880.245 210.650 2880.265 ;
        RECT 212.070 2880.245 212.350 2920.305 ;
        RECT 213.960 2912.425 214.210 3128.085 ;
        RECT 214.460 3074.975 214.710 3290.635 ;
        RECT 214.960 3090.165 215.210 3305.825 ;
        RECT 3369.830 3238.185 3370.080 3463.845 ;
        RECT 3370.330 3253.365 3370.580 3479.025 ;
        RECT 3370.830 3426.925 3371.080 3651.585 ;
        RECT 3375.290 3642.385 3375.570 3682.405 ;
      LAYER met2 ;
        RECT 3379.715 3682.155 3588.000 3682.995 ;
        RECT 3379.435 3679.775 3588.000 3682.155 ;
        RECT 3379.715 3678.935 3588.000 3679.775 ;
        RECT 3379.435 3677.015 3588.000 3678.935 ;
        RECT 3379.715 3676.175 3588.000 3677.015 ;
        RECT 3379.435 3673.795 3588.000 3676.175 ;
        RECT 3379.715 3672.955 3588.000 3673.795 ;
        RECT 3379.435 3670.575 3588.000 3672.955 ;
        RECT 3379.715 3669.735 3588.000 3670.575 ;
        RECT 3379.435 3667.815 3588.000 3669.735 ;
        RECT 3379.715 3666.975 3588.000 3667.815 ;
        RECT 3379.435 3664.595 3588.000 3666.975 ;
        RECT 3379.715 3663.755 3588.000 3664.595 ;
        RECT 3379.435 3661.375 3588.000 3663.755 ;
      LAYER met2 ;
        RECT 3377.035 3660.815 3379.435 3661.095 ;
      LAYER met2 ;
        RECT 3379.715 3660.535 3588.000 3661.375 ;
        RECT 3379.435 3658.615 3588.000 3660.535 ;
        RECT 3379.715 3657.775 3588.000 3658.615 ;
        RECT 3379.435 3655.395 3588.000 3657.775 ;
        RECT 3379.715 3654.555 3588.000 3655.395 ;
        RECT 3379.435 3652.175 3588.000 3654.555 ;
      LAYER met2 ;
        RECT 3377.035 3651.615 3379.435 3651.895 ;
      LAYER met2 ;
        RECT 3379.715 3651.335 3588.000 3652.175 ;
        RECT 3379.435 3649.415 3588.000 3651.335 ;
      LAYER met2 ;
        RECT 3377.035 3648.855 3379.435 3649.135 ;
      LAYER met2 ;
        RECT 3379.715 3648.575 3588.000 3649.415 ;
        RECT 3379.435 3646.195 3588.000 3648.575 ;
        RECT 3379.715 3645.355 3588.000 3646.195 ;
        RECT 3379.435 3642.975 3588.000 3645.355 ;
      LAYER met2 ;
        RECT 3377.525 3642.695 3377.785 3642.705 ;
        RECT 3377.035 3642.415 3379.435 3642.695 ;
        RECT 3377.525 3642.385 3377.785 3642.415 ;
      LAYER met2 ;
        RECT 3379.715 3642.135 3588.000 3642.975 ;
        RECT 3379.435 3641.085 3588.000 3642.135 ;
        RECT 3379.435 3494.795 3588.000 3495.790 ;
        RECT 3379.715 3493.955 3588.000 3494.795 ;
        RECT 3379.435 3492.035 3588.000 3493.955 ;
        RECT 3379.715 3491.195 3588.000 3492.035 ;
        RECT 3379.435 3488.815 3588.000 3491.195 ;
        RECT 3379.715 3487.975 3588.000 3488.815 ;
        RECT 3379.435 3485.595 3588.000 3487.975 ;
        RECT 3379.715 3484.755 3588.000 3485.595 ;
        RECT 3379.435 3482.835 3588.000 3484.755 ;
        RECT 3379.715 3481.995 3588.000 3482.835 ;
        RECT 3379.435 3479.615 3588.000 3481.995 ;
      LAYER met2 ;
        RECT 3377.035 3479.055 3379.435 3479.335 ;
      LAYER met2 ;
        RECT 3379.715 3478.775 3588.000 3479.615 ;
        RECT 3379.435 3476.395 3588.000 3478.775 ;
        RECT 3379.715 3475.555 3588.000 3476.395 ;
        RECT 3379.435 3473.635 3588.000 3475.555 ;
        RECT 3379.715 3472.795 3588.000 3473.635 ;
        RECT 3379.435 3470.415 3588.000 3472.795 ;
        RECT 3379.715 3469.575 3588.000 3470.415 ;
        RECT 3379.435 3467.195 3588.000 3469.575 ;
        RECT 3379.715 3466.355 3588.000 3467.195 ;
        RECT 3379.435 3464.435 3588.000 3466.355 ;
      LAYER met2 ;
        RECT 3377.035 3463.875 3379.435 3464.155 ;
      LAYER met2 ;
        RECT 3379.715 3463.595 3588.000 3464.435 ;
        RECT 3379.435 3461.215 3588.000 3463.595 ;
        RECT 3379.715 3460.375 3588.000 3461.215 ;
        RECT 3379.435 3457.995 3588.000 3460.375 ;
      LAYER met2 ;
        RECT 3374.290 3457.745 3374.570 3457.840 ;
        RECT 3374.255 3457.405 3374.570 3457.745 ;
        RECT 3377.035 3457.435 3379.435 3457.715 ;
        RECT 3370.830 3426.585 3371.130 3426.925 ;
        RECT 3370.330 3253.025 3370.640 3253.365 ;
        RECT 3369.805 3237.845 3370.105 3238.185 ;
        RECT 214.955 3089.825 215.235 3090.165 ;
        RECT 214.430 3074.635 214.710 3074.975 ;
        RECT 213.920 2912.085 214.210 2912.425 ;
      LAYER met2 ;
        RECT 0.000 2877.625 208.565 2880.005 ;
        RECT 0.000 2876.785 208.285 2877.625 ;
        RECT 0.000 2874.405 208.565 2876.785 ;
        RECT 0.000 2873.565 208.285 2874.405 ;
      LAYER met2 ;
        RECT 210.370 2874.135 210.650 2874.165 ;
        RECT 210.145 2874.125 210.965 2874.135 ;
        RECT 208.565 2873.845 210.965 2874.125 ;
        RECT 210.370 2873.825 210.650 2873.845 ;
      LAYER met2 ;
        RECT 0.000 2871.645 208.565 2873.565 ;
        RECT 0.000 2870.805 208.285 2871.645 ;
        RECT 0.000 2868.425 208.565 2870.805 ;
        RECT 0.000 2867.585 208.285 2868.425 ;
        RECT 0.000 2865.205 208.565 2867.585 ;
        RECT 0.000 2864.365 208.285 2865.205 ;
        RECT 0.000 2862.445 208.565 2864.365 ;
        RECT 0.000 2861.605 208.285 2862.445 ;
        RECT 0.000 2859.225 208.565 2861.605 ;
        RECT 0.000 2858.385 208.285 2859.225 ;
      LAYER met2 ;
        RECT 210.370 2858.945 210.650 2858.975 ;
        RECT 208.565 2858.665 210.965 2858.945 ;
        RECT 210.370 2858.635 210.650 2858.665 ;
      LAYER met2 ;
        RECT 0.000 2856.005 208.565 2858.385 ;
        RECT 0.000 2855.165 208.285 2856.005 ;
        RECT 0.000 2853.245 208.565 2855.165 ;
        RECT 0.000 2852.405 208.285 2853.245 ;
        RECT 0.000 2850.025 208.565 2852.405 ;
        RECT 0.000 2849.185 208.285 2850.025 ;
        RECT 0.000 2846.805 208.565 2849.185 ;
        RECT 0.000 2845.965 208.285 2846.805 ;
        RECT 0.000 2844.045 208.565 2845.965 ;
        RECT 0.000 2843.205 208.285 2844.045 ;
        RECT 0.000 2842.210 208.565 2843.205 ;
        RECT 0.000 2704.865 208.565 2705.915 ;
        RECT 0.000 2704.025 208.285 2704.865 ;
      LAYER met2 ;
        RECT 211.970 2704.645 212.250 2704.720 ;
        RECT 210.370 2704.625 210.650 2704.645 ;
        RECT 209.945 2704.605 210.965 2704.625 ;
        RECT 209.910 2704.585 210.965 2704.605 ;
        RECT 208.565 2704.305 210.965 2704.585 ;
        RECT 211.970 2704.305 212.265 2704.645 ;
      LAYER met2 ;
        RECT 0.000 2701.645 208.565 2704.025 ;
        RECT 0.000 2700.805 208.285 2701.645 ;
        RECT 0.000 2698.425 208.565 2700.805 ;
        RECT 0.000 2697.585 208.285 2698.425 ;
      LAYER met2 ;
        RECT 208.565 2697.865 210.965 2698.145 ;
      LAYER met2 ;
        RECT 0.000 2695.665 208.565 2697.585 ;
        RECT 0.000 2694.825 208.285 2695.665 ;
      LAYER met2 ;
        RECT 210.370 2695.405 210.650 2695.425 ;
        RECT 209.945 2695.385 210.965 2695.405 ;
        RECT 208.565 2695.105 210.965 2695.385 ;
        RECT 210.370 2695.085 210.650 2695.105 ;
      LAYER met2 ;
        RECT 0.000 2692.445 208.565 2694.825 ;
        RECT 0.000 2691.605 208.285 2692.445 ;
        RECT 0.000 2689.225 208.565 2691.605 ;
        RECT 0.000 2688.385 208.285 2689.225 ;
        RECT 0.000 2686.465 208.565 2688.385 ;
        RECT 0.000 2685.625 208.285 2686.465 ;
      LAYER met2 ;
        RECT 208.565 2685.905 210.965 2686.185 ;
      LAYER met2 ;
        RECT 0.000 2683.245 208.565 2685.625 ;
        RECT 0.000 2682.405 208.285 2683.245 ;
        RECT 0.000 2680.025 208.565 2682.405 ;
        RECT 0.000 2679.185 208.285 2680.025 ;
        RECT 0.000 2677.265 208.565 2679.185 ;
        RECT 0.000 2676.425 208.285 2677.265 ;
        RECT 0.000 2674.045 208.565 2676.425 ;
        RECT 0.000 2673.205 208.285 2674.045 ;
        RECT 0.000 2670.825 208.565 2673.205 ;
        RECT 0.000 2669.985 208.285 2670.825 ;
        RECT 0.000 2668.065 208.565 2669.985 ;
        RECT 0.000 2667.225 208.285 2668.065 ;
        RECT 0.000 2664.845 208.565 2667.225 ;
        RECT 0.000 2664.005 208.285 2664.845 ;
      LAYER met2 ;
        RECT 210.370 2664.565 210.650 2664.585 ;
        RECT 208.565 2664.285 210.965 2664.565 ;
        RECT 209.400 2664.265 210.965 2664.285 ;
        RECT 210.370 2664.245 210.650 2664.265 ;
        RECT 211.970 2664.245 212.250 2704.305 ;
        RECT 213.960 2695.425 214.210 2912.085 ;
        RECT 214.460 2858.975 214.710 3074.635 ;
        RECT 214.960 2874.165 215.210 3089.825 ;
        RECT 3369.830 3013.185 3370.080 3237.845 ;
        RECT 3370.330 3028.365 3370.580 3253.025 ;
        RECT 3370.830 3200.925 3371.080 3426.585 ;
        RECT 3374.290 3417.385 3374.570 3457.405 ;
      LAYER met2 ;
        RECT 3379.715 3457.155 3588.000 3457.995 ;
        RECT 3379.435 3454.775 3588.000 3457.155 ;
        RECT 3379.715 3453.935 3588.000 3454.775 ;
        RECT 3379.435 3452.015 3588.000 3453.935 ;
        RECT 3379.715 3451.175 3588.000 3452.015 ;
        RECT 3379.435 3448.795 3588.000 3451.175 ;
        RECT 3379.715 3447.955 3588.000 3448.795 ;
        RECT 3379.435 3445.575 3588.000 3447.955 ;
        RECT 3379.715 3444.735 3588.000 3445.575 ;
        RECT 3379.435 3442.815 3588.000 3444.735 ;
        RECT 3379.715 3441.975 3588.000 3442.815 ;
        RECT 3379.435 3439.595 3588.000 3441.975 ;
        RECT 3379.715 3438.755 3588.000 3439.595 ;
        RECT 3379.435 3436.375 3588.000 3438.755 ;
      LAYER met2 ;
        RECT 3377.035 3435.815 3379.435 3436.095 ;
      LAYER met2 ;
        RECT 3379.715 3435.535 3588.000 3436.375 ;
        RECT 3379.435 3433.615 3588.000 3435.535 ;
        RECT 3379.715 3432.775 3588.000 3433.615 ;
        RECT 3379.435 3430.395 3588.000 3432.775 ;
        RECT 3379.715 3429.555 3588.000 3430.395 ;
        RECT 3379.435 3427.175 3588.000 3429.555 ;
      LAYER met2 ;
        RECT 3377.035 3426.615 3379.435 3426.895 ;
      LAYER met2 ;
        RECT 3379.715 3426.335 3588.000 3427.175 ;
        RECT 3379.435 3424.415 3588.000 3426.335 ;
      LAYER met2 ;
        RECT 3377.035 3423.855 3379.435 3424.135 ;
      LAYER met2 ;
        RECT 3379.715 3423.575 3588.000 3424.415 ;
        RECT 3379.435 3421.195 3588.000 3423.575 ;
        RECT 3379.715 3420.355 3588.000 3421.195 ;
        RECT 3379.435 3417.975 3588.000 3420.355 ;
      LAYER met2 ;
        RECT 3377.525 3417.695 3377.785 3417.705 ;
        RECT 3377.035 3417.415 3379.435 3417.695 ;
        RECT 3377.525 3417.385 3377.785 3417.415 ;
      LAYER met2 ;
        RECT 3379.715 3417.135 3588.000 3417.975 ;
        RECT 3379.435 3416.085 3588.000 3417.135 ;
        RECT 3379.435 3268.795 3588.000 3269.790 ;
        RECT 3379.715 3267.955 3588.000 3268.795 ;
        RECT 3379.435 3266.035 3588.000 3267.955 ;
        RECT 3379.715 3265.195 3588.000 3266.035 ;
        RECT 3379.435 3262.815 3588.000 3265.195 ;
        RECT 3379.715 3261.975 3588.000 3262.815 ;
        RECT 3379.435 3259.595 3588.000 3261.975 ;
        RECT 3379.715 3258.755 3588.000 3259.595 ;
        RECT 3379.435 3256.835 3588.000 3258.755 ;
        RECT 3379.715 3255.995 3588.000 3256.835 ;
        RECT 3379.435 3253.615 3588.000 3255.995 ;
      LAYER met2 ;
        RECT 3377.035 3253.055 3379.435 3253.335 ;
      LAYER met2 ;
        RECT 3379.715 3252.775 3588.000 3253.615 ;
        RECT 3379.435 3250.395 3588.000 3252.775 ;
        RECT 3379.715 3249.555 3588.000 3250.395 ;
        RECT 3379.435 3247.635 3588.000 3249.555 ;
        RECT 3379.715 3246.795 3588.000 3247.635 ;
        RECT 3379.435 3244.415 3588.000 3246.795 ;
        RECT 3379.715 3243.575 3588.000 3244.415 ;
        RECT 3379.435 3241.195 3588.000 3243.575 ;
        RECT 3379.715 3240.355 3588.000 3241.195 ;
        RECT 3379.435 3238.435 3588.000 3240.355 ;
      LAYER met2 ;
        RECT 3377.035 3237.875 3379.435 3238.155 ;
      LAYER met2 ;
        RECT 3379.715 3237.595 3588.000 3238.435 ;
        RECT 3379.435 3235.215 3588.000 3237.595 ;
        RECT 3379.715 3234.375 3588.000 3235.215 ;
        RECT 3379.435 3231.995 3588.000 3234.375 ;
      LAYER met2 ;
        RECT 3374.290 3231.745 3374.570 3231.840 ;
        RECT 3374.255 3231.405 3374.570 3231.745 ;
        RECT 3377.035 3231.435 3379.435 3231.715 ;
        RECT 3370.830 3200.585 3371.130 3200.925 ;
        RECT 3370.330 3028.025 3370.640 3028.365 ;
        RECT 3369.805 3012.845 3370.105 3013.185 ;
        RECT 214.955 2873.825 215.235 2874.165 ;
        RECT 214.430 2858.635 214.710 2858.975 ;
        RECT 213.920 2695.085 214.210 2695.425 ;
      LAYER met2 ;
        RECT 0.000 2661.625 208.565 2664.005 ;
        RECT 0.000 2660.785 208.285 2661.625 ;
        RECT 0.000 2658.405 208.565 2660.785 ;
        RECT 0.000 2657.565 208.285 2658.405 ;
      LAYER met2 ;
        RECT 210.370 2658.135 210.650 2658.165 ;
        RECT 210.145 2658.125 210.965 2658.135 ;
        RECT 208.565 2657.845 210.965 2658.125 ;
        RECT 210.370 2657.825 210.650 2657.845 ;
      LAYER met2 ;
        RECT 0.000 2655.645 208.565 2657.565 ;
        RECT 0.000 2654.805 208.285 2655.645 ;
        RECT 0.000 2652.425 208.565 2654.805 ;
        RECT 0.000 2651.585 208.285 2652.425 ;
        RECT 0.000 2649.205 208.565 2651.585 ;
        RECT 0.000 2648.365 208.285 2649.205 ;
        RECT 0.000 2646.445 208.565 2648.365 ;
        RECT 0.000 2645.605 208.285 2646.445 ;
        RECT 0.000 2643.225 208.565 2645.605 ;
        RECT 0.000 2642.385 208.285 2643.225 ;
      LAYER met2 ;
        RECT 210.370 2642.945 210.650 2642.975 ;
        RECT 208.565 2642.665 210.965 2642.945 ;
        RECT 210.370 2642.635 210.650 2642.665 ;
      LAYER met2 ;
        RECT 0.000 2640.005 208.565 2642.385 ;
        RECT 0.000 2639.165 208.285 2640.005 ;
        RECT 0.000 2637.245 208.565 2639.165 ;
        RECT 0.000 2636.405 208.285 2637.245 ;
        RECT 0.000 2634.025 208.565 2636.405 ;
        RECT 0.000 2633.185 208.285 2634.025 ;
        RECT 0.000 2630.805 208.565 2633.185 ;
        RECT 0.000 2629.965 208.285 2630.805 ;
        RECT 0.000 2628.045 208.565 2629.965 ;
        RECT 0.000 2627.205 208.285 2628.045 ;
        RECT 0.000 2626.210 208.565 2627.205 ;
        RECT 4.925 2465.390 200.000 2489.290 ;
        RECT 4.925 2439.395 197.965 2465.390 ;
        RECT 198.080 2440.895 200.000 2442.895 ;
        RECT 4.925 2415.495 200.000 2439.395 ;
        RECT 4.925 2415.265 197.965 2415.495 ;
        RECT 0.000 2066.865 208.565 2067.915 ;
        RECT 0.000 2066.025 208.285 2066.865 ;
      LAYER met2 ;
        RECT 212.370 2066.645 212.650 2066.720 ;
        RECT 210.370 2066.625 210.650 2066.645 ;
        RECT 209.945 2066.605 210.965 2066.625 ;
        RECT 209.910 2066.585 210.965 2066.605 ;
        RECT 208.565 2066.305 210.965 2066.585 ;
        RECT 212.370 2066.305 212.665 2066.645 ;
      LAYER met2 ;
        RECT 0.000 2063.645 208.565 2066.025 ;
        RECT 0.000 2062.805 208.285 2063.645 ;
        RECT 0.000 2060.425 208.565 2062.805 ;
        RECT 0.000 2059.585 208.285 2060.425 ;
      LAYER met2 ;
        RECT 208.565 2059.865 210.965 2060.145 ;
      LAYER met2 ;
        RECT 0.000 2057.665 208.565 2059.585 ;
        RECT 0.000 2056.825 208.285 2057.665 ;
      LAYER met2 ;
        RECT 210.370 2057.405 210.650 2057.425 ;
        RECT 209.945 2057.385 210.965 2057.405 ;
        RECT 208.565 2057.105 210.965 2057.385 ;
        RECT 210.370 2057.085 210.650 2057.105 ;
      LAYER met2 ;
        RECT 0.000 2054.445 208.565 2056.825 ;
        RECT 0.000 2053.605 208.285 2054.445 ;
        RECT 0.000 2051.225 208.565 2053.605 ;
        RECT 0.000 2050.385 208.285 2051.225 ;
        RECT 0.000 2048.465 208.565 2050.385 ;
        RECT 0.000 2047.625 208.285 2048.465 ;
      LAYER met2 ;
        RECT 208.565 2047.905 210.965 2048.185 ;
      LAYER met2 ;
        RECT 0.000 2045.245 208.565 2047.625 ;
        RECT 0.000 2044.405 208.285 2045.245 ;
        RECT 0.000 2042.025 208.565 2044.405 ;
        RECT 0.000 2041.185 208.285 2042.025 ;
        RECT 0.000 2039.265 208.565 2041.185 ;
        RECT 0.000 2038.425 208.285 2039.265 ;
        RECT 0.000 2036.045 208.565 2038.425 ;
        RECT 0.000 2035.205 208.285 2036.045 ;
        RECT 0.000 2032.825 208.565 2035.205 ;
        RECT 0.000 2031.985 208.285 2032.825 ;
        RECT 0.000 2030.065 208.565 2031.985 ;
        RECT 0.000 2029.225 208.285 2030.065 ;
        RECT 0.000 2026.845 208.565 2029.225 ;
        RECT 0.000 2026.005 208.285 2026.845 ;
      LAYER met2 ;
        RECT 210.370 2026.565 210.650 2026.585 ;
        RECT 208.565 2026.285 210.965 2026.565 ;
        RECT 209.400 2026.265 210.965 2026.285 ;
        RECT 210.370 2026.245 210.650 2026.265 ;
        RECT 212.370 2026.245 212.650 2066.305 ;
        RECT 213.960 2057.425 214.210 2695.085 ;
        RECT 214.460 2642.975 214.710 2858.635 ;
        RECT 214.960 2658.165 215.210 2873.825 ;
        RECT 3369.830 2787.185 3370.080 3012.845 ;
        RECT 3370.330 2802.365 3370.580 3028.025 ;
        RECT 3370.830 2975.925 3371.080 3200.585 ;
        RECT 3374.290 3191.385 3374.570 3231.405 ;
      LAYER met2 ;
        RECT 3379.715 3231.155 3588.000 3231.995 ;
        RECT 3379.435 3228.775 3588.000 3231.155 ;
        RECT 3379.715 3227.935 3588.000 3228.775 ;
        RECT 3379.435 3226.015 3588.000 3227.935 ;
        RECT 3379.715 3225.175 3588.000 3226.015 ;
        RECT 3379.435 3222.795 3588.000 3225.175 ;
        RECT 3379.715 3221.955 3588.000 3222.795 ;
        RECT 3379.435 3219.575 3588.000 3221.955 ;
        RECT 3379.715 3218.735 3588.000 3219.575 ;
        RECT 3379.435 3216.815 3588.000 3218.735 ;
        RECT 3379.715 3215.975 3588.000 3216.815 ;
        RECT 3379.435 3213.595 3588.000 3215.975 ;
        RECT 3379.715 3212.755 3588.000 3213.595 ;
        RECT 3379.435 3210.375 3588.000 3212.755 ;
      LAYER met2 ;
        RECT 3377.035 3209.815 3379.435 3210.095 ;
      LAYER met2 ;
        RECT 3379.715 3209.535 3588.000 3210.375 ;
        RECT 3379.435 3207.615 3588.000 3209.535 ;
        RECT 3379.715 3206.775 3588.000 3207.615 ;
        RECT 3379.435 3204.395 3588.000 3206.775 ;
        RECT 3379.715 3203.555 3588.000 3204.395 ;
        RECT 3379.435 3201.175 3588.000 3203.555 ;
      LAYER met2 ;
        RECT 3377.035 3200.615 3379.435 3200.895 ;
      LAYER met2 ;
        RECT 3379.715 3200.335 3588.000 3201.175 ;
        RECT 3379.435 3198.415 3588.000 3200.335 ;
      LAYER met2 ;
        RECT 3377.035 3197.855 3379.435 3198.135 ;
      LAYER met2 ;
        RECT 3379.715 3197.575 3588.000 3198.415 ;
        RECT 3379.435 3195.195 3588.000 3197.575 ;
        RECT 3379.715 3194.355 3588.000 3195.195 ;
        RECT 3379.435 3191.975 3588.000 3194.355 ;
      LAYER met2 ;
        RECT 3377.525 3191.695 3377.785 3191.705 ;
        RECT 3377.035 3191.415 3379.435 3191.695 ;
        RECT 3377.525 3191.385 3377.785 3191.415 ;
      LAYER met2 ;
        RECT 3379.715 3191.135 3588.000 3191.975 ;
        RECT 3379.435 3190.085 3588.000 3191.135 ;
        RECT 3379.435 3043.795 3588.000 3044.790 ;
        RECT 3379.715 3042.955 3588.000 3043.795 ;
        RECT 3379.435 3041.035 3588.000 3042.955 ;
        RECT 3379.715 3040.195 3588.000 3041.035 ;
        RECT 3379.435 3037.815 3588.000 3040.195 ;
        RECT 3379.715 3036.975 3588.000 3037.815 ;
        RECT 3379.435 3034.595 3588.000 3036.975 ;
        RECT 3379.715 3033.755 3588.000 3034.595 ;
        RECT 3379.435 3031.835 3588.000 3033.755 ;
        RECT 3379.715 3030.995 3588.000 3031.835 ;
        RECT 3379.435 3028.615 3588.000 3030.995 ;
      LAYER met2 ;
        RECT 3377.035 3028.055 3379.435 3028.335 ;
      LAYER met2 ;
        RECT 3379.715 3027.775 3588.000 3028.615 ;
        RECT 3379.435 3025.395 3588.000 3027.775 ;
        RECT 3379.715 3024.555 3588.000 3025.395 ;
        RECT 3379.435 3022.635 3588.000 3024.555 ;
        RECT 3379.715 3021.795 3588.000 3022.635 ;
        RECT 3379.435 3019.415 3588.000 3021.795 ;
        RECT 3379.715 3018.575 3588.000 3019.415 ;
        RECT 3379.435 3016.195 3588.000 3018.575 ;
        RECT 3379.715 3015.355 3588.000 3016.195 ;
        RECT 3379.435 3013.435 3588.000 3015.355 ;
      LAYER met2 ;
        RECT 3377.035 3012.875 3379.435 3013.155 ;
      LAYER met2 ;
        RECT 3379.715 3012.595 3588.000 3013.435 ;
        RECT 3379.435 3010.215 3588.000 3012.595 ;
        RECT 3379.715 3009.375 3588.000 3010.215 ;
        RECT 3379.435 3006.995 3588.000 3009.375 ;
      LAYER met2 ;
        RECT 3374.140 3006.745 3374.405 3006.840 ;
        RECT 3374.105 3006.405 3374.405 3006.745 ;
        RECT 3377.035 3006.435 3379.435 3006.715 ;
        RECT 3370.830 2975.585 3371.130 2975.925 ;
        RECT 3370.330 2802.025 3370.640 2802.365 ;
        RECT 3369.805 2786.845 3370.105 2787.185 ;
        RECT 214.955 2657.825 215.235 2658.165 ;
        RECT 214.430 2642.635 214.710 2642.975 ;
        RECT 213.920 2057.085 214.210 2057.425 ;
      LAYER met2 ;
        RECT 0.000 2023.625 208.565 2026.005 ;
        RECT 0.000 2022.785 208.285 2023.625 ;
        RECT 0.000 2020.405 208.565 2022.785 ;
        RECT 0.000 2019.565 208.285 2020.405 ;
      LAYER met2 ;
        RECT 210.370 2020.135 210.650 2020.165 ;
        RECT 210.145 2020.125 210.965 2020.135 ;
        RECT 208.565 2019.845 210.965 2020.125 ;
        RECT 210.370 2019.825 210.650 2019.845 ;
      LAYER met2 ;
        RECT 0.000 2017.645 208.565 2019.565 ;
        RECT 0.000 2016.805 208.285 2017.645 ;
        RECT 0.000 2014.425 208.565 2016.805 ;
        RECT 0.000 2013.585 208.285 2014.425 ;
        RECT 0.000 2011.205 208.565 2013.585 ;
        RECT 0.000 2010.365 208.285 2011.205 ;
        RECT 0.000 2008.445 208.565 2010.365 ;
        RECT 0.000 2007.605 208.285 2008.445 ;
        RECT 0.000 2005.225 208.565 2007.605 ;
        RECT 0.000 2004.385 208.285 2005.225 ;
      LAYER met2 ;
        RECT 210.370 2004.945 210.650 2004.975 ;
        RECT 208.565 2004.665 210.965 2004.945 ;
        RECT 210.370 2004.635 210.650 2004.665 ;
      LAYER met2 ;
        RECT 0.000 2002.005 208.565 2004.385 ;
        RECT 0.000 2001.165 208.285 2002.005 ;
        RECT 0.000 1999.245 208.565 2001.165 ;
        RECT 0.000 1998.405 208.285 1999.245 ;
        RECT 0.000 1996.025 208.565 1998.405 ;
        RECT 0.000 1995.185 208.285 1996.025 ;
        RECT 0.000 1992.805 208.565 1995.185 ;
        RECT 0.000 1991.965 208.285 1992.805 ;
        RECT 0.000 1990.045 208.565 1991.965 ;
        RECT 0.000 1989.205 208.285 1990.045 ;
        RECT 0.000 1988.210 208.565 1989.205 ;
        RECT 0.000 1850.865 208.565 1851.915 ;
        RECT 0.000 1850.025 208.285 1850.865 ;
      LAYER met2 ;
        RECT 212.370 1850.645 212.650 1850.720 ;
        RECT 210.370 1850.625 210.650 1850.645 ;
        RECT 209.945 1850.605 210.965 1850.625 ;
        RECT 209.910 1850.585 210.965 1850.605 ;
        RECT 208.565 1850.305 210.965 1850.585 ;
        RECT 212.370 1850.305 212.665 1850.645 ;
      LAYER met2 ;
        RECT 0.000 1847.645 208.565 1850.025 ;
        RECT 0.000 1846.805 208.285 1847.645 ;
        RECT 0.000 1844.425 208.565 1846.805 ;
        RECT 0.000 1843.585 208.285 1844.425 ;
      LAYER met2 ;
        RECT 208.565 1843.865 210.965 1844.145 ;
      LAYER met2 ;
        RECT 0.000 1841.665 208.565 1843.585 ;
        RECT 0.000 1840.825 208.285 1841.665 ;
      LAYER met2 ;
        RECT 210.370 1841.405 210.650 1841.425 ;
        RECT 209.945 1841.385 210.965 1841.405 ;
        RECT 208.565 1841.105 210.965 1841.385 ;
        RECT 210.370 1841.085 210.650 1841.105 ;
      LAYER met2 ;
        RECT 0.000 1838.445 208.565 1840.825 ;
        RECT 0.000 1837.605 208.285 1838.445 ;
        RECT 0.000 1835.225 208.565 1837.605 ;
        RECT 0.000 1834.385 208.285 1835.225 ;
        RECT 0.000 1832.465 208.565 1834.385 ;
        RECT 0.000 1831.625 208.285 1832.465 ;
      LAYER met2 ;
        RECT 208.565 1831.905 210.965 1832.185 ;
      LAYER met2 ;
        RECT 0.000 1829.245 208.565 1831.625 ;
        RECT 0.000 1828.405 208.285 1829.245 ;
        RECT 0.000 1826.025 208.565 1828.405 ;
        RECT 0.000 1825.185 208.285 1826.025 ;
        RECT 0.000 1823.265 208.565 1825.185 ;
        RECT 0.000 1822.425 208.285 1823.265 ;
        RECT 0.000 1820.045 208.565 1822.425 ;
        RECT 0.000 1819.205 208.285 1820.045 ;
        RECT 0.000 1816.825 208.565 1819.205 ;
        RECT 0.000 1815.985 208.285 1816.825 ;
        RECT 0.000 1814.065 208.565 1815.985 ;
        RECT 0.000 1813.225 208.285 1814.065 ;
        RECT 0.000 1810.845 208.565 1813.225 ;
        RECT 0.000 1810.005 208.285 1810.845 ;
      LAYER met2 ;
        RECT 210.370 1810.565 210.650 1810.585 ;
        RECT 208.565 1810.285 210.965 1810.565 ;
        RECT 209.400 1810.265 210.965 1810.285 ;
        RECT 210.370 1810.245 210.650 1810.265 ;
        RECT 212.370 1810.245 212.650 1850.305 ;
        RECT 213.960 1841.425 214.210 2057.085 ;
        RECT 214.460 2004.975 214.710 2642.635 ;
        RECT 214.960 2020.165 215.210 2657.825 ;
        RECT 214.955 2019.825 215.235 2020.165 ;
        RECT 214.430 2004.635 214.710 2004.975 ;
        RECT 213.920 1841.085 214.210 1841.425 ;
      LAYER met2 ;
        RECT 0.000 1807.625 208.565 1810.005 ;
        RECT 0.000 1806.785 208.285 1807.625 ;
        RECT 0.000 1804.405 208.565 1806.785 ;
        RECT 0.000 1803.565 208.285 1804.405 ;
      LAYER met2 ;
        RECT 210.370 1804.135 210.650 1804.165 ;
        RECT 210.145 1804.125 210.965 1804.135 ;
        RECT 208.565 1803.845 210.965 1804.125 ;
        RECT 210.370 1803.825 210.650 1803.845 ;
      LAYER met2 ;
        RECT 0.000 1801.645 208.565 1803.565 ;
        RECT 0.000 1800.805 208.285 1801.645 ;
        RECT 0.000 1798.425 208.565 1800.805 ;
        RECT 0.000 1797.585 208.285 1798.425 ;
        RECT 0.000 1795.205 208.565 1797.585 ;
        RECT 0.000 1794.365 208.285 1795.205 ;
        RECT 0.000 1792.445 208.565 1794.365 ;
        RECT 0.000 1791.605 208.285 1792.445 ;
        RECT 0.000 1789.225 208.565 1791.605 ;
        RECT 0.000 1788.385 208.285 1789.225 ;
      LAYER met2 ;
        RECT 210.370 1788.945 210.650 1788.975 ;
        RECT 208.565 1788.665 210.965 1788.945 ;
        RECT 210.370 1788.635 210.650 1788.665 ;
      LAYER met2 ;
        RECT 0.000 1786.005 208.565 1788.385 ;
        RECT 0.000 1785.165 208.285 1786.005 ;
        RECT 0.000 1783.245 208.565 1785.165 ;
        RECT 0.000 1782.405 208.285 1783.245 ;
        RECT 0.000 1780.025 208.565 1782.405 ;
        RECT 0.000 1779.185 208.285 1780.025 ;
        RECT 0.000 1776.805 208.565 1779.185 ;
        RECT 0.000 1775.965 208.285 1776.805 ;
        RECT 0.000 1774.045 208.565 1775.965 ;
        RECT 0.000 1773.205 208.285 1774.045 ;
        RECT 0.000 1772.210 208.565 1773.205 ;
        RECT 0.000 1634.865 208.565 1635.915 ;
        RECT 0.000 1634.025 208.285 1634.865 ;
      LAYER met2 ;
        RECT 212.370 1634.645 212.650 1634.720 ;
        RECT 210.370 1634.625 210.650 1634.645 ;
        RECT 209.945 1634.605 210.965 1634.625 ;
        RECT 209.910 1634.585 210.965 1634.605 ;
        RECT 208.565 1634.305 210.965 1634.585 ;
        RECT 212.370 1634.305 212.665 1634.645 ;
      LAYER met2 ;
        RECT 0.000 1631.645 208.565 1634.025 ;
        RECT 0.000 1630.805 208.285 1631.645 ;
        RECT 0.000 1628.425 208.565 1630.805 ;
        RECT 0.000 1627.585 208.285 1628.425 ;
      LAYER met2 ;
        RECT 208.565 1627.865 210.965 1628.145 ;
      LAYER met2 ;
        RECT 0.000 1625.665 208.565 1627.585 ;
        RECT 0.000 1624.825 208.285 1625.665 ;
      LAYER met2 ;
        RECT 210.370 1625.405 210.650 1625.425 ;
        RECT 209.945 1625.385 210.965 1625.405 ;
        RECT 208.565 1625.105 210.965 1625.385 ;
        RECT 210.370 1625.085 210.650 1625.105 ;
      LAYER met2 ;
        RECT 0.000 1622.445 208.565 1624.825 ;
        RECT 0.000 1621.605 208.285 1622.445 ;
        RECT 0.000 1619.225 208.565 1621.605 ;
        RECT 0.000 1618.385 208.285 1619.225 ;
        RECT 0.000 1616.465 208.565 1618.385 ;
        RECT 0.000 1615.625 208.285 1616.465 ;
      LAYER met2 ;
        RECT 208.565 1615.905 210.965 1616.185 ;
      LAYER met2 ;
        RECT 0.000 1613.245 208.565 1615.625 ;
        RECT 0.000 1612.405 208.285 1613.245 ;
        RECT 0.000 1610.025 208.565 1612.405 ;
        RECT 0.000 1609.185 208.285 1610.025 ;
        RECT 0.000 1607.265 208.565 1609.185 ;
        RECT 0.000 1606.425 208.285 1607.265 ;
        RECT 0.000 1604.045 208.565 1606.425 ;
        RECT 0.000 1603.205 208.285 1604.045 ;
        RECT 0.000 1600.825 208.565 1603.205 ;
        RECT 0.000 1599.985 208.285 1600.825 ;
        RECT 0.000 1598.065 208.565 1599.985 ;
        RECT 0.000 1597.225 208.285 1598.065 ;
        RECT 0.000 1594.845 208.565 1597.225 ;
        RECT 0.000 1594.005 208.285 1594.845 ;
      LAYER met2 ;
        RECT 210.370 1594.565 210.650 1594.585 ;
        RECT 208.565 1594.285 210.965 1594.565 ;
        RECT 209.400 1594.265 210.965 1594.285 ;
        RECT 210.370 1594.245 210.650 1594.265 ;
        RECT 212.370 1594.245 212.650 1634.305 ;
        RECT 213.960 1625.425 214.210 1841.085 ;
        RECT 214.460 1788.975 214.710 2004.635 ;
        RECT 214.960 1804.165 215.210 2019.825 ;
        RECT 3369.830 1901.185 3370.080 2786.845 ;
        RECT 3370.330 1916.365 3370.580 2802.025 ;
        RECT 3370.830 2749.925 3371.080 2975.585 ;
        RECT 3374.140 2966.385 3374.405 3006.405 ;
      LAYER met2 ;
        RECT 3379.715 3006.155 3588.000 3006.995 ;
        RECT 3379.435 3003.775 3588.000 3006.155 ;
        RECT 3379.715 3002.935 3588.000 3003.775 ;
        RECT 3379.435 3001.015 3588.000 3002.935 ;
        RECT 3379.715 3000.175 3588.000 3001.015 ;
        RECT 3379.435 2997.795 3588.000 3000.175 ;
        RECT 3379.715 2996.955 3588.000 2997.795 ;
        RECT 3379.435 2994.575 3588.000 2996.955 ;
        RECT 3379.715 2993.735 3588.000 2994.575 ;
        RECT 3379.435 2991.815 3588.000 2993.735 ;
        RECT 3379.715 2990.975 3588.000 2991.815 ;
        RECT 3379.435 2988.595 3588.000 2990.975 ;
        RECT 3379.715 2987.755 3588.000 2988.595 ;
        RECT 3379.435 2985.375 3588.000 2987.755 ;
      LAYER met2 ;
        RECT 3377.035 2984.815 3379.435 2985.095 ;
      LAYER met2 ;
        RECT 3379.715 2984.535 3588.000 2985.375 ;
        RECT 3379.435 2982.615 3588.000 2984.535 ;
        RECT 3379.715 2981.775 3588.000 2982.615 ;
        RECT 3379.435 2979.395 3588.000 2981.775 ;
        RECT 3379.715 2978.555 3588.000 2979.395 ;
        RECT 3379.435 2976.175 3588.000 2978.555 ;
      LAYER met2 ;
        RECT 3377.035 2975.615 3379.435 2975.895 ;
      LAYER met2 ;
        RECT 3379.715 2975.335 3588.000 2976.175 ;
        RECT 3379.435 2973.415 3588.000 2975.335 ;
      LAYER met2 ;
        RECT 3377.035 2972.855 3379.435 2973.135 ;
      LAYER met2 ;
        RECT 3379.715 2972.575 3588.000 2973.415 ;
        RECT 3379.435 2970.195 3588.000 2972.575 ;
        RECT 3379.715 2969.355 3588.000 2970.195 ;
        RECT 3379.435 2966.975 3588.000 2969.355 ;
      LAYER met2 ;
        RECT 3377.525 2966.695 3377.785 2966.705 ;
        RECT 3377.035 2966.415 3379.435 2966.695 ;
        RECT 3377.525 2966.385 3377.785 2966.415 ;
      LAYER met2 ;
        RECT 3379.715 2966.135 3588.000 2966.975 ;
        RECT 3379.435 2965.085 3588.000 2966.135 ;
        RECT 3379.435 2817.795 3588.000 2818.790 ;
        RECT 3379.715 2816.955 3588.000 2817.795 ;
        RECT 3379.435 2815.035 3588.000 2816.955 ;
        RECT 3379.715 2814.195 3588.000 2815.035 ;
        RECT 3379.435 2811.815 3588.000 2814.195 ;
        RECT 3379.715 2810.975 3588.000 2811.815 ;
        RECT 3379.435 2808.595 3588.000 2810.975 ;
        RECT 3379.715 2807.755 3588.000 2808.595 ;
        RECT 3379.435 2805.835 3588.000 2807.755 ;
        RECT 3379.715 2804.995 3588.000 2805.835 ;
        RECT 3379.435 2802.615 3588.000 2804.995 ;
      LAYER met2 ;
        RECT 3377.035 2802.055 3379.435 2802.335 ;
      LAYER met2 ;
        RECT 3379.715 2801.775 3588.000 2802.615 ;
        RECT 3379.435 2799.395 3588.000 2801.775 ;
        RECT 3379.715 2798.555 3588.000 2799.395 ;
        RECT 3379.435 2796.635 3588.000 2798.555 ;
        RECT 3379.715 2795.795 3588.000 2796.635 ;
        RECT 3379.435 2793.415 3588.000 2795.795 ;
        RECT 3379.715 2792.575 3588.000 2793.415 ;
        RECT 3379.435 2790.195 3588.000 2792.575 ;
        RECT 3379.715 2789.355 3588.000 2790.195 ;
        RECT 3379.435 2787.435 3588.000 2789.355 ;
      LAYER met2 ;
        RECT 3377.035 2786.875 3379.435 2787.155 ;
      LAYER met2 ;
        RECT 3379.715 2786.595 3588.000 2787.435 ;
        RECT 3379.435 2784.215 3588.000 2786.595 ;
        RECT 3379.715 2783.375 3588.000 2784.215 ;
        RECT 3379.435 2780.995 3588.000 2783.375 ;
      LAYER met2 ;
        RECT 3374.290 2780.745 3374.570 2780.840 ;
        RECT 3374.255 2780.405 3374.570 2780.745 ;
        RECT 3377.035 2780.435 3379.435 2780.715 ;
        RECT 3370.830 2749.585 3371.130 2749.925 ;
        RECT 3370.330 1916.025 3370.640 1916.365 ;
        RECT 3369.805 1900.845 3370.105 1901.185 ;
        RECT 214.955 1803.825 215.235 1804.165 ;
        RECT 214.430 1788.635 214.710 1788.975 ;
        RECT 213.920 1625.085 214.210 1625.425 ;
      LAYER met2 ;
        RECT 0.000 1591.625 208.565 1594.005 ;
        RECT 0.000 1590.785 208.285 1591.625 ;
        RECT 0.000 1588.405 208.565 1590.785 ;
        RECT 0.000 1587.565 208.285 1588.405 ;
      LAYER met2 ;
        RECT 210.370 1588.135 210.650 1588.165 ;
        RECT 210.145 1588.125 210.965 1588.135 ;
        RECT 208.565 1587.845 210.965 1588.125 ;
        RECT 210.370 1587.825 210.650 1587.845 ;
      LAYER met2 ;
        RECT 0.000 1585.645 208.565 1587.565 ;
        RECT 0.000 1584.805 208.285 1585.645 ;
        RECT 0.000 1582.425 208.565 1584.805 ;
        RECT 0.000 1581.585 208.285 1582.425 ;
        RECT 0.000 1579.205 208.565 1581.585 ;
        RECT 0.000 1578.365 208.285 1579.205 ;
        RECT 0.000 1576.445 208.565 1578.365 ;
        RECT 0.000 1575.605 208.285 1576.445 ;
        RECT 0.000 1573.225 208.565 1575.605 ;
        RECT 0.000 1572.385 208.285 1573.225 ;
      LAYER met2 ;
        RECT 210.370 1572.945 210.650 1572.975 ;
        RECT 208.565 1572.665 210.965 1572.945 ;
        RECT 210.370 1572.635 210.650 1572.665 ;
      LAYER met2 ;
        RECT 0.000 1570.005 208.565 1572.385 ;
        RECT 0.000 1569.165 208.285 1570.005 ;
        RECT 0.000 1567.245 208.565 1569.165 ;
        RECT 0.000 1566.405 208.285 1567.245 ;
        RECT 0.000 1564.025 208.565 1566.405 ;
        RECT 0.000 1563.185 208.285 1564.025 ;
        RECT 0.000 1560.805 208.565 1563.185 ;
        RECT 0.000 1559.965 208.285 1560.805 ;
        RECT 0.000 1558.045 208.565 1559.965 ;
        RECT 0.000 1557.205 208.285 1558.045 ;
        RECT 0.000 1556.210 208.565 1557.205 ;
        RECT 0.000 1418.865 208.565 1419.915 ;
        RECT 0.000 1418.025 208.285 1418.865 ;
      LAYER met2 ;
        RECT 212.370 1418.645 212.650 1418.720 ;
        RECT 210.370 1418.625 210.650 1418.645 ;
        RECT 209.945 1418.605 210.965 1418.625 ;
        RECT 209.910 1418.585 210.965 1418.605 ;
        RECT 208.565 1418.305 210.965 1418.585 ;
        RECT 212.370 1418.305 212.665 1418.645 ;
      LAYER met2 ;
        RECT 0.000 1415.645 208.565 1418.025 ;
        RECT 0.000 1414.805 208.285 1415.645 ;
        RECT 0.000 1412.425 208.565 1414.805 ;
        RECT 0.000 1411.585 208.285 1412.425 ;
      LAYER met2 ;
        RECT 208.565 1411.865 210.965 1412.145 ;
      LAYER met2 ;
        RECT 0.000 1409.665 208.565 1411.585 ;
        RECT 0.000 1408.825 208.285 1409.665 ;
      LAYER met2 ;
        RECT 210.370 1409.405 210.650 1409.425 ;
        RECT 209.945 1409.385 210.965 1409.405 ;
        RECT 208.565 1409.105 210.965 1409.385 ;
        RECT 210.370 1409.085 210.650 1409.105 ;
      LAYER met2 ;
        RECT 0.000 1406.445 208.565 1408.825 ;
        RECT 0.000 1405.605 208.285 1406.445 ;
        RECT 0.000 1403.225 208.565 1405.605 ;
        RECT 0.000 1402.385 208.285 1403.225 ;
        RECT 0.000 1400.465 208.565 1402.385 ;
        RECT 0.000 1399.625 208.285 1400.465 ;
      LAYER met2 ;
        RECT 208.565 1399.905 210.965 1400.185 ;
      LAYER met2 ;
        RECT 0.000 1397.245 208.565 1399.625 ;
        RECT 0.000 1396.405 208.285 1397.245 ;
        RECT 0.000 1394.025 208.565 1396.405 ;
        RECT 0.000 1393.185 208.285 1394.025 ;
        RECT 0.000 1391.265 208.565 1393.185 ;
        RECT 0.000 1390.425 208.285 1391.265 ;
        RECT 0.000 1388.045 208.565 1390.425 ;
        RECT 0.000 1387.205 208.285 1388.045 ;
        RECT 0.000 1384.825 208.565 1387.205 ;
        RECT 0.000 1383.985 208.285 1384.825 ;
        RECT 0.000 1382.065 208.565 1383.985 ;
        RECT 0.000 1381.225 208.285 1382.065 ;
        RECT 0.000 1378.845 208.565 1381.225 ;
        RECT 0.000 1378.005 208.285 1378.845 ;
      LAYER met2 ;
        RECT 210.370 1378.565 210.650 1378.585 ;
        RECT 208.565 1378.285 210.965 1378.565 ;
        RECT 209.400 1378.265 210.965 1378.285 ;
        RECT 210.370 1378.245 210.650 1378.265 ;
        RECT 212.370 1378.245 212.650 1418.305 ;
        RECT 213.960 1409.425 214.210 1625.085 ;
        RECT 214.460 1572.975 214.710 1788.635 ;
        RECT 214.960 1588.165 215.210 1803.825 ;
        RECT 3369.830 1675.185 3370.080 1900.845 ;
        RECT 3370.330 1690.365 3370.580 1916.025 ;
        RECT 3370.830 1863.925 3371.080 2749.585 ;
        RECT 3374.290 2740.385 3374.570 2780.405 ;
      LAYER met2 ;
        RECT 3379.715 2780.155 3588.000 2780.995 ;
        RECT 3379.435 2777.775 3588.000 2780.155 ;
        RECT 3379.715 2776.935 3588.000 2777.775 ;
        RECT 3379.435 2775.015 3588.000 2776.935 ;
        RECT 3379.715 2774.175 3588.000 2775.015 ;
        RECT 3379.435 2771.795 3588.000 2774.175 ;
        RECT 3379.715 2770.955 3588.000 2771.795 ;
        RECT 3379.435 2768.575 3588.000 2770.955 ;
        RECT 3379.715 2767.735 3588.000 2768.575 ;
        RECT 3379.435 2765.815 3588.000 2767.735 ;
        RECT 3379.715 2764.975 3588.000 2765.815 ;
        RECT 3379.435 2762.595 3588.000 2764.975 ;
        RECT 3379.715 2761.755 3588.000 2762.595 ;
        RECT 3379.435 2759.375 3588.000 2761.755 ;
      LAYER met2 ;
        RECT 3377.035 2758.815 3379.435 2759.095 ;
      LAYER met2 ;
        RECT 3379.715 2758.535 3588.000 2759.375 ;
        RECT 3379.435 2756.615 3588.000 2758.535 ;
        RECT 3379.715 2755.775 3588.000 2756.615 ;
        RECT 3379.435 2753.395 3588.000 2755.775 ;
        RECT 3379.715 2752.555 3588.000 2753.395 ;
        RECT 3379.435 2750.175 3588.000 2752.555 ;
      LAYER met2 ;
        RECT 3377.035 2749.615 3379.435 2749.895 ;
      LAYER met2 ;
        RECT 3379.715 2749.335 3588.000 2750.175 ;
        RECT 3379.435 2747.415 3588.000 2749.335 ;
      LAYER met2 ;
        RECT 3377.035 2746.855 3379.435 2747.135 ;
      LAYER met2 ;
        RECT 3379.715 2746.575 3588.000 2747.415 ;
        RECT 3379.435 2744.195 3588.000 2746.575 ;
        RECT 3379.715 2743.355 3588.000 2744.195 ;
        RECT 3379.435 2740.975 3588.000 2743.355 ;
      LAYER met2 ;
        RECT 3377.525 2740.695 3377.785 2740.705 ;
        RECT 3377.035 2740.415 3379.435 2740.695 ;
        RECT 3377.525 2740.385 3377.785 2740.415 ;
      LAYER met2 ;
        RECT 3379.715 2740.135 3588.000 2740.975 ;
        RECT 3379.435 2739.085 3588.000 2740.135 ;
        RECT 3390.035 2593.505 3583.075 2593.735 ;
        RECT 3388.000 2569.605 3583.075 2593.505 ;
        RECT 3388.000 2566.105 3389.920 2568.105 ;
        RECT 3390.035 2543.610 3583.075 2569.605 ;
        RECT 3388.000 2519.710 3583.075 2543.610 ;
        RECT 3390.035 2152.505 3583.075 2152.735 ;
        RECT 3388.000 2128.605 3583.075 2152.505 ;
        RECT 3388.000 2125.105 3389.920 2127.105 ;
        RECT 3390.035 2102.610 3583.075 2128.605 ;
        RECT 3388.000 2078.710 3583.075 2102.610 ;
        RECT 3379.435 1931.795 3588.000 1932.790 ;
        RECT 3379.715 1930.955 3588.000 1931.795 ;
        RECT 3379.435 1929.035 3588.000 1930.955 ;
        RECT 3379.715 1928.195 3588.000 1929.035 ;
        RECT 3379.435 1925.815 3588.000 1928.195 ;
        RECT 3379.715 1924.975 3588.000 1925.815 ;
        RECT 3379.435 1922.595 3588.000 1924.975 ;
        RECT 3379.715 1921.755 3588.000 1922.595 ;
        RECT 3379.435 1919.835 3588.000 1921.755 ;
        RECT 3379.715 1918.995 3588.000 1919.835 ;
        RECT 3379.435 1916.615 3588.000 1918.995 ;
      LAYER met2 ;
        RECT 3377.035 1916.055 3379.435 1916.335 ;
      LAYER met2 ;
        RECT 3379.715 1915.775 3588.000 1916.615 ;
        RECT 3379.435 1913.395 3588.000 1915.775 ;
        RECT 3379.715 1912.555 3588.000 1913.395 ;
        RECT 3379.435 1910.635 3588.000 1912.555 ;
        RECT 3379.715 1909.795 3588.000 1910.635 ;
        RECT 3379.435 1907.415 3588.000 1909.795 ;
        RECT 3379.715 1906.575 3588.000 1907.415 ;
        RECT 3379.435 1904.195 3588.000 1906.575 ;
        RECT 3379.715 1903.355 3588.000 1904.195 ;
        RECT 3379.435 1901.435 3588.000 1903.355 ;
      LAYER met2 ;
        RECT 3377.035 1900.875 3379.435 1901.155 ;
      LAYER met2 ;
        RECT 3379.715 1900.595 3588.000 1901.435 ;
        RECT 3379.435 1898.215 3588.000 1900.595 ;
        RECT 3379.715 1897.375 3588.000 1898.215 ;
        RECT 3379.435 1894.995 3588.000 1897.375 ;
      LAYER met2 ;
        RECT 3374.290 1894.745 3374.570 1894.840 ;
        RECT 3374.255 1894.405 3374.570 1894.745 ;
        RECT 3377.035 1894.435 3379.435 1894.715 ;
        RECT 3370.830 1863.585 3371.130 1863.925 ;
        RECT 3370.330 1690.025 3370.640 1690.365 ;
        RECT 3369.805 1674.845 3370.105 1675.185 ;
        RECT 214.955 1587.825 215.235 1588.165 ;
        RECT 214.430 1572.635 214.710 1572.975 ;
        RECT 213.920 1409.085 214.210 1409.425 ;
      LAYER met2 ;
        RECT 0.000 1375.625 208.565 1378.005 ;
        RECT 0.000 1374.785 208.285 1375.625 ;
        RECT 0.000 1372.405 208.565 1374.785 ;
        RECT 0.000 1371.565 208.285 1372.405 ;
      LAYER met2 ;
        RECT 210.370 1372.135 210.650 1372.165 ;
        RECT 210.145 1372.125 210.965 1372.135 ;
        RECT 208.565 1371.845 210.965 1372.125 ;
        RECT 210.370 1371.825 210.650 1371.845 ;
      LAYER met2 ;
        RECT 0.000 1369.645 208.565 1371.565 ;
        RECT 0.000 1368.805 208.285 1369.645 ;
        RECT 0.000 1366.425 208.565 1368.805 ;
        RECT 0.000 1365.585 208.285 1366.425 ;
        RECT 0.000 1363.205 208.565 1365.585 ;
        RECT 0.000 1362.365 208.285 1363.205 ;
        RECT 0.000 1360.445 208.565 1362.365 ;
        RECT 0.000 1359.605 208.285 1360.445 ;
        RECT 0.000 1357.225 208.565 1359.605 ;
        RECT 0.000 1356.385 208.285 1357.225 ;
      LAYER met2 ;
        RECT 210.370 1356.945 210.650 1356.975 ;
        RECT 208.565 1356.665 210.965 1356.945 ;
        RECT 210.370 1356.635 210.650 1356.665 ;
      LAYER met2 ;
        RECT 0.000 1354.005 208.565 1356.385 ;
        RECT 0.000 1353.165 208.285 1354.005 ;
        RECT 0.000 1351.245 208.565 1353.165 ;
        RECT 0.000 1350.405 208.285 1351.245 ;
        RECT 0.000 1348.025 208.565 1350.405 ;
        RECT 0.000 1347.185 208.285 1348.025 ;
        RECT 0.000 1344.805 208.565 1347.185 ;
        RECT 0.000 1343.965 208.285 1344.805 ;
        RECT 0.000 1342.045 208.565 1343.965 ;
        RECT 0.000 1341.205 208.285 1342.045 ;
        RECT 0.000 1340.210 208.565 1341.205 ;
        RECT 0.000 1202.865 208.565 1203.915 ;
        RECT 0.000 1202.025 208.285 1202.865 ;
      LAYER met2 ;
        RECT 212.370 1202.645 212.650 1202.720 ;
        RECT 210.370 1202.625 210.650 1202.645 ;
        RECT 209.945 1202.605 210.965 1202.625 ;
        RECT 209.910 1202.585 210.965 1202.605 ;
        RECT 208.565 1202.305 210.965 1202.585 ;
        RECT 212.370 1202.305 212.665 1202.645 ;
      LAYER met2 ;
        RECT 0.000 1199.645 208.565 1202.025 ;
        RECT 0.000 1198.805 208.285 1199.645 ;
        RECT 0.000 1196.425 208.565 1198.805 ;
        RECT 0.000 1195.585 208.285 1196.425 ;
      LAYER met2 ;
        RECT 208.565 1195.865 210.965 1196.145 ;
      LAYER met2 ;
        RECT 0.000 1193.665 208.565 1195.585 ;
        RECT 0.000 1192.825 208.285 1193.665 ;
      LAYER met2 ;
        RECT 210.370 1193.405 210.650 1193.425 ;
        RECT 209.945 1193.385 210.965 1193.405 ;
        RECT 208.565 1193.105 210.965 1193.385 ;
        RECT 210.370 1193.085 210.650 1193.105 ;
      LAYER met2 ;
        RECT 0.000 1190.445 208.565 1192.825 ;
        RECT 0.000 1189.605 208.285 1190.445 ;
        RECT 0.000 1187.225 208.565 1189.605 ;
        RECT 0.000 1186.385 208.285 1187.225 ;
      LAYER met2 ;
        RECT 208.565 1186.665 210.965 1186.945 ;
      LAYER met2 ;
        RECT 0.000 1184.465 208.565 1186.385 ;
        RECT 0.000 1183.625 208.285 1184.465 ;
      LAYER met2 ;
        RECT 208.565 1183.905 210.965 1184.185 ;
      LAYER met2 ;
        RECT 0.000 1181.245 208.565 1183.625 ;
        RECT 0.000 1180.405 208.285 1181.245 ;
        RECT 0.000 1178.025 208.565 1180.405 ;
        RECT 0.000 1177.185 208.285 1178.025 ;
      LAYER met2 ;
        RECT 208.565 1177.465 210.965 1177.745 ;
      LAYER met2 ;
        RECT 0.000 1175.265 208.565 1177.185 ;
        RECT 0.000 1174.425 208.285 1175.265 ;
        RECT 0.000 1172.045 208.565 1174.425 ;
        RECT 0.000 1171.205 208.285 1172.045 ;
        RECT 0.000 1168.825 208.565 1171.205 ;
        RECT 0.000 1167.985 208.285 1168.825 ;
        RECT 0.000 1166.065 208.565 1167.985 ;
        RECT 0.000 1165.225 208.285 1166.065 ;
        RECT 0.000 1162.845 208.565 1165.225 ;
        RECT 0.000 1162.005 208.285 1162.845 ;
      LAYER met2 ;
        RECT 210.370 1162.565 210.650 1162.585 ;
        RECT 208.565 1162.285 210.965 1162.565 ;
        RECT 209.400 1162.265 210.965 1162.285 ;
        RECT 210.370 1162.245 210.650 1162.265 ;
        RECT 212.370 1162.245 212.650 1202.305 ;
        RECT 213.960 1193.425 214.210 1409.085 ;
        RECT 214.460 1356.975 214.710 1572.635 ;
        RECT 214.960 1372.165 215.210 1587.825 ;
        RECT 3369.830 1450.185 3370.080 1674.845 ;
        RECT 3370.330 1465.365 3370.580 1690.025 ;
        RECT 3370.830 1637.925 3371.080 1863.585 ;
        RECT 3374.290 1854.385 3374.570 1894.405 ;
      LAYER met2 ;
        RECT 3379.715 1894.155 3588.000 1894.995 ;
        RECT 3379.435 1891.775 3588.000 1894.155 ;
        RECT 3379.715 1890.935 3588.000 1891.775 ;
        RECT 3379.435 1889.015 3588.000 1890.935 ;
        RECT 3379.715 1888.175 3588.000 1889.015 ;
        RECT 3379.435 1885.795 3588.000 1888.175 ;
        RECT 3379.715 1884.955 3588.000 1885.795 ;
        RECT 3379.435 1882.575 3588.000 1884.955 ;
        RECT 3379.715 1881.735 3588.000 1882.575 ;
        RECT 3379.435 1879.815 3588.000 1881.735 ;
      LAYER met2 ;
        RECT 3377.035 1879.255 3379.435 1879.535 ;
      LAYER met2 ;
        RECT 3379.715 1878.975 3588.000 1879.815 ;
        RECT 3379.435 1876.595 3588.000 1878.975 ;
        RECT 3379.715 1875.755 3588.000 1876.595 ;
        RECT 3379.435 1873.375 3588.000 1875.755 ;
      LAYER met2 ;
        RECT 3377.035 1872.815 3379.435 1873.095 ;
      LAYER met2 ;
        RECT 3379.715 1872.535 3588.000 1873.375 ;
        RECT 3379.435 1870.615 3588.000 1872.535 ;
      LAYER met2 ;
        RECT 3377.035 1870.055 3379.435 1870.335 ;
      LAYER met2 ;
        RECT 3379.715 1869.775 3588.000 1870.615 ;
        RECT 3379.435 1867.395 3588.000 1869.775 ;
        RECT 3379.715 1866.555 3588.000 1867.395 ;
        RECT 3379.435 1864.175 3588.000 1866.555 ;
      LAYER met2 ;
        RECT 3377.035 1863.615 3379.435 1863.895 ;
      LAYER met2 ;
        RECT 3379.715 1863.335 3588.000 1864.175 ;
        RECT 3379.435 1861.415 3588.000 1863.335 ;
      LAYER met2 ;
        RECT 3377.035 1860.855 3379.435 1861.135 ;
      LAYER met2 ;
        RECT 3379.715 1860.575 3588.000 1861.415 ;
        RECT 3379.435 1858.195 3588.000 1860.575 ;
        RECT 3379.715 1857.355 3588.000 1858.195 ;
        RECT 3379.435 1854.975 3588.000 1857.355 ;
      LAYER met2 ;
        RECT 3377.525 1854.695 3377.785 1854.705 ;
        RECT 3377.035 1854.415 3379.435 1854.695 ;
        RECT 3377.525 1854.385 3377.785 1854.415 ;
      LAYER met2 ;
        RECT 3379.715 1854.135 3588.000 1854.975 ;
        RECT 3379.435 1853.085 3588.000 1854.135 ;
        RECT 3379.435 1705.795 3588.000 1706.790 ;
        RECT 3379.715 1704.955 3588.000 1705.795 ;
        RECT 3379.435 1703.035 3588.000 1704.955 ;
        RECT 3379.715 1702.195 3588.000 1703.035 ;
        RECT 3379.435 1699.815 3588.000 1702.195 ;
        RECT 3379.715 1698.975 3588.000 1699.815 ;
        RECT 3379.435 1696.595 3588.000 1698.975 ;
        RECT 3379.715 1695.755 3588.000 1696.595 ;
        RECT 3379.435 1693.835 3588.000 1695.755 ;
        RECT 3379.715 1692.995 3588.000 1693.835 ;
        RECT 3379.435 1690.615 3588.000 1692.995 ;
      LAYER met2 ;
        RECT 3377.035 1690.055 3379.435 1690.335 ;
      LAYER met2 ;
        RECT 3379.715 1689.775 3588.000 1690.615 ;
        RECT 3379.435 1687.395 3588.000 1689.775 ;
        RECT 3379.715 1686.555 3588.000 1687.395 ;
        RECT 3379.435 1684.635 3588.000 1686.555 ;
        RECT 3379.715 1683.795 3588.000 1684.635 ;
        RECT 3379.435 1681.415 3588.000 1683.795 ;
        RECT 3379.715 1680.575 3588.000 1681.415 ;
        RECT 3379.435 1678.195 3588.000 1680.575 ;
        RECT 3379.715 1677.355 3588.000 1678.195 ;
        RECT 3379.435 1675.435 3588.000 1677.355 ;
      LAYER met2 ;
        RECT 3377.035 1674.875 3379.435 1675.155 ;
      LAYER met2 ;
        RECT 3379.715 1674.595 3588.000 1675.435 ;
        RECT 3379.435 1672.215 3588.000 1674.595 ;
        RECT 3379.715 1671.375 3588.000 1672.215 ;
        RECT 3379.435 1668.995 3588.000 1671.375 ;
      LAYER met2 ;
        RECT 3373.290 1668.745 3373.570 1668.840 ;
        RECT 3373.255 1668.405 3373.570 1668.745 ;
        RECT 3377.035 1668.435 3379.435 1668.715 ;
        RECT 3370.830 1637.585 3371.130 1637.925 ;
        RECT 3370.330 1465.025 3370.640 1465.365 ;
        RECT 3369.805 1449.845 3370.105 1450.185 ;
        RECT 214.955 1371.825 215.235 1372.165 ;
        RECT 214.430 1356.635 214.710 1356.975 ;
        RECT 213.920 1193.085 214.210 1193.425 ;
      LAYER met2 ;
        RECT 0.000 1159.625 208.565 1162.005 ;
        RECT 0.000 1158.785 208.285 1159.625 ;
        RECT 0.000 1156.405 208.565 1158.785 ;
        RECT 0.000 1155.565 208.285 1156.405 ;
      LAYER met2 ;
        RECT 210.370 1156.135 210.650 1156.165 ;
        RECT 210.145 1156.125 210.965 1156.135 ;
        RECT 208.565 1155.845 210.965 1156.125 ;
        RECT 210.370 1155.825 210.650 1155.845 ;
      LAYER met2 ;
        RECT 0.000 1153.645 208.565 1155.565 ;
        RECT 0.000 1152.805 208.285 1153.645 ;
        RECT 0.000 1150.425 208.565 1152.805 ;
        RECT 0.000 1149.585 208.285 1150.425 ;
        RECT 0.000 1147.205 208.565 1149.585 ;
        RECT 0.000 1146.365 208.285 1147.205 ;
        RECT 0.000 1144.445 208.565 1146.365 ;
        RECT 0.000 1143.605 208.285 1144.445 ;
        RECT 0.000 1141.225 208.565 1143.605 ;
        RECT 0.000 1140.385 208.285 1141.225 ;
      LAYER met2 ;
        RECT 210.370 1140.945 210.650 1140.975 ;
        RECT 208.565 1140.665 210.965 1140.945 ;
        RECT 210.370 1140.635 210.650 1140.665 ;
      LAYER met2 ;
        RECT 0.000 1138.005 208.565 1140.385 ;
        RECT 0.000 1137.165 208.285 1138.005 ;
        RECT 0.000 1135.245 208.565 1137.165 ;
        RECT 0.000 1134.405 208.285 1135.245 ;
        RECT 0.000 1132.025 208.565 1134.405 ;
        RECT 0.000 1131.185 208.285 1132.025 ;
        RECT 0.000 1128.805 208.565 1131.185 ;
        RECT 0.000 1127.965 208.285 1128.805 ;
        RECT 0.000 1126.045 208.565 1127.965 ;
        RECT 0.000 1125.205 208.285 1126.045 ;
        RECT 0.000 1124.210 208.565 1125.205 ;
        RECT 0.000 986.865 208.565 987.915 ;
        RECT 0.000 986.025 208.285 986.865 ;
      LAYER met2 ;
        RECT 212.370 986.645 212.650 986.720 ;
        RECT 210.370 986.625 210.650 986.645 ;
        RECT 209.945 986.605 210.965 986.625 ;
        RECT 209.910 986.585 210.965 986.605 ;
        RECT 208.565 986.305 210.965 986.585 ;
        RECT 212.370 986.305 212.665 986.645 ;
      LAYER met2 ;
        RECT 0.000 983.645 208.565 986.025 ;
        RECT 0.000 982.805 208.285 983.645 ;
        RECT 0.000 980.425 208.565 982.805 ;
        RECT 0.000 979.585 208.285 980.425 ;
      LAYER met2 ;
        RECT 208.565 979.865 210.965 980.145 ;
      LAYER met2 ;
        RECT 0.000 977.665 208.565 979.585 ;
        RECT 0.000 976.825 208.285 977.665 ;
      LAYER met2 ;
        RECT 210.370 977.405 210.650 977.425 ;
        RECT 209.945 977.385 210.965 977.405 ;
        RECT 208.565 977.105 210.965 977.385 ;
        RECT 210.370 977.085 210.650 977.105 ;
      LAYER met2 ;
        RECT 0.000 974.445 208.565 976.825 ;
        RECT 0.000 973.605 208.285 974.445 ;
        RECT 0.000 971.225 208.565 973.605 ;
        RECT 0.000 970.385 208.285 971.225 ;
      LAYER met2 ;
        RECT 208.565 970.665 210.965 970.945 ;
      LAYER met2 ;
        RECT 0.000 968.465 208.565 970.385 ;
        RECT 0.000 967.625 208.285 968.465 ;
      LAYER met2 ;
        RECT 208.565 967.905 210.965 968.185 ;
      LAYER met2 ;
        RECT 0.000 965.245 208.565 967.625 ;
        RECT 0.000 964.405 208.285 965.245 ;
        RECT 0.000 962.025 208.565 964.405 ;
        RECT 0.000 961.185 208.285 962.025 ;
      LAYER met2 ;
        RECT 208.565 961.465 210.965 961.745 ;
      LAYER met2 ;
        RECT 0.000 959.265 208.565 961.185 ;
        RECT 0.000 958.425 208.285 959.265 ;
        RECT 0.000 956.045 208.565 958.425 ;
        RECT 0.000 955.205 208.285 956.045 ;
        RECT 0.000 952.825 208.565 955.205 ;
        RECT 0.000 951.985 208.285 952.825 ;
        RECT 0.000 950.065 208.565 951.985 ;
        RECT 0.000 949.225 208.285 950.065 ;
        RECT 0.000 946.845 208.565 949.225 ;
        RECT 0.000 946.005 208.285 946.845 ;
      LAYER met2 ;
        RECT 210.370 946.565 210.650 946.585 ;
        RECT 208.565 946.285 210.965 946.565 ;
        RECT 209.400 946.265 210.965 946.285 ;
        RECT 210.370 946.245 210.650 946.265 ;
        RECT 212.370 946.245 212.650 986.305 ;
        RECT 213.960 977.425 214.210 1193.085 ;
        RECT 214.460 1140.975 214.710 1356.635 ;
        RECT 214.960 1156.165 215.210 1371.825 ;
        RECT 3369.830 1225.185 3370.080 1449.845 ;
        RECT 3370.330 1240.365 3370.580 1465.025 ;
        RECT 3370.830 1412.925 3371.080 1637.585 ;
        RECT 3373.290 1628.385 3373.570 1668.405 ;
      LAYER met2 ;
        RECT 3379.715 1668.155 3588.000 1668.995 ;
        RECT 3379.435 1665.775 3588.000 1668.155 ;
        RECT 3379.715 1664.935 3588.000 1665.775 ;
        RECT 3379.435 1663.015 3588.000 1664.935 ;
        RECT 3379.715 1662.175 3588.000 1663.015 ;
        RECT 3379.435 1659.795 3588.000 1662.175 ;
        RECT 3379.715 1658.955 3588.000 1659.795 ;
        RECT 3379.435 1656.575 3588.000 1658.955 ;
        RECT 3379.715 1655.735 3588.000 1656.575 ;
        RECT 3379.435 1653.815 3588.000 1655.735 ;
      LAYER met2 ;
        RECT 3377.035 1653.255 3379.435 1653.535 ;
      LAYER met2 ;
        RECT 3379.715 1652.975 3588.000 1653.815 ;
        RECT 3379.435 1650.595 3588.000 1652.975 ;
        RECT 3379.715 1649.755 3588.000 1650.595 ;
        RECT 3379.435 1647.375 3588.000 1649.755 ;
      LAYER met2 ;
        RECT 3377.035 1646.815 3379.435 1647.095 ;
      LAYER met2 ;
        RECT 3379.715 1646.535 3588.000 1647.375 ;
        RECT 3379.435 1644.615 3588.000 1646.535 ;
      LAYER met2 ;
        RECT 3377.035 1644.055 3379.435 1644.335 ;
      LAYER met2 ;
        RECT 3379.715 1643.775 3588.000 1644.615 ;
        RECT 3379.435 1641.395 3588.000 1643.775 ;
        RECT 3379.715 1640.555 3588.000 1641.395 ;
        RECT 3379.435 1638.175 3588.000 1640.555 ;
      LAYER met2 ;
        RECT 3377.035 1637.615 3379.435 1637.895 ;
      LAYER met2 ;
        RECT 3379.715 1637.335 3588.000 1638.175 ;
        RECT 3379.435 1635.415 3588.000 1637.335 ;
      LAYER met2 ;
        RECT 3377.035 1634.855 3379.435 1635.135 ;
      LAYER met2 ;
        RECT 3379.715 1634.575 3588.000 1635.415 ;
        RECT 3379.435 1632.195 3588.000 1634.575 ;
        RECT 3379.715 1631.355 3588.000 1632.195 ;
        RECT 3379.435 1628.975 3588.000 1631.355 ;
      LAYER met2 ;
        RECT 3377.525 1628.695 3377.785 1628.705 ;
        RECT 3377.035 1628.415 3379.435 1628.695 ;
        RECT 3377.525 1628.385 3377.785 1628.415 ;
      LAYER met2 ;
        RECT 3379.715 1628.135 3588.000 1628.975 ;
        RECT 3379.435 1627.085 3588.000 1628.135 ;
        RECT 3379.435 1480.795 3588.000 1481.790 ;
        RECT 3379.715 1479.955 3588.000 1480.795 ;
        RECT 3379.435 1478.035 3588.000 1479.955 ;
        RECT 3379.715 1477.195 3588.000 1478.035 ;
        RECT 3379.435 1474.815 3588.000 1477.195 ;
        RECT 3379.715 1473.975 3588.000 1474.815 ;
        RECT 3379.435 1471.595 3588.000 1473.975 ;
        RECT 3379.715 1470.755 3588.000 1471.595 ;
        RECT 3379.435 1468.835 3588.000 1470.755 ;
        RECT 3379.715 1467.995 3588.000 1468.835 ;
        RECT 3379.435 1465.615 3588.000 1467.995 ;
      LAYER met2 ;
        RECT 3377.035 1465.055 3379.435 1465.335 ;
      LAYER met2 ;
        RECT 3379.715 1464.775 3588.000 1465.615 ;
        RECT 3379.435 1462.395 3588.000 1464.775 ;
        RECT 3379.715 1461.555 3588.000 1462.395 ;
        RECT 3379.435 1459.635 3588.000 1461.555 ;
        RECT 3379.715 1458.795 3588.000 1459.635 ;
        RECT 3379.435 1456.415 3588.000 1458.795 ;
        RECT 3379.715 1455.575 3588.000 1456.415 ;
        RECT 3379.435 1453.195 3588.000 1455.575 ;
        RECT 3379.715 1452.355 3588.000 1453.195 ;
        RECT 3379.435 1450.435 3588.000 1452.355 ;
      LAYER met2 ;
        RECT 3377.035 1449.875 3379.435 1450.155 ;
      LAYER met2 ;
        RECT 3379.715 1449.595 3588.000 1450.435 ;
        RECT 3379.435 1447.215 3588.000 1449.595 ;
        RECT 3379.715 1446.375 3588.000 1447.215 ;
        RECT 3379.435 1443.995 3588.000 1446.375 ;
      LAYER met2 ;
        RECT 3373.290 1443.745 3373.570 1443.840 ;
        RECT 3373.255 1443.405 3373.570 1443.745 ;
        RECT 3377.035 1443.435 3379.435 1443.715 ;
        RECT 3370.830 1412.585 3371.130 1412.925 ;
        RECT 3370.330 1240.025 3370.640 1240.365 ;
        RECT 3369.805 1224.845 3370.105 1225.185 ;
        RECT 214.955 1155.825 215.235 1156.165 ;
        RECT 214.430 1140.635 214.710 1140.975 ;
        RECT 213.920 977.085 214.210 977.425 ;
      LAYER met2 ;
        RECT 0.000 943.625 208.565 946.005 ;
        RECT 0.000 942.785 208.285 943.625 ;
        RECT 0.000 940.405 208.565 942.785 ;
        RECT 0.000 939.565 208.285 940.405 ;
      LAYER met2 ;
        RECT 210.370 940.135 210.650 940.165 ;
        RECT 209.935 940.125 210.965 940.135 ;
        RECT 208.565 939.845 210.965 940.125 ;
        RECT 210.370 939.825 210.650 939.845 ;
      LAYER met2 ;
        RECT 0.000 937.645 208.565 939.565 ;
        RECT 0.000 936.805 208.285 937.645 ;
        RECT 0.000 934.425 208.565 936.805 ;
        RECT 0.000 933.585 208.285 934.425 ;
        RECT 0.000 931.205 208.565 933.585 ;
        RECT 0.000 930.365 208.285 931.205 ;
        RECT 0.000 928.445 208.565 930.365 ;
        RECT 0.000 927.605 208.285 928.445 ;
        RECT 0.000 925.225 208.565 927.605 ;
        RECT 0.000 924.385 208.285 925.225 ;
      LAYER met2 ;
        RECT 210.370 924.945 210.650 924.975 ;
        RECT 208.565 924.665 210.965 924.945 ;
        RECT 210.370 924.635 210.650 924.665 ;
      LAYER met2 ;
        RECT 0.000 922.005 208.565 924.385 ;
        RECT 0.000 921.165 208.285 922.005 ;
        RECT 0.000 919.245 208.565 921.165 ;
        RECT 0.000 918.405 208.285 919.245 ;
        RECT 0.000 916.025 208.565 918.405 ;
        RECT 0.000 915.185 208.285 916.025 ;
        RECT 0.000 912.805 208.565 915.185 ;
        RECT 0.000 911.965 208.285 912.805 ;
        RECT 0.000 910.045 208.565 911.965 ;
        RECT 0.000 909.205 208.285 910.045 ;
        RECT 0.000 908.210 208.565 909.205 ;
      LAYER met2 ;
        RECT 213.960 905.430 214.210 977.085 ;
        RECT 214.460 924.975 214.710 1140.635 ;
        RECT 214.960 940.165 215.210 1155.825 ;
        RECT 3369.830 999.185 3370.080 1224.845 ;
        RECT 3370.330 1014.365 3370.580 1240.025 ;
        RECT 3370.830 1187.925 3371.080 1412.585 ;
        RECT 3373.290 1403.385 3373.570 1443.405 ;
      LAYER met2 ;
        RECT 3379.715 1443.155 3588.000 1443.995 ;
        RECT 3379.435 1440.775 3588.000 1443.155 ;
        RECT 3379.715 1439.935 3588.000 1440.775 ;
        RECT 3379.435 1438.015 3588.000 1439.935 ;
        RECT 3379.715 1437.175 3588.000 1438.015 ;
        RECT 3379.435 1434.795 3588.000 1437.175 ;
        RECT 3379.715 1433.955 3588.000 1434.795 ;
        RECT 3379.435 1431.575 3588.000 1433.955 ;
        RECT 3379.715 1430.735 3588.000 1431.575 ;
        RECT 3379.435 1428.815 3588.000 1430.735 ;
      LAYER met2 ;
        RECT 3377.035 1428.255 3379.435 1428.535 ;
      LAYER met2 ;
        RECT 3379.715 1427.975 3588.000 1428.815 ;
        RECT 3379.435 1425.595 3588.000 1427.975 ;
        RECT 3379.715 1424.755 3588.000 1425.595 ;
        RECT 3379.435 1422.375 3588.000 1424.755 ;
      LAYER met2 ;
        RECT 3377.035 1421.815 3379.435 1422.095 ;
      LAYER met2 ;
        RECT 3379.715 1421.535 3588.000 1422.375 ;
        RECT 3379.435 1419.615 3588.000 1421.535 ;
      LAYER met2 ;
        RECT 3377.035 1419.055 3379.435 1419.335 ;
      LAYER met2 ;
        RECT 3379.715 1418.775 3588.000 1419.615 ;
        RECT 3379.435 1416.395 3588.000 1418.775 ;
        RECT 3379.715 1415.555 3588.000 1416.395 ;
        RECT 3379.435 1413.175 3588.000 1415.555 ;
      LAYER met2 ;
        RECT 3377.035 1412.615 3379.435 1412.895 ;
      LAYER met2 ;
        RECT 3379.715 1412.335 3588.000 1413.175 ;
        RECT 3379.435 1410.415 3588.000 1412.335 ;
      LAYER met2 ;
        RECT 3377.035 1409.855 3379.435 1410.135 ;
      LAYER met2 ;
        RECT 3379.715 1409.575 3588.000 1410.415 ;
        RECT 3379.435 1407.195 3588.000 1409.575 ;
        RECT 3379.715 1406.355 3588.000 1407.195 ;
        RECT 3379.435 1403.975 3588.000 1406.355 ;
      LAYER met2 ;
        RECT 3377.525 1403.695 3377.785 1403.705 ;
        RECT 3377.035 1403.415 3379.435 1403.695 ;
        RECT 3377.525 1403.385 3377.785 1403.415 ;
      LAYER met2 ;
        RECT 3379.715 1403.135 3588.000 1403.975 ;
        RECT 3379.435 1402.085 3588.000 1403.135 ;
        RECT 3379.435 1255.795 3588.000 1256.790 ;
        RECT 3379.715 1254.955 3588.000 1255.795 ;
        RECT 3379.435 1253.035 3588.000 1254.955 ;
        RECT 3379.715 1252.195 3588.000 1253.035 ;
        RECT 3379.435 1249.815 3588.000 1252.195 ;
        RECT 3379.715 1248.975 3588.000 1249.815 ;
        RECT 3379.435 1246.595 3588.000 1248.975 ;
        RECT 3379.715 1245.755 3588.000 1246.595 ;
        RECT 3379.435 1243.835 3588.000 1245.755 ;
        RECT 3379.715 1242.995 3588.000 1243.835 ;
        RECT 3379.435 1240.615 3588.000 1242.995 ;
      LAYER met2 ;
        RECT 3377.035 1240.055 3379.435 1240.335 ;
      LAYER met2 ;
        RECT 3379.715 1239.775 3588.000 1240.615 ;
        RECT 3379.435 1237.395 3588.000 1239.775 ;
        RECT 3379.715 1236.555 3588.000 1237.395 ;
        RECT 3379.435 1234.635 3588.000 1236.555 ;
        RECT 3379.715 1233.795 3588.000 1234.635 ;
        RECT 3379.435 1231.415 3588.000 1233.795 ;
        RECT 3379.715 1230.575 3588.000 1231.415 ;
        RECT 3379.435 1228.195 3588.000 1230.575 ;
        RECT 3379.715 1227.355 3588.000 1228.195 ;
        RECT 3379.435 1225.435 3588.000 1227.355 ;
      LAYER met2 ;
        RECT 3377.035 1224.875 3379.435 1225.155 ;
      LAYER met2 ;
        RECT 3379.715 1224.595 3588.000 1225.435 ;
        RECT 3379.435 1222.215 3588.000 1224.595 ;
        RECT 3379.715 1221.375 3588.000 1222.215 ;
        RECT 3379.435 1218.995 3588.000 1221.375 ;
      LAYER met2 ;
        RECT 3373.290 1218.745 3373.570 1218.840 ;
        RECT 3373.255 1218.405 3373.570 1218.745 ;
        RECT 3377.035 1218.435 3379.435 1218.715 ;
        RECT 3370.830 1187.585 3371.130 1187.925 ;
        RECT 3370.330 1014.025 3370.640 1014.365 ;
        RECT 3369.805 998.845 3370.105 999.185 ;
        RECT 214.955 939.825 215.235 940.165 ;
        RECT 214.430 924.635 214.710 924.975 ;
        RECT 213.950 905.110 214.210 905.430 ;
        RECT 213.960 905.090 214.210 905.110 ;
        RECT 214.460 904.930 214.710 924.635 ;
        RECT 214.460 904.610 214.720 904.930 ;
        RECT 214.460 904.535 214.710 904.610 ;
        RECT 214.960 904.430 215.210 939.825 ;
        RECT 214.950 904.110 215.210 904.430 ;
        RECT 214.960 904.040 215.210 904.110 ;
        RECT 3369.830 774.185 3370.080 998.845 ;
        RECT 3370.330 789.365 3370.580 1014.025 ;
        RECT 3370.830 961.925 3371.080 1187.585 ;
        RECT 3373.290 1178.385 3373.570 1218.405 ;
      LAYER met2 ;
        RECT 3379.715 1218.155 3588.000 1218.995 ;
        RECT 3379.435 1215.775 3588.000 1218.155 ;
        RECT 3379.715 1214.935 3588.000 1215.775 ;
        RECT 3379.435 1213.015 3588.000 1214.935 ;
        RECT 3379.715 1212.175 3588.000 1213.015 ;
        RECT 3379.435 1209.795 3588.000 1212.175 ;
        RECT 3379.715 1208.955 3588.000 1209.795 ;
        RECT 3379.435 1206.575 3588.000 1208.955 ;
        RECT 3379.715 1205.735 3588.000 1206.575 ;
        RECT 3379.435 1203.815 3588.000 1205.735 ;
      LAYER met2 ;
        RECT 3377.035 1203.255 3379.435 1203.535 ;
      LAYER met2 ;
        RECT 3379.715 1202.975 3588.000 1203.815 ;
        RECT 3379.435 1200.595 3588.000 1202.975 ;
        RECT 3379.715 1199.755 3588.000 1200.595 ;
        RECT 3379.435 1197.375 3588.000 1199.755 ;
      LAYER met2 ;
        RECT 3377.035 1196.815 3379.435 1197.095 ;
      LAYER met2 ;
        RECT 3379.715 1196.535 3588.000 1197.375 ;
        RECT 3379.435 1194.615 3588.000 1196.535 ;
      LAYER met2 ;
        RECT 3377.035 1194.055 3379.435 1194.335 ;
      LAYER met2 ;
        RECT 3379.715 1193.775 3588.000 1194.615 ;
        RECT 3379.435 1191.395 3588.000 1193.775 ;
        RECT 3379.715 1190.555 3588.000 1191.395 ;
        RECT 3379.435 1188.175 3588.000 1190.555 ;
      LAYER met2 ;
        RECT 3377.035 1187.615 3379.435 1187.895 ;
      LAYER met2 ;
        RECT 3379.715 1187.335 3588.000 1188.175 ;
        RECT 3379.435 1185.415 3588.000 1187.335 ;
      LAYER met2 ;
        RECT 3377.035 1184.855 3379.435 1185.135 ;
      LAYER met2 ;
        RECT 3379.715 1184.575 3588.000 1185.415 ;
        RECT 3379.435 1182.195 3588.000 1184.575 ;
        RECT 3379.715 1181.355 3588.000 1182.195 ;
        RECT 3379.435 1178.975 3588.000 1181.355 ;
      LAYER met2 ;
        RECT 3377.525 1178.695 3377.785 1178.705 ;
        RECT 3377.035 1178.415 3379.435 1178.695 ;
        RECT 3377.525 1178.385 3377.785 1178.415 ;
      LAYER met2 ;
        RECT 3379.715 1178.135 3588.000 1178.975 ;
        RECT 3379.435 1177.085 3588.000 1178.135 ;
        RECT 3379.435 1029.795 3588.000 1030.790 ;
        RECT 3379.715 1028.955 3588.000 1029.795 ;
        RECT 3379.435 1027.035 3588.000 1028.955 ;
        RECT 3379.715 1026.195 3588.000 1027.035 ;
        RECT 3379.435 1023.815 3588.000 1026.195 ;
        RECT 3379.715 1022.975 3588.000 1023.815 ;
        RECT 3379.435 1020.595 3588.000 1022.975 ;
        RECT 3379.715 1019.755 3588.000 1020.595 ;
        RECT 3379.435 1017.835 3588.000 1019.755 ;
        RECT 3379.715 1016.995 3588.000 1017.835 ;
        RECT 3379.435 1014.615 3588.000 1016.995 ;
      LAYER met2 ;
        RECT 3377.035 1014.055 3379.435 1014.335 ;
      LAYER met2 ;
        RECT 3379.715 1013.775 3588.000 1014.615 ;
        RECT 3379.435 1011.395 3588.000 1013.775 ;
        RECT 3379.715 1010.555 3588.000 1011.395 ;
        RECT 3379.435 1008.635 3588.000 1010.555 ;
        RECT 3379.715 1007.795 3588.000 1008.635 ;
        RECT 3379.435 1005.415 3588.000 1007.795 ;
        RECT 3379.715 1004.575 3588.000 1005.415 ;
        RECT 3379.435 1002.195 3588.000 1004.575 ;
        RECT 3379.715 1001.355 3588.000 1002.195 ;
        RECT 3379.435 999.435 3588.000 1001.355 ;
      LAYER met2 ;
        RECT 3377.035 998.875 3379.435 999.155 ;
      LAYER met2 ;
        RECT 3379.715 998.595 3588.000 999.435 ;
        RECT 3379.435 996.215 3588.000 998.595 ;
        RECT 3379.715 995.375 3588.000 996.215 ;
        RECT 3379.435 992.995 3588.000 995.375 ;
      LAYER met2 ;
        RECT 3373.290 992.745 3373.570 992.840 ;
        RECT 3373.255 992.405 3373.570 992.745 ;
        RECT 3377.035 992.435 3379.435 992.715 ;
        RECT 3370.830 961.585 3371.130 961.925 ;
        RECT 3370.330 789.025 3370.640 789.365 ;
        RECT 3369.805 773.845 3370.105 774.185 ;
      LAYER met2 ;
        RECT 4.925 601.390 200.000 625.290 ;
        RECT 4.925 575.395 197.965 601.390 ;
        RECT 198.080 576.895 200.000 578.895 ;
        RECT 4.925 551.495 200.000 575.395 ;
      LAYER met2 ;
        RECT 212.070 561.770 212.595 563.775 ;
      LAYER met2 ;
        RECT 4.925 551.265 197.965 551.495 ;
      LAYER met2 ;
        RECT 3369.830 548.185 3370.080 773.845 ;
        RECT 3370.330 563.365 3370.580 789.025 ;
        RECT 3370.830 736.925 3371.080 961.585 ;
        RECT 3373.290 952.385 3373.570 992.405 ;
      LAYER met2 ;
        RECT 3379.715 992.155 3588.000 992.995 ;
        RECT 3379.435 989.775 3588.000 992.155 ;
        RECT 3379.715 988.935 3588.000 989.775 ;
        RECT 3379.435 987.015 3588.000 988.935 ;
        RECT 3379.715 986.175 3588.000 987.015 ;
        RECT 3379.435 983.795 3588.000 986.175 ;
        RECT 3379.715 982.955 3588.000 983.795 ;
        RECT 3379.435 980.575 3588.000 982.955 ;
        RECT 3379.715 979.735 3588.000 980.575 ;
        RECT 3379.435 977.815 3588.000 979.735 ;
      LAYER met2 ;
        RECT 3377.035 977.255 3379.435 977.535 ;
      LAYER met2 ;
        RECT 3379.715 976.975 3588.000 977.815 ;
        RECT 3379.435 974.595 3588.000 976.975 ;
        RECT 3379.715 973.755 3588.000 974.595 ;
        RECT 3379.435 971.375 3588.000 973.755 ;
      LAYER met2 ;
        RECT 3377.035 970.815 3379.435 971.095 ;
      LAYER met2 ;
        RECT 3379.715 970.535 3588.000 971.375 ;
        RECT 3379.435 968.615 3588.000 970.535 ;
      LAYER met2 ;
        RECT 3377.035 968.055 3379.435 968.335 ;
      LAYER met2 ;
        RECT 3379.715 967.775 3588.000 968.615 ;
        RECT 3379.435 965.395 3588.000 967.775 ;
        RECT 3379.715 964.555 3588.000 965.395 ;
        RECT 3379.435 962.175 3588.000 964.555 ;
      LAYER met2 ;
        RECT 3377.035 961.615 3379.435 961.895 ;
      LAYER met2 ;
        RECT 3379.715 961.335 3588.000 962.175 ;
        RECT 3379.435 959.415 3588.000 961.335 ;
      LAYER met2 ;
        RECT 3377.035 958.855 3379.435 959.135 ;
      LAYER met2 ;
        RECT 3379.715 958.575 3588.000 959.415 ;
        RECT 3379.435 956.195 3588.000 958.575 ;
        RECT 3379.715 955.355 3588.000 956.195 ;
        RECT 3379.435 952.975 3588.000 955.355 ;
      LAYER met2 ;
        RECT 3377.525 952.695 3377.785 952.705 ;
        RECT 3377.035 952.415 3379.435 952.695 ;
        RECT 3377.525 952.385 3377.785 952.415 ;
      LAYER met2 ;
        RECT 3379.715 952.135 3588.000 952.975 ;
        RECT 3379.435 951.085 3588.000 952.135 ;
        RECT 3379.435 804.795 3588.000 805.790 ;
        RECT 3379.715 803.955 3588.000 804.795 ;
        RECT 3379.435 802.035 3588.000 803.955 ;
        RECT 3379.715 801.195 3588.000 802.035 ;
        RECT 3379.435 798.815 3588.000 801.195 ;
        RECT 3379.715 797.975 3588.000 798.815 ;
        RECT 3379.435 795.595 3588.000 797.975 ;
        RECT 3379.715 794.755 3588.000 795.595 ;
        RECT 3379.435 792.835 3588.000 794.755 ;
        RECT 3379.715 791.995 3588.000 792.835 ;
        RECT 3379.435 789.615 3588.000 791.995 ;
      LAYER met2 ;
        RECT 3377.035 789.055 3379.435 789.335 ;
      LAYER met2 ;
        RECT 3379.715 788.775 3588.000 789.615 ;
        RECT 3379.435 786.395 3588.000 788.775 ;
        RECT 3379.715 785.555 3588.000 786.395 ;
        RECT 3379.435 783.635 3588.000 785.555 ;
        RECT 3379.715 782.795 3588.000 783.635 ;
        RECT 3379.435 780.415 3588.000 782.795 ;
        RECT 3379.715 779.575 3588.000 780.415 ;
        RECT 3379.435 777.195 3588.000 779.575 ;
        RECT 3379.715 776.355 3588.000 777.195 ;
        RECT 3379.435 774.435 3588.000 776.355 ;
      LAYER met2 ;
        RECT 3377.035 773.875 3379.435 774.155 ;
      LAYER met2 ;
        RECT 3379.715 773.595 3588.000 774.435 ;
        RECT 3379.435 771.215 3588.000 773.595 ;
        RECT 3379.715 770.375 3588.000 771.215 ;
        RECT 3379.435 767.995 3588.000 770.375 ;
      LAYER met2 ;
        RECT 3373.290 767.745 3373.570 767.840 ;
        RECT 3373.255 767.405 3373.570 767.745 ;
        RECT 3377.035 767.435 3379.435 767.715 ;
        RECT 3370.830 736.585 3371.130 736.925 ;
        RECT 3370.330 563.025 3370.640 563.365 ;
        RECT 3369.805 547.845 3370.105 548.185 ;
      LAYER met2 ;
        RECT 153.765 415.000 158.415 426.140 ;
        RECT 159.640 415.245 163.510 426.195 ;
        RECT 3.570 414.700 197.965 415.000 ;
        RECT 3.570 394.095 198.000 414.700 ;
        RECT 3.570 393.535 197.965 394.095 ;
        RECT 3.570 360.925 198.000 393.535 ;
        RECT 3.570 360.495 197.965 360.925 ;
        RECT 3.570 340.500 198.000 360.495 ;
      LAYER met2 ;
        RECT 211.050 347.125 211.480 349.935 ;
      LAYER met2 ;
        RECT 3.570 340.490 197.965 340.500 ;
      LAYER met2 ;
        RECT 2856.605 212.915 2858.820 214.920 ;
        RECT 211.575 212.320 211.905 212.720 ;
        RECT 212.910 212.320 213.670 212.350 ;
        RECT 211.575 212.060 213.670 212.320 ;
        RECT 212.910 212.030 213.670 212.060 ;
        RECT 454.315 210.870 455.470 211.225 ;
        RECT 665.020 201.170 665.260 201.190 ;
        RECT 664.990 200.850 665.260 201.170 ;
        RECT 665.020 200.000 665.260 200.850 ;
      LAYER met2 ;
        RECT 394.710 197.965 418.610 200.000 ;
        RECT 441.105 198.080 443.105 200.000 ;
        RECT 444.605 197.965 468.505 200.000 ;
        RECT 663.085 199.390 664.485 200.000 ;
      LAYER met2 ;
        RECT 664.765 199.670 665.785 200.000 ;
      LAYER met2 ;
        RECT 666.065 199.390 704.700 200.000 ;
        RECT 663.085 199.080 704.700 199.390 ;
      LAYER met2 ;
        RECT 704.980 199.360 705.240 212.350 ;
        RECT 712.850 200.610 713.110 212.500 ;
        RECT 715.375 212.345 715.635 212.350 ;
        RECT 712.820 200.350 713.140 200.610 ;
      LAYER met2 ;
        RECT 705.520 199.390 706.565 200.000 ;
      LAYER met2 ;
        RECT 706.845 199.670 707.495 200.000 ;
      LAYER met2 ;
        RECT 707.775 199.390 708.055 200.000 ;
        RECT 709.345 199.390 709.490 200.000 ;
      LAYER met2 ;
        RECT 709.770 199.670 710.420 200.000 ;
      LAYER met2 ;
        RECT 710.700 199.390 715.060 200.000 ;
        RECT 705.520 199.080 715.060 199.390 ;
        RECT 394.710 4.925 468.735 197.965 ;
        RECT 663.085 196.020 715.060 199.080 ;
        RECT 663.085 195.735 714.775 196.020 ;
      LAYER met2 ;
        RECT 715.340 195.755 715.640 212.345 ;
        RECT 717.145 201.600 717.425 212.420 ;
        RECT 717.100 201.320 717.470 201.600 ;
        RECT 719.625 200.850 719.885 201.170 ;
        RECT 719.660 200.000 719.850 200.850 ;
        RECT 723.005 200.000 723.275 212.415 ;
        RECT 979.875 211.705 980.155 211.840 ;
        RECT 979.875 211.385 980.170 211.705 ;
        RECT 729.265 200.000 729.535 210.710 ;
        RECT 933.415 208.565 933.695 210.965 ;
        RECT 939.855 208.565 940.135 210.965 ;
        RECT 942.615 208.565 942.895 210.965 ;
        RECT 945.835 208.565 946.115 210.965 ;
        RECT 949.055 208.565 949.335 210.965 ;
        RECT 951.815 208.565 952.095 210.965 ;
        RECT 955.035 208.565 955.315 210.965 ;
        RECT 958.255 208.565 958.535 210.965 ;
        RECT 961.015 210.205 961.295 210.965 ;
        RECT 964.235 210.705 964.515 210.965 ;
        RECT 964.230 210.385 964.515 210.705 ;
        RECT 961.000 209.885 961.295 210.205 ;
        RECT 961.015 208.565 961.295 209.885 ;
        RECT 964.235 208.565 964.515 210.385 ;
        RECT 967.455 210.205 967.735 210.965 ;
        RECT 967.455 209.885 967.760 210.205 ;
        RECT 967.455 208.565 967.735 209.885 ;
        RECT 973.435 208.565 973.715 210.965 ;
        RECT 979.875 208.565 980.155 211.385 ;
        RECT 995.055 211.205 995.335 211.320 ;
        RECT 982.635 210.205 982.915 210.965 ;
        RECT 982.620 209.885 982.915 210.205 ;
        RECT 982.635 208.565 982.915 209.885 ;
        RECT 985.855 210.205 986.135 210.965 ;
        RECT 985.855 209.885 986.140 210.205 ;
        RECT 985.855 208.565 986.135 209.885 ;
        RECT 989.075 208.565 989.355 210.965 ;
        RECT 991.835 210.205 992.115 210.965 ;
        RECT 995.055 210.885 995.370 211.205 ;
        RECT 991.835 209.885 992.130 210.205 ;
        RECT 991.835 208.565 992.115 209.885 ;
        RECT 995.055 208.565 995.335 210.885 ;
        RECT 1001.035 210.205 1001.315 210.965 ;
        RECT 1001.035 209.885 1001.330 210.205 ;
        RECT 1001.035 208.565 1001.315 209.885 ;
        RECT 1004.255 208.565 1004.535 210.965 ;
        RECT 1007.475 210.705 1007.755 210.965 ;
        RECT 1007.460 210.385 1007.755 210.705 ;
        RECT 1007.475 208.565 1007.755 210.385 ;
        RECT 1010.235 208.565 1010.515 210.965 ;
        RECT 1268.065 209.755 1269.135 210.215 ;
        RECT 1476.415 208.565 1476.695 212.840 ;
        RECT 1479.635 208.565 1479.915 210.965 ;
        RECT 1482.855 208.565 1483.135 210.965 ;
        RECT 1485.615 208.565 1485.895 210.965 ;
        RECT 1488.835 208.565 1489.115 210.965 ;
        RECT 1492.055 208.565 1492.335 210.965 ;
        RECT 1494.815 208.565 1495.095 210.965 ;
        RECT 1498.035 208.565 1498.315 210.965 ;
        RECT 1501.255 208.565 1501.535 210.965 ;
        RECT 1504.015 210.205 1504.295 210.965 ;
        RECT 1504.000 209.885 1504.295 210.205 ;
        RECT 1504.015 208.565 1504.295 209.885 ;
        RECT 1507.235 208.565 1507.515 210.965 ;
        RECT 1510.455 210.205 1510.735 210.965 ;
        RECT 1510.455 209.885 1510.760 210.205 ;
        RECT 1510.455 208.565 1510.735 209.885 ;
        RECT 1516.435 208.565 1516.715 212.840 ;
        RECT 1522.875 211.705 1523.155 211.815 ;
        RECT 1522.875 211.385 1523.170 211.705 ;
        RECT 1522.875 208.565 1523.155 211.385 ;
        RECT 1538.055 211.210 1538.340 211.230 ;
        RECT 1525.635 210.205 1525.915 210.965 ;
        RECT 1525.620 209.885 1525.915 210.205 ;
        RECT 1525.635 208.565 1525.915 209.885 ;
        RECT 1528.855 208.565 1529.135 210.965 ;
        RECT 1532.075 208.565 1532.355 210.965 ;
        RECT 1538.050 210.880 1538.340 211.210 ;
        RECT 1538.055 208.565 1538.335 210.880 ;
        RECT 1544.035 210.205 1544.315 210.965 ;
        RECT 1544.035 209.885 1544.330 210.205 ;
        RECT 1544.035 208.565 1544.315 209.885 ;
        RECT 1547.255 208.565 1547.535 210.965 ;
        RECT 1553.235 208.565 1553.515 210.965 ;
        RECT 1750.415 208.565 1750.695 212.840 ;
        RECT 1753.635 208.565 1753.915 210.965 ;
        RECT 1756.855 208.565 1757.135 210.965 ;
        RECT 1759.615 208.565 1759.895 210.965 ;
        RECT 1762.835 208.565 1763.115 210.965 ;
        RECT 1766.055 208.565 1766.335 210.965 ;
        RECT 1768.815 208.565 1769.095 210.965 ;
        RECT 1772.035 208.565 1772.315 210.965 ;
        RECT 1775.255 208.565 1775.535 210.965 ;
        RECT 1778.015 210.205 1778.295 210.965 ;
        RECT 1778.000 209.885 1778.295 210.205 ;
        RECT 1778.015 208.565 1778.295 209.885 ;
        RECT 1781.235 208.565 1781.515 210.965 ;
        RECT 1784.455 210.205 1784.735 210.965 ;
        RECT 1784.455 209.885 1784.760 210.205 ;
        RECT 1784.455 208.565 1784.735 209.885 ;
        RECT 1790.435 208.565 1790.715 212.840 ;
        RECT 1796.875 211.705 1797.155 211.815 ;
        RECT 1796.875 211.385 1797.170 211.705 ;
        RECT 1796.875 208.565 1797.155 211.385 ;
        RECT 1812.055 211.210 1812.340 211.230 ;
        RECT 1799.635 210.205 1799.915 210.965 ;
        RECT 1799.620 209.885 1799.915 210.205 ;
        RECT 1799.635 208.565 1799.915 209.885 ;
        RECT 1802.855 208.565 1803.135 210.965 ;
        RECT 1806.075 208.565 1806.355 210.965 ;
        RECT 1812.050 210.880 1812.340 211.210 ;
        RECT 1812.055 208.565 1812.335 210.880 ;
        RECT 1818.035 210.205 1818.315 210.965 ;
        RECT 1818.035 209.885 1818.330 210.205 ;
        RECT 1818.035 208.565 1818.315 209.885 ;
        RECT 1821.255 208.565 1821.535 210.965 ;
        RECT 1827.235 208.565 1827.515 210.965 ;
        RECT 2024.415 208.565 2024.695 212.840 ;
        RECT 2030.855 208.565 2031.135 210.965 ;
        RECT 2033.615 208.565 2033.895 210.965 ;
        RECT 2036.835 208.565 2037.115 210.965 ;
        RECT 2040.055 208.565 2040.335 210.965 ;
        RECT 2042.815 208.565 2043.095 210.965 ;
        RECT 2049.255 208.565 2049.535 210.965 ;
        RECT 2052.015 210.205 2052.295 210.965 ;
        RECT 2052.000 209.885 2052.295 210.205 ;
        RECT 2052.015 208.565 2052.295 209.885 ;
        RECT 2058.455 210.205 2058.735 210.965 ;
        RECT 2058.455 209.885 2058.760 210.205 ;
        RECT 2058.455 208.565 2058.735 209.885 ;
        RECT 2064.435 208.565 2064.715 212.840 ;
        RECT 2618.875 212.575 2619.155 212.710 ;
        RECT 3369.830 212.575 3370.080 547.845 ;
        RECT 3370.330 213.215 3370.580 563.025 ;
        RECT 3370.830 510.925 3371.080 736.585 ;
        RECT 3373.290 727.385 3373.570 767.405 ;
      LAYER met2 ;
        RECT 3379.715 767.155 3588.000 767.995 ;
        RECT 3379.435 764.775 3588.000 767.155 ;
        RECT 3379.715 763.935 3588.000 764.775 ;
        RECT 3379.435 762.015 3588.000 763.935 ;
        RECT 3379.715 761.175 3588.000 762.015 ;
        RECT 3379.435 758.795 3588.000 761.175 ;
        RECT 3379.715 757.955 3588.000 758.795 ;
        RECT 3379.435 755.575 3588.000 757.955 ;
        RECT 3379.715 754.735 3588.000 755.575 ;
        RECT 3379.435 752.815 3588.000 754.735 ;
      LAYER met2 ;
        RECT 3377.035 752.255 3379.435 752.535 ;
      LAYER met2 ;
        RECT 3379.715 751.975 3588.000 752.815 ;
        RECT 3379.435 749.595 3588.000 751.975 ;
        RECT 3379.715 748.755 3588.000 749.595 ;
        RECT 3379.435 746.375 3588.000 748.755 ;
      LAYER met2 ;
        RECT 3377.035 745.815 3379.435 746.095 ;
      LAYER met2 ;
        RECT 3379.715 745.535 3588.000 746.375 ;
        RECT 3379.435 743.615 3588.000 745.535 ;
      LAYER met2 ;
        RECT 3377.035 743.055 3379.435 743.335 ;
      LAYER met2 ;
        RECT 3379.715 742.775 3588.000 743.615 ;
        RECT 3379.435 740.395 3588.000 742.775 ;
        RECT 3379.715 739.555 3588.000 740.395 ;
        RECT 3379.435 737.175 3588.000 739.555 ;
      LAYER met2 ;
        RECT 3377.035 736.615 3379.435 736.895 ;
      LAYER met2 ;
        RECT 3379.715 736.335 3588.000 737.175 ;
        RECT 3379.435 734.415 3588.000 736.335 ;
      LAYER met2 ;
        RECT 3377.035 733.855 3379.435 734.135 ;
      LAYER met2 ;
        RECT 3379.715 733.575 3588.000 734.415 ;
        RECT 3379.435 731.195 3588.000 733.575 ;
        RECT 3379.715 730.355 3588.000 731.195 ;
        RECT 3379.435 727.975 3588.000 730.355 ;
      LAYER met2 ;
        RECT 3377.525 727.695 3377.785 727.705 ;
        RECT 3377.035 727.415 3379.435 727.695 ;
        RECT 3377.525 727.385 3377.785 727.415 ;
      LAYER met2 ;
        RECT 3379.715 727.135 3588.000 727.975 ;
        RECT 3379.435 726.085 3588.000 727.135 ;
        RECT 3379.435 578.795 3588.000 579.790 ;
        RECT 3379.715 577.955 3588.000 578.795 ;
        RECT 3379.435 576.035 3588.000 577.955 ;
        RECT 3379.715 575.195 3588.000 576.035 ;
        RECT 3379.435 572.815 3588.000 575.195 ;
        RECT 3379.715 571.975 3588.000 572.815 ;
        RECT 3379.435 569.595 3588.000 571.975 ;
        RECT 3379.715 568.755 3588.000 569.595 ;
        RECT 3379.435 566.835 3588.000 568.755 ;
        RECT 3379.715 565.995 3588.000 566.835 ;
        RECT 3379.435 563.615 3588.000 565.995 ;
      LAYER met2 ;
        RECT 3377.035 563.055 3379.435 563.335 ;
      LAYER met2 ;
        RECT 3379.715 562.775 3588.000 563.615 ;
        RECT 3379.435 560.395 3588.000 562.775 ;
        RECT 3379.715 559.555 3588.000 560.395 ;
        RECT 3379.435 557.635 3588.000 559.555 ;
        RECT 3379.715 556.795 3588.000 557.635 ;
        RECT 3379.435 554.415 3588.000 556.795 ;
        RECT 3379.715 553.575 3588.000 554.415 ;
        RECT 3379.435 551.195 3588.000 553.575 ;
        RECT 3379.715 550.355 3588.000 551.195 ;
        RECT 3379.435 548.435 3588.000 550.355 ;
      LAYER met2 ;
        RECT 3377.035 547.875 3379.435 548.155 ;
      LAYER met2 ;
        RECT 3379.715 547.595 3588.000 548.435 ;
        RECT 3379.435 545.215 3588.000 547.595 ;
        RECT 3379.715 544.375 3588.000 545.215 ;
        RECT 3379.435 541.995 3588.000 544.375 ;
      LAYER met2 ;
        RECT 3373.290 541.745 3373.570 541.840 ;
        RECT 3373.255 541.405 3373.570 541.745 ;
        RECT 3377.035 541.435 3379.435 541.715 ;
        RECT 3370.830 510.585 3371.130 510.925 ;
        RECT 3370.330 212.895 3370.615 213.215 ;
        RECT 3370.330 212.850 3370.580 212.895 ;
        RECT 2618.875 212.255 2619.170 212.575 ;
        RECT 3369.830 212.255 3370.090 212.575 ;
        RECT 2070.875 211.705 2071.155 211.840 ;
        RECT 2344.875 211.705 2345.155 211.840 ;
        RECT 2070.875 211.385 2071.170 211.705 ;
        RECT 2344.875 211.385 2345.170 211.705 ;
        RECT 2070.875 208.565 2071.155 211.385 ;
        RECT 2086.055 211.210 2086.340 211.230 ;
        RECT 2073.635 210.205 2073.915 210.965 ;
        RECT 2073.620 209.885 2073.915 210.205 ;
        RECT 2073.635 208.565 2073.915 209.885 ;
        RECT 2080.075 208.565 2080.355 210.965 ;
        RECT 2086.050 210.880 2086.340 211.210 ;
        RECT 2086.055 208.565 2086.335 210.880 ;
        RECT 2092.035 210.205 2092.315 210.965 ;
        RECT 2092.035 209.885 2092.330 210.205 ;
        RECT 2092.035 208.565 2092.315 209.885 ;
        RECT 2095.255 208.565 2095.535 210.965 ;
        RECT 2101.235 208.565 2101.515 210.965 ;
        RECT 2298.415 208.565 2298.695 210.965 ;
        RECT 2304.855 208.565 2305.135 210.965 ;
        RECT 2307.615 208.565 2307.895 210.965 ;
        RECT 2310.835 208.565 2311.115 210.965 ;
        RECT 2314.055 208.565 2314.335 210.965 ;
        RECT 2316.815 208.565 2317.095 210.965 ;
        RECT 2323.255 208.565 2323.535 210.965 ;
        RECT 2326.015 210.205 2326.295 210.965 ;
        RECT 2326.000 209.885 2326.295 210.205 ;
        RECT 2326.015 208.565 2326.295 209.885 ;
        RECT 2332.455 210.205 2332.735 210.965 ;
        RECT 2332.455 209.885 2332.760 210.205 ;
        RECT 2332.455 208.565 2332.735 209.885 ;
        RECT 2338.435 208.565 2338.715 210.965 ;
        RECT 2344.875 208.565 2345.155 211.385 ;
        RECT 2360.055 211.210 2360.340 211.230 ;
        RECT 2347.635 210.205 2347.915 210.965 ;
        RECT 2347.620 209.885 2347.915 210.205 ;
        RECT 2347.635 208.565 2347.915 209.885 ;
        RECT 2354.075 208.565 2354.355 210.965 ;
        RECT 2360.050 210.880 2360.340 211.210 ;
        RECT 2360.055 208.565 2360.335 210.880 ;
        RECT 2366.035 210.205 2366.315 210.965 ;
        RECT 2366.035 209.885 2366.330 210.205 ;
        RECT 2366.035 208.565 2366.315 209.885 ;
        RECT 2369.255 208.565 2369.535 210.965 ;
        RECT 2375.235 208.565 2375.515 210.965 ;
        RECT 2572.415 208.565 2572.695 210.965 ;
        RECT 2578.855 208.565 2579.135 210.965 ;
        RECT 2581.615 208.565 2581.895 211.610 ;
        RECT 2584.840 210.965 2585.100 211.075 ;
        RECT 2600.000 210.965 2600.260 211.075 ;
        RECT 2606.500 210.965 2606.760 211.075 ;
        RECT 2584.835 208.565 2585.115 210.965 ;
        RECT 2588.055 208.565 2588.335 210.965 ;
        RECT 2590.815 208.565 2591.095 210.965 ;
        RECT 2597.255 208.565 2597.535 210.965 ;
        RECT 2600.000 210.755 2600.295 210.965 ;
        RECT 2600.015 208.565 2600.295 210.755 ;
        RECT 2606.455 210.755 2606.760 210.965 ;
        RECT 2606.455 208.565 2606.735 210.755 ;
        RECT 2612.435 208.565 2612.715 210.965 ;
        RECT 2618.875 208.565 2619.155 212.255 ;
        RECT 3369.830 212.155 3370.080 212.255 ;
        RECT 2634.055 212.080 2634.340 212.100 ;
        RECT 2634.050 211.750 2634.340 212.080 ;
        RECT 2621.620 210.965 2621.880 211.075 ;
        RECT 2628.080 210.965 2628.340 211.075 ;
        RECT 2621.620 210.755 2621.915 210.965 ;
        RECT 2621.635 208.565 2621.915 210.755 ;
        RECT 2628.075 208.565 2628.355 210.965 ;
        RECT 2634.055 208.565 2634.335 211.750 ;
        RECT 3370.830 211.575 3371.080 510.585 ;
        RECT 3373.290 501.385 3373.570 541.405 ;
      LAYER met2 ;
        RECT 3379.715 541.155 3588.000 541.995 ;
        RECT 3379.435 538.775 3588.000 541.155 ;
        RECT 3379.715 537.935 3588.000 538.775 ;
        RECT 3379.435 536.015 3588.000 537.935 ;
        RECT 3379.715 535.175 3588.000 536.015 ;
        RECT 3379.435 532.795 3588.000 535.175 ;
        RECT 3379.715 531.955 3588.000 532.795 ;
        RECT 3379.435 529.575 3588.000 531.955 ;
        RECT 3379.715 528.735 3588.000 529.575 ;
        RECT 3379.435 526.815 3588.000 528.735 ;
      LAYER met2 ;
        RECT 3377.035 526.255 3379.435 526.535 ;
      LAYER met2 ;
        RECT 3379.715 525.975 3588.000 526.815 ;
        RECT 3379.435 523.595 3588.000 525.975 ;
        RECT 3379.715 522.755 3588.000 523.595 ;
        RECT 3379.435 520.375 3588.000 522.755 ;
      LAYER met2 ;
        RECT 3377.035 519.815 3379.435 520.095 ;
      LAYER met2 ;
        RECT 3379.715 519.535 3588.000 520.375 ;
        RECT 3379.435 517.615 3588.000 519.535 ;
      LAYER met2 ;
        RECT 3377.035 517.055 3379.435 517.335 ;
      LAYER met2 ;
        RECT 3379.715 516.775 3588.000 517.615 ;
        RECT 3379.435 514.395 3588.000 516.775 ;
        RECT 3379.715 513.555 3588.000 514.395 ;
        RECT 3379.435 511.175 3588.000 513.555 ;
      LAYER met2 ;
        RECT 3377.035 510.615 3379.435 510.895 ;
      LAYER met2 ;
        RECT 3379.715 510.335 3588.000 511.175 ;
        RECT 3379.435 508.415 3588.000 510.335 ;
      LAYER met2 ;
        RECT 3377.035 507.855 3379.435 508.135 ;
      LAYER met2 ;
        RECT 3379.715 507.575 3588.000 508.415 ;
        RECT 3379.435 505.195 3588.000 507.575 ;
        RECT 3379.715 504.355 3588.000 505.195 ;
        RECT 3379.435 501.975 3588.000 504.355 ;
      LAYER met2 ;
        RECT 3377.525 501.695 3377.785 501.705 ;
        RECT 3377.035 501.415 3379.435 501.695 ;
        RECT 3377.525 501.385 3377.785 501.415 ;
      LAYER met2 ;
        RECT 3379.715 501.135 3588.000 501.975 ;
        RECT 3379.435 500.085 3588.000 501.135 ;
      LAYER met2 ;
        RECT 3370.830 211.255 3371.090 211.575 ;
        RECT 3370.830 211.215 3371.080 211.255 ;
        RECT 2640.070 210.965 2640.330 211.075 ;
        RECT 2643.260 210.965 2643.520 211.075 ;
        RECT 2640.035 210.755 2640.330 210.965 ;
        RECT 2640.035 208.565 2640.315 210.755 ;
        RECT 2643.255 208.565 2643.535 210.965 ;
        RECT 2649.235 208.565 2649.515 210.965 ;
      LAYER met2 ;
        RECT 932.085 208.285 933.135 208.565 ;
        RECT 933.975 208.285 936.355 208.565 ;
        RECT 937.195 208.285 939.575 208.565 ;
        RECT 940.415 208.285 942.335 208.565 ;
        RECT 943.175 208.285 945.555 208.565 ;
        RECT 946.395 208.285 948.775 208.565 ;
        RECT 949.615 208.285 951.535 208.565 ;
        RECT 952.375 208.285 954.755 208.565 ;
        RECT 955.595 208.285 957.975 208.565 ;
        RECT 958.815 208.285 960.735 208.565 ;
        RECT 961.575 208.285 963.955 208.565 ;
        RECT 964.795 208.285 967.175 208.565 ;
        RECT 968.015 208.285 969.935 208.565 ;
        RECT 970.775 208.285 973.155 208.565 ;
        RECT 973.995 208.285 976.375 208.565 ;
        RECT 977.215 208.285 979.595 208.565 ;
        RECT 980.435 208.285 982.355 208.565 ;
        RECT 983.195 208.285 985.575 208.565 ;
        RECT 986.415 208.285 988.795 208.565 ;
        RECT 989.635 208.285 991.555 208.565 ;
        RECT 992.395 208.285 994.775 208.565 ;
        RECT 995.615 208.285 997.995 208.565 ;
        RECT 998.835 208.285 1000.755 208.565 ;
        RECT 1001.595 208.285 1003.975 208.565 ;
        RECT 1004.815 208.285 1007.195 208.565 ;
        RECT 1008.035 208.285 1009.955 208.565 ;
        RECT 1010.795 208.285 1011.790 208.565 ;
        RECT 715.920 198.310 716.495 200.000 ;
      LAYER met2 ;
        RECT 716.775 198.590 717.925 200.000 ;
      LAYER met2 ;
        RECT 718.205 199.155 718.810 200.000 ;
      LAYER met2 ;
        RECT 719.090 199.435 720.755 200.000 ;
      LAYER met2 ;
        RECT 721.035 199.155 722.585 200.000 ;
        RECT 718.205 198.735 722.585 199.155 ;
      LAYER met2 ;
        RECT 722.865 199.015 723.445 200.000 ;
      LAYER met2 ;
        RECT 723.725 198.735 725.175 200.000 ;
        RECT 718.205 198.310 725.175 198.735 ;
        RECT 715.920 198.250 725.175 198.310 ;
        RECT 725.995 199.390 728.825 200.000 ;
      LAYER met2 ;
        RECT 729.105 199.670 729.575 200.000 ;
      LAYER met2 ;
        RECT 729.855 199.390 737.660 200.000 ;
        RECT 725.995 198.250 737.660 199.390 ;
        RECT 715.920 196.845 737.660 198.250 ;
        RECT 715.920 196.485 722.475 196.845 ;
        RECT 727.600 196.705 737.660 196.845 ;
        RECT 715.920 196.215 722.205 196.485 ;
      LAYER met2 ;
        RECT 722.755 196.425 727.320 196.565 ;
        RECT 722.755 196.355 727.650 196.425 ;
      LAYER met2 ;
        RECT 727.930 196.375 737.660 196.705 ;
      LAYER met2 ;
        RECT 722.755 196.305 727.180 196.355 ;
      LAYER met2 ;
        RECT 715.920 196.035 721.835 196.215 ;
      LAYER met2 ;
        RECT 722.755 196.205 723.115 196.305 ;
        RECT 723.125 196.205 723.225 196.305 ;
        RECT 727.070 196.235 727.305 196.305 ;
        RECT 727.320 196.235 727.650 196.355 ;
      LAYER met2 ;
        RECT 716.220 195.845 721.835 196.035 ;
      LAYER met2 ;
        RECT 722.485 196.165 722.755 196.205 ;
        RECT 722.855 196.165 723.125 196.205 ;
        RECT 722.485 196.025 723.125 196.165 ;
        RECT 727.070 196.095 727.650 196.235 ;
        RECT 727.070 196.070 727.305 196.095 ;
        RECT 722.485 195.935 722.755 196.025 ;
        RECT 722.855 195.935 723.125 196.025 ;
        RECT 715.340 195.740 715.940 195.755 ;
      LAYER met2 ;
        RECT 663.085 195.380 708.600 195.735 ;
      LAYER met2 ;
        RECT 715.055 195.455 715.940 195.740 ;
      LAYER met2 ;
        RECT 716.220 195.735 721.725 195.845 ;
      LAYER met2 ;
        RECT 722.115 195.565 722.855 195.935 ;
      LAYER met2 ;
        RECT 723.505 195.925 726.790 196.025 ;
        RECT 723.405 195.790 726.790 195.925 ;
      LAYER met2 ;
        RECT 727.305 195.955 727.625 196.070 ;
        RECT 727.650 195.955 727.995 196.095 ;
      LAYER met2 ;
        RECT 728.275 196.030 737.660 196.375 ;
      LAYER met2 ;
        RECT 727.305 195.815 727.995 195.955 ;
      LAYER met2 ;
        RECT 723.405 195.655 727.025 195.790 ;
      LAYER met2 ;
        RECT 727.305 195.750 727.625 195.815 ;
        RECT 727.650 195.750 727.995 195.815 ;
        RECT 722.005 195.455 722.485 195.565 ;
      LAYER met2 ;
        RECT 663.085 195.050 708.270 195.380 ;
      LAYER met2 ;
        RECT 708.880 195.315 722.485 195.455 ;
        RECT 708.880 195.245 709.235 195.315 ;
        RECT 715.340 195.245 715.640 195.315 ;
        RECT 722.115 195.245 722.485 195.315 ;
      LAYER met2 ;
        RECT 723.135 195.470 727.025 195.655 ;
      LAYER met2 ;
        RECT 727.625 195.675 727.955 195.750 ;
        RECT 727.995 195.675 728.265 195.750 ;
      LAYER met2 ;
        RECT 723.135 195.285 727.345 195.470 ;
      LAYER met2 ;
        RECT 727.625 195.425 728.265 195.675 ;
        RECT 727.625 195.420 727.955 195.425 ;
        RECT 708.880 195.195 722.485 195.245 ;
        RECT 708.880 195.100 709.235 195.195 ;
        RECT 709.250 195.100 709.345 195.195 ;
      LAYER met2 ;
        RECT 722.765 195.140 727.345 195.285 ;
      LAYER met2 ;
        RECT 708.550 195.055 708.880 195.100 ;
        RECT 708.920 195.055 709.250 195.100 ;
      LAYER met2 ;
        RECT 663.085 189.305 708.140 195.050 ;
      LAYER met2 ;
        RECT 708.550 194.845 709.250 195.055 ;
      LAYER met2 ;
        RECT 722.765 194.915 727.725 195.140 ;
      LAYER met2 ;
        RECT 708.550 194.770 708.880 194.845 ;
        RECT 708.920 194.770 709.250 194.845 ;
      LAYER met2 ;
        RECT 709.625 194.820 727.725 194.915 ;
      LAYER met2 ;
        RECT 708.420 194.640 708.550 194.770 ;
        RECT 708.680 194.640 708.920 194.770 ;
        RECT 708.420 194.530 708.920 194.640 ;
      LAYER met2 ;
        RECT 663.085 189.115 707.950 189.305 ;
        RECT 663.085 184.635 707.690 189.115 ;
      LAYER met2 ;
        RECT 708.420 189.025 708.680 194.530 ;
      LAYER met2 ;
        RECT 709.530 194.490 727.725 194.820 ;
        RECT 709.200 194.250 727.725 194.490 ;
      LAYER met2 ;
        RECT 708.230 188.915 708.680 189.025 ;
        RECT 708.230 188.835 708.420 188.915 ;
        RECT 708.600 188.835 708.680 188.915 ;
      LAYER met2 ;
        RECT 708.960 191.420 727.725 194.250 ;
        RECT 708.960 191.080 727.385 191.420 ;
      LAYER met2 ;
        RECT 728.005 191.140 728.265 195.425 ;
      LAYER met2 ;
        RECT 708.960 190.880 727.185 191.080 ;
      LAYER met2 ;
        RECT 727.665 190.890 728.265 191.140 ;
      LAYER met2 ;
        RECT 708.960 190.550 726.855 190.880 ;
      LAYER met2 ;
        RECT 727.665 190.800 728.005 190.890 ;
        RECT 728.035 190.800 728.265 190.890 ;
        RECT 727.465 190.750 727.665 190.800 ;
        RECT 727.835 190.750 728.035 190.800 ;
        RECT 727.465 190.680 728.035 190.750 ;
        RECT 727.465 190.600 727.665 190.680 ;
        RECT 727.835 190.600 728.035 190.680 ;
        RECT 707.970 188.465 708.600 188.835 ;
      LAYER met2 ;
        RECT 708.960 188.555 726.595 190.550 ;
      LAYER met2 ;
        RECT 727.135 190.540 727.465 190.600 ;
        RECT 727.505 190.540 727.835 190.600 ;
        RECT 727.135 190.400 727.835 190.540 ;
      LAYER met2 ;
        RECT 728.545 190.520 737.660 196.030 ;
      LAYER met2 ;
        RECT 727.135 190.270 727.465 190.400 ;
        RECT 727.505 190.270 727.835 190.400 ;
      LAYER met2 ;
        RECT 728.315 190.320 737.660 190.520 ;
        RECT 663.085 184.300 707.355 184.635 ;
      LAYER met2 ;
        RECT 707.970 184.355 708.230 188.465 ;
      LAYER met2 ;
        RECT 708.880 188.185 726.595 188.555 ;
        RECT 663.085 179.225 707.095 184.300 ;
      LAYER met2 ;
        RECT 707.635 184.105 708.230 184.355 ;
        RECT 707.635 184.020 707.970 184.105 ;
        RECT 708.005 184.020 708.230 184.105 ;
        RECT 707.375 183.650 708.005 184.020 ;
      LAYER met2 ;
        RECT 708.510 183.740 726.595 188.185 ;
      LAYER met2 ;
        RECT 707.375 179.505 707.635 183.650 ;
      LAYER met2 ;
        RECT 708.285 183.370 726.595 183.740 ;
        RECT 707.915 179.225 726.595 183.370 ;
        RECT 663.085 172.420 726.595 179.225 ;
      LAYER met2 ;
        RECT 726.875 189.900 727.505 190.270 ;
      LAYER met2 ;
        RECT 728.115 189.990 737.660 190.320 ;
      LAYER met2 ;
        RECT 726.875 173.390 727.135 189.900 ;
      LAYER met2 ;
        RECT 727.785 189.620 737.660 189.990 ;
        RECT 727.415 173.670 737.660 189.620 ;
      LAYER met2 ;
        RECT 726.875 172.700 727.350 173.390 ;
      LAYER met2 ;
        RECT 663.085 172.345 726.810 172.420 ;
        RECT 663.085 169.195 726.595 172.345 ;
      LAYER met2 ;
        RECT 727.090 172.065 727.350 172.700 ;
        RECT 726.875 171.855 727.350 172.065 ;
        RECT 726.875 171.850 727.090 171.855 ;
        RECT 726.875 171.375 727.350 171.850 ;
      LAYER met2 ;
        RECT 663.085 169.050 726.450 169.195 ;
        RECT 663.085 168.825 726.225 169.050 ;
      LAYER met2 ;
        RECT 726.875 168.915 727.135 171.375 ;
      LAYER met2 ;
        RECT 727.630 171.095 737.660 173.670 ;
        RECT 663.085 164.260 726.200 168.825 ;
      LAYER met2 ;
        RECT 726.730 168.770 727.135 168.915 ;
        RECT 726.505 168.735 726.730 168.770 ;
        RECT 726.875 168.735 727.135 168.770 ;
        RECT 726.505 168.665 727.135 168.735 ;
        RECT 726.505 168.545 726.730 168.665 ;
        RECT 726.875 168.545 727.135 168.665 ;
        RECT 726.480 168.520 726.505 168.545 ;
        RECT 726.740 168.520 726.875 168.545 ;
        RECT 726.480 168.410 726.875 168.520 ;
      LAYER met2 ;
        RECT 663.085 163.440 725.570 164.260 ;
      LAYER met2 ;
        RECT 726.480 163.980 726.740 168.410 ;
      LAYER met2 ;
        RECT 727.415 168.265 737.660 171.095 ;
        RECT 727.155 168.130 737.660 168.265 ;
      LAYER met2 ;
        RECT 725.850 163.720 726.740 163.980 ;
      LAYER met2 ;
        RECT 727.020 163.440 737.660 168.130 ;
        RECT 663.085 0.790 737.660 163.440 ;
        RECT 932.085 0.000 1011.790 208.285 ;
        RECT 1475.085 208.285 1476.135 208.565 ;
        RECT 1476.975 208.285 1479.355 208.565 ;
        RECT 1480.195 208.285 1482.575 208.565 ;
        RECT 1483.415 208.285 1485.335 208.565 ;
        RECT 1486.175 208.285 1488.555 208.565 ;
        RECT 1489.395 208.285 1491.775 208.565 ;
        RECT 1492.615 208.285 1494.535 208.565 ;
        RECT 1495.375 208.285 1497.755 208.565 ;
        RECT 1498.595 208.285 1500.975 208.565 ;
        RECT 1501.815 208.285 1503.735 208.565 ;
        RECT 1504.575 208.285 1506.955 208.565 ;
        RECT 1507.795 208.285 1510.175 208.565 ;
        RECT 1511.015 208.285 1512.935 208.565 ;
        RECT 1513.775 208.285 1516.155 208.565 ;
        RECT 1516.995 208.285 1519.375 208.565 ;
        RECT 1520.215 208.285 1522.595 208.565 ;
        RECT 1523.435 208.285 1525.355 208.565 ;
        RECT 1526.195 208.285 1528.575 208.565 ;
        RECT 1529.415 208.285 1531.795 208.565 ;
        RECT 1532.635 208.285 1534.555 208.565 ;
        RECT 1535.395 208.285 1537.775 208.565 ;
        RECT 1538.615 208.285 1540.995 208.565 ;
        RECT 1541.835 208.285 1543.755 208.565 ;
        RECT 1544.595 208.285 1546.975 208.565 ;
        RECT 1547.815 208.285 1550.195 208.565 ;
        RECT 1551.035 208.285 1552.955 208.565 ;
        RECT 1553.795 208.285 1554.790 208.565 ;
        RECT 1206.300 197.965 1226.905 198.000 ;
        RECT 1227.465 197.965 1260.075 198.000 ;
        RECT 1260.505 197.965 1280.500 198.000 ;
        RECT 1194.805 159.640 1205.755 163.510 ;
        RECT 1206.000 158.415 1280.500 197.965 ;
        RECT 1194.860 153.765 1280.500 158.415 ;
        RECT 1206.000 3.570 1280.500 153.765 ;
        RECT 1475.085 0.000 1554.790 208.285 ;
        RECT 1749.085 208.285 1750.135 208.565 ;
        RECT 1750.975 208.285 1753.355 208.565 ;
        RECT 1754.195 208.285 1756.575 208.565 ;
        RECT 1757.415 208.285 1759.335 208.565 ;
        RECT 1760.175 208.285 1762.555 208.565 ;
        RECT 1763.395 208.285 1765.775 208.565 ;
        RECT 1766.615 208.285 1768.535 208.565 ;
        RECT 1769.375 208.285 1771.755 208.565 ;
        RECT 1772.595 208.285 1774.975 208.565 ;
        RECT 1775.815 208.285 1777.735 208.565 ;
        RECT 1778.575 208.285 1780.955 208.565 ;
        RECT 1781.795 208.285 1784.175 208.565 ;
        RECT 1785.015 208.285 1786.935 208.565 ;
        RECT 1787.775 208.285 1790.155 208.565 ;
        RECT 1790.995 208.285 1793.375 208.565 ;
        RECT 1794.215 208.285 1796.595 208.565 ;
        RECT 1797.435 208.285 1799.355 208.565 ;
        RECT 1800.195 208.285 1802.575 208.565 ;
        RECT 1803.415 208.285 1805.795 208.565 ;
        RECT 1806.635 208.285 1808.555 208.565 ;
        RECT 1809.395 208.285 1811.775 208.565 ;
        RECT 1812.615 208.285 1814.995 208.565 ;
        RECT 1815.835 208.285 1817.755 208.565 ;
        RECT 1818.595 208.285 1820.975 208.565 ;
        RECT 1821.815 208.285 1824.195 208.565 ;
        RECT 1825.035 208.285 1826.955 208.565 ;
        RECT 1827.795 208.285 1828.790 208.565 ;
        RECT 1749.085 0.000 1828.790 208.285 ;
        RECT 2023.085 208.285 2024.135 208.565 ;
        RECT 2024.975 208.285 2027.355 208.565 ;
        RECT 2028.195 208.285 2030.575 208.565 ;
        RECT 2031.415 208.285 2033.335 208.565 ;
        RECT 2034.175 208.285 2036.555 208.565 ;
        RECT 2037.395 208.285 2039.775 208.565 ;
        RECT 2040.615 208.285 2042.535 208.565 ;
        RECT 2043.375 208.285 2045.755 208.565 ;
        RECT 2046.595 208.285 2048.975 208.565 ;
        RECT 2049.815 208.285 2051.735 208.565 ;
        RECT 2052.575 208.285 2054.955 208.565 ;
        RECT 2055.795 208.285 2058.175 208.565 ;
        RECT 2059.015 208.285 2060.935 208.565 ;
        RECT 2061.775 208.285 2064.155 208.565 ;
        RECT 2064.995 208.285 2067.375 208.565 ;
        RECT 2068.215 208.285 2070.595 208.565 ;
        RECT 2071.435 208.285 2073.355 208.565 ;
        RECT 2074.195 208.285 2076.575 208.565 ;
        RECT 2077.415 208.285 2079.795 208.565 ;
        RECT 2080.635 208.285 2082.555 208.565 ;
        RECT 2083.395 208.285 2085.775 208.565 ;
        RECT 2086.615 208.285 2088.995 208.565 ;
        RECT 2089.835 208.285 2091.755 208.565 ;
        RECT 2092.595 208.285 2094.975 208.565 ;
        RECT 2095.815 208.285 2098.195 208.565 ;
        RECT 2099.035 208.285 2100.955 208.565 ;
        RECT 2101.795 208.285 2102.790 208.565 ;
        RECT 2023.085 0.000 2102.790 208.285 ;
        RECT 2297.085 208.285 2298.135 208.565 ;
        RECT 2298.975 208.285 2301.355 208.565 ;
        RECT 2302.195 208.285 2304.575 208.565 ;
        RECT 2305.415 208.285 2307.335 208.565 ;
        RECT 2308.175 208.285 2310.555 208.565 ;
        RECT 2311.395 208.285 2313.775 208.565 ;
        RECT 2314.615 208.285 2316.535 208.565 ;
        RECT 2317.375 208.285 2319.755 208.565 ;
        RECT 2320.595 208.285 2322.975 208.565 ;
        RECT 2323.815 208.285 2325.735 208.565 ;
        RECT 2326.575 208.285 2328.955 208.565 ;
        RECT 2329.795 208.285 2332.175 208.565 ;
        RECT 2333.015 208.285 2334.935 208.565 ;
        RECT 2335.775 208.285 2338.155 208.565 ;
        RECT 2338.995 208.285 2341.375 208.565 ;
        RECT 2342.215 208.285 2344.595 208.565 ;
        RECT 2345.435 208.285 2347.355 208.565 ;
        RECT 2348.195 208.285 2350.575 208.565 ;
        RECT 2351.415 208.285 2353.795 208.565 ;
        RECT 2354.635 208.285 2356.555 208.565 ;
        RECT 2357.395 208.285 2359.775 208.565 ;
        RECT 2360.615 208.285 2362.995 208.565 ;
        RECT 2363.835 208.285 2365.755 208.565 ;
        RECT 2366.595 208.285 2368.975 208.565 ;
        RECT 2369.815 208.285 2372.195 208.565 ;
        RECT 2373.035 208.285 2374.955 208.565 ;
        RECT 2375.795 208.285 2376.790 208.565 ;
        RECT 2297.085 0.000 2376.790 208.285 ;
        RECT 2571.085 208.285 2572.135 208.565 ;
        RECT 2572.975 208.285 2575.355 208.565 ;
        RECT 2576.195 208.285 2578.575 208.565 ;
        RECT 2579.415 208.285 2581.335 208.565 ;
        RECT 2582.175 208.285 2584.555 208.565 ;
        RECT 2585.395 208.285 2587.775 208.565 ;
        RECT 2588.615 208.285 2590.535 208.565 ;
        RECT 2591.375 208.285 2593.755 208.565 ;
        RECT 2594.595 208.285 2596.975 208.565 ;
        RECT 2597.815 208.285 2599.735 208.565 ;
        RECT 2600.575 208.285 2602.955 208.565 ;
        RECT 2603.795 208.285 2606.175 208.565 ;
        RECT 2607.015 208.285 2608.935 208.565 ;
        RECT 2609.775 208.285 2612.155 208.565 ;
        RECT 2612.995 208.285 2615.375 208.565 ;
        RECT 2616.215 208.285 2618.595 208.565 ;
        RECT 2619.435 208.285 2621.355 208.565 ;
        RECT 2622.195 208.285 2624.575 208.565 ;
        RECT 2625.415 208.285 2627.795 208.565 ;
        RECT 2628.635 208.285 2630.555 208.565 ;
        RECT 2631.395 208.285 2633.775 208.565 ;
        RECT 2634.615 208.285 2636.995 208.565 ;
        RECT 2637.835 208.285 2639.755 208.565 ;
        RECT 2640.595 208.285 2642.975 208.565 ;
        RECT 2643.815 208.285 2646.195 208.565 ;
        RECT 2647.035 208.285 2648.955 208.565 ;
        RECT 2649.795 208.285 2650.790 208.565 ;
        RECT 2571.085 0.000 2650.790 208.285 ;
        RECT 2845.710 197.965 2869.610 200.000 ;
        RECT 2892.105 198.080 2894.105 200.000 ;
        RECT 2895.605 197.965 2919.505 200.000 ;
        RECT 3114.710 197.965 3138.610 200.000 ;
        RECT 3161.105 198.080 3163.105 200.000 ;
        RECT 3164.605 197.965 3188.505 200.000 ;
        RECT 2845.710 4.925 2919.735 197.965 ;
        RECT 3114.710 4.925 3188.735 197.965 ;
      LAYER via2 ;
        RECT 212.140 561.855 212.550 563.670 ;
        RECT 211.080 347.205 211.445 349.835 ;
        RECT 2856.730 213.005 2858.685 214.805 ;
        RECT 454.360 210.915 455.425 211.195 ;
        RECT 717.145 201.320 717.425 201.600 ;
        RECT 1268.110 209.810 1269.075 210.170 ;
      LAYER met3 ;
        RECT 386.455 5070.750 460.250 5161.315 ;
        RECT 386.455 5002.905 410.320 5070.750 ;
        RECT 436.120 5002.905 460.250 5070.750 ;
        RECT 643.455 5070.750 717.250 5161.315 ;
        RECT 643.455 5002.905 667.320 5070.750 ;
        RECT 693.120 5002.905 717.250 5070.750 ;
        RECT 900.455 5070.750 974.250 5161.315 ;
        RECT 900.455 5002.905 924.320 5070.750 ;
        RECT 950.120 5002.905 974.250 5070.750 ;
        RECT 1105.000 5004.085 1274.000 5188.000 ;
        RECT 1368.000 5004.085 1537.000 5188.000 ;
        RECT 1667.240 5014.250 1741.290 5188.000 ;
      LAYER met3 ;
        RECT 1105.000 4988.000 1176.395 5003.685 ;
      LAYER met3 ;
        RECT 1176.795 4999.730 1201.990 5004.085 ;
        RECT 1176.795 4991.125 1189.490 4999.730 ;
        RECT 1176.795 4990.725 1177.495 4991.125 ;
        RECT 1189.295 4990.725 1189.490 4991.125 ;
      LAYER met3 ;
        RECT 1177.895 4988.000 1188.895 4990.725 ;
        RECT 1189.890 4988.000 1200.890 4999.330 ;
      LAYER met3 ;
        RECT 1201.290 4990.725 1201.990 4999.730 ;
      LAYER met3 ;
        RECT 1368.000 4988.000 1439.395 5003.685 ;
      LAYER met3 ;
        RECT 1439.795 4999.730 1464.990 5004.085 ;
        RECT 1439.795 4991.125 1452.490 4999.730 ;
        RECT 1439.795 4990.725 1440.495 4991.125 ;
        RECT 1452.295 4990.725 1452.490 4991.125 ;
      LAYER met3 ;
        RECT 1440.895 4988.000 1451.895 4990.725 ;
        RECT 1452.890 4988.000 1463.890 4999.330 ;
      LAYER met3 ;
        RECT 1464.290 4990.725 1464.990 4999.730 ;
      LAYER met3 ;
        RECT 1667.495 4988.000 1691.395 5013.850 ;
      LAYER met3 ;
        RECT 1691.795 4990.035 1716.990 5014.250 ;
        RECT 1692.895 4988.000 1703.895 4990.035 ;
        RECT 1704.890 4988.000 1715.890 4990.035 ;
      LAYER met3 ;
        RECT 1717.390 4988.000 1741.290 5013.850 ;
      LAYER met3 ;
        RECT 1877.000 5004.085 2046.000 5188.000 ;
        RECT 2369.455 5070.750 2443.250 5161.315 ;
      LAYER met3 ;
        RECT 1877.000 4988.000 1948.395 5003.685 ;
      LAYER met3 ;
        RECT 1948.795 4999.730 1973.990 5004.085 ;
        RECT 2369.455 5002.905 2393.320 5070.750 ;
        RECT 2419.120 5002.905 2443.250 5070.750 ;
        RECT 2626.455 5070.750 2700.250 5161.315 ;
        RECT 2626.455 5002.905 2650.320 5070.750 ;
        RECT 2676.120 5002.905 2700.250 5070.750 ;
        RECT 2878.240 5025.160 2952.290 5183.100 ;
        RECT 3135.455 5070.750 3209.250 5161.315 ;
        RECT 2878.240 5020.915 2927.990 5025.160 ;
        RECT 1948.795 4991.125 1961.490 4999.730 ;
        RECT 1948.795 4990.725 1949.495 4991.125 ;
        RECT 1961.295 4990.725 1961.490 4991.125 ;
      LAYER met3 ;
        RECT 1949.895 4988.000 1960.895 4990.725 ;
        RECT 1961.890 4988.000 1972.890 4999.330 ;
      LAYER met3 ;
        RECT 1973.290 4990.725 1973.990 4999.730 ;
      LAYER met3 ;
        RECT 2878.495 4988.000 2902.395 5020.515 ;
      LAYER met3 ;
        RECT 2902.795 4990.035 2927.990 5020.915 ;
        RECT 2903.895 4988.000 2914.895 4990.035 ;
        RECT 2915.890 4988.000 2926.890 4990.035 ;
      LAYER met3 ;
        RECT 2928.390 4988.000 2952.290 5024.760 ;
      LAYER met3 ;
        RECT 3135.455 5002.905 3159.320 5070.750 ;
        RECT 3185.120 5002.905 3209.250 5070.750 ;
        RECT 26.685 4826.120 185.095 4850.250 ;
        RECT 26.685 4800.320 117.250 4826.120 ;
        RECT 3402.905 4808.680 3561.315 4832.545 ;
        RECT 26.685 4776.455 185.095 4800.320 ;
        RECT 3470.750 4782.880 3561.315 4808.680 ;
        RECT 3402.905 4758.750 3561.315 4782.880 ;
        RECT 0.000 4398.990 179.800 4423.290 ;
      LAYER met3 ;
        RECT 180.200 4399.390 200.000 4423.290 ;
      LAYER met3 ;
        RECT 0.000 4397.890 197.965 4398.990 ;
        RECT 0.000 4386.890 200.000 4397.890 ;
        RECT 0.000 4385.895 197.965 4386.890 ;
        RECT 0.000 4374.895 200.000 4385.895 ;
        RECT 0.000 4373.795 197.965 4374.895 ;
        RECT 0.000 4349.240 179.800 4373.795 ;
      LAYER met3 ;
        RECT 180.200 4349.495 200.000 4373.395 ;
      LAYER met3 ;
        RECT 3386.690 4312.430 3588.000 4391.690 ;
        RECT 4.900 4187.990 162.840 4212.290 ;
      LAYER met3 ;
        RECT 163.240 4188.390 200.000 4212.290 ;
      LAYER met3 ;
        RECT 4.900 4186.890 197.965 4187.990 ;
        RECT 4.900 4175.890 200.000 4186.890 ;
        RECT 4.900 4174.895 197.965 4175.890 ;
        RECT 4.900 4163.895 200.000 4174.895 ;
        RECT 4.900 4162.795 197.965 4163.895 ;
        RECT 4.900 4138.240 167.085 4162.795 ;
      LAYER met3 ;
        RECT 167.485 4138.495 200.000 4162.395 ;
        RECT 3388.000 4142.605 3402.960 4166.505 ;
      LAYER met3 ;
        RECT 3403.360 4142.205 3588.000 4166.760 ;
        RECT 3390.035 4141.105 3588.000 4142.205 ;
        RECT 3388.000 4130.105 3588.000 4141.105 ;
        RECT 3390.035 4129.110 3588.000 4130.105 ;
        RECT 3388.000 4118.110 3588.000 4129.110 ;
        RECT 3390.035 4117.010 3588.000 4118.110 ;
      LAYER met3 ;
        RECT 3388.000 4092.710 3402.960 4116.610 ;
      LAYER met3 ;
        RECT 3403.360 4092.710 3588.000 4117.010 ;
        RECT 0.000 3922.310 201.310 4001.570 ;
        RECT 3386.690 3866.430 3588.000 3945.690 ;
        RECT 0.000 3706.310 201.310 3785.570 ;
        RECT 3386.690 3641.430 3588.000 3720.690 ;
        RECT 0.000 3490.310 201.310 3569.570 ;
        RECT 3386.690 3416.430 3588.000 3495.690 ;
        RECT 0.000 3274.310 201.310 3353.570 ;
        RECT 3386.690 3190.430 3588.000 3269.690 ;
        RECT 0.000 3058.310 201.310 3137.570 ;
        RECT 3386.690 2965.430 3588.000 3044.690 ;
        RECT 0.000 2842.310 201.310 2921.570 ;
        RECT 3386.690 2739.430 3588.000 2818.690 ;
        RECT 0.000 2626.310 201.310 2705.570 ;
      LAYER met3 ;
        RECT 3388.000 2569.605 3402.960 2593.505 ;
      LAYER met3 ;
        RECT 3403.360 2569.205 3588.000 2593.760 ;
        RECT 3390.035 2568.105 3588.000 2569.205 ;
        RECT 3388.000 2557.105 3588.000 2568.105 ;
        RECT 3390.035 2556.110 3588.000 2557.105 ;
        RECT 3388.000 2545.110 3588.000 2556.110 ;
        RECT 3390.035 2544.010 3588.000 2545.110 ;
      LAYER met3 ;
        RECT 3388.000 2519.710 3402.960 2543.610 ;
      LAYER met3 ;
        RECT 3403.360 2519.710 3588.000 2544.010 ;
        RECT 0.000 2464.990 184.640 2489.290 ;
      LAYER met3 ;
        RECT 185.040 2465.390 200.000 2489.290 ;
      LAYER met3 ;
        RECT 0.000 2463.890 197.965 2464.990 ;
        RECT 0.000 2452.890 200.000 2463.890 ;
        RECT 0.000 2451.895 197.965 2452.890 ;
        RECT 0.000 2440.895 200.000 2451.895 ;
        RECT 0.000 2439.795 197.965 2440.895 ;
        RECT 0.000 2415.240 184.640 2439.795 ;
      LAYER met3 ;
        RECT 185.040 2415.495 200.000 2439.395 ;
        RECT 3390.000 2349.500 3416.435 2373.500 ;
        RECT 171.165 2204.500 198.000 2228.500 ;
        RECT 3388.000 2128.605 3420.515 2152.505 ;
      LAYER met3 ;
        RECT 3420.915 2128.205 3583.100 2152.760 ;
        RECT 3390.035 2127.105 3583.100 2128.205 ;
        RECT 3388.000 2116.105 3583.100 2127.105 ;
        RECT 3390.035 2115.110 3583.100 2116.105 ;
        RECT 3388.000 2104.110 3583.100 2115.110 ;
        RECT 3390.035 2103.010 3583.100 2104.110 ;
      LAYER met3 ;
        RECT 3388.000 2078.710 3424.760 2102.610 ;
      LAYER met3 ;
        RECT 3425.160 2078.710 3583.100 2103.010 ;
        RECT 0.000 1988.310 201.310 2067.570 ;
        RECT 3386.690 1853.430 3588.000 1932.690 ;
        RECT 0.000 1772.310 201.310 1851.570 ;
        RECT 0.000 1556.310 201.310 1635.570 ;
        RECT 3386.690 1627.430 3588.000 1706.690 ;
        RECT 0.000 1340.310 201.310 1419.570 ;
        RECT 3386.690 1402.430 3588.000 1481.690 ;
        RECT 0.000 1124.310 201.310 1203.570 ;
        RECT 3386.690 1177.430 3588.000 1256.690 ;
        RECT 0.000 908.310 201.310 987.570 ;
        RECT 3386.690 951.430 3588.000 1030.690 ;
        RECT 3386.690 726.430 3588.000 805.690 ;
        RECT 0.000 600.990 179.800 625.290 ;
      LAYER met3 ;
        RECT 180.200 601.390 200.000 625.290 ;
      LAYER met3 ;
        RECT 0.000 599.890 197.965 600.990 ;
        RECT 0.000 588.890 200.000 599.890 ;
        RECT 0.000 587.895 197.965 588.890 ;
        RECT 0.000 576.895 200.000 587.895 ;
        RECT 0.000 575.795 197.965 576.895 ;
        RECT 0.000 551.240 179.800 575.795 ;
      LAYER met3 ;
        RECT 180.200 563.625 200.000 575.395 ;
        RECT 212.070 563.625 212.595 563.775 ;
        RECT 180.200 561.900 212.595 563.625 ;
        RECT 180.200 551.495 200.000 561.900 ;
        RECT 212.070 561.770 212.595 561.900 ;
      LAYER met3 ;
        RECT 3386.690 500.430 3588.000 579.690 ;
        RECT 153.765 415.605 158.415 426.140 ;
        RECT 159.805 415.440 163.270 426.140 ;
        RECT 4.395 390.355 190.700 415.000 ;
      LAYER met3 ;
        RECT 191.100 390.755 198.000 414.700 ;
      LAYER met3 ;
        RECT 4.395 389.255 197.965 390.355 ;
        RECT 4.395 378.380 198.000 389.255 ;
        RECT 4.395 376.880 197.965 378.380 ;
        RECT 4.395 366.000 198.000 376.880 ;
        RECT 4.395 364.900 197.965 366.000 ;
        RECT 4.395 340.490 190.700 364.900 ;
      LAYER met3 ;
        RECT 191.100 349.830 198.000 364.500 ;
        RECT 211.050 349.830 211.480 349.935 ;
        RECT 191.100 347.205 211.480 349.830 ;
        RECT 191.100 340.500 198.000 347.205 ;
        RECT 211.050 347.125 211.480 347.205 ;
        RECT 2856.605 212.915 2858.820 214.920 ;
        RECT 454.330 211.225 455.460 211.920 ;
        RECT 454.315 210.870 455.470 211.225 ;
        RECT 454.330 200.000 455.460 210.870 ;
        RECT 717.120 200.000 717.450 201.625 ;
        RECT 238.000 164.765 256.010 180.085 ;
        RECT 258.000 164.765 276.010 180.085 ;
        RECT 278.000 164.765 296.010 180.085 ;
        RECT 298.000 164.765 316.010 180.085 ;
        RECT 318.000 164.765 336.010 180.085 ;
        RECT 338.000 164.765 356.010 180.085 ;
        RECT 394.710 163.240 418.610 200.000 ;
      LAYER met3 ;
        RECT 420.110 197.965 431.110 200.000 ;
        RECT 432.105 197.965 443.105 200.000 ;
        RECT 419.010 167.085 444.205 197.965 ;
      LAYER met3 ;
        RECT 444.605 167.485 468.505 200.000 ;
      LAYER met3 ;
        RECT 419.010 162.840 468.760 167.085 ;
      LAYER met3 ;
        RECT 507.000 164.765 525.010 180.085 ;
        RECT 527.000 164.765 545.010 180.085 ;
        RECT 547.000 164.765 565.010 180.085 ;
        RECT 567.000 164.765 585.010 180.085 ;
        RECT 587.000 164.765 605.010 180.085 ;
        RECT 607.000 164.765 625.010 180.085 ;
      LAYER met3 ;
        RECT 394.710 4.900 468.760 162.840 ;
        RECT 663.300 151.080 664.340 199.375 ;
        RECT 663.300 133.400 663.675 151.080 ;
      LAYER met3 ;
        RECT 664.740 150.680 665.810 200.000 ;
        RECT 664.075 135.400 665.810 150.680 ;
      LAYER met3 ;
        RECT 666.210 188.690 707.935 199.375 ;
      LAYER met3 ;
        RECT 708.335 190.155 709.065 200.000 ;
      LAYER met3 ;
        RECT 709.465 193.730 716.375 199.375 ;
        RECT 709.465 192.265 714.910 193.730 ;
      LAYER met3 ;
        RECT 716.775 193.330 717.925 200.000 ;
      LAYER met3 ;
        RECT 709.465 191.985 714.630 192.265 ;
        RECT 709.465 190.555 713.550 191.985 ;
      LAYER met3 ;
        RECT 715.310 191.950 717.925 193.330 ;
        RECT 715.310 191.865 716.875 191.950 ;
        RECT 716.940 191.865 717.925 191.950 ;
      LAYER met3 ;
        RECT 718.325 196.465 718.690 199.375 ;
      LAYER met3 ;
        RECT 719.090 196.865 720.755 200.000 ;
      LAYER met3 ;
        RECT 721.155 196.465 728.680 199.375 ;
      LAYER met3 ;
        RECT 715.030 191.800 715.310 191.865 ;
        RECT 715.395 191.800 716.940 191.865 ;
        RECT 715.030 191.650 716.940 191.800 ;
        RECT 715.030 191.585 716.575 191.650 ;
        RECT 716.660 191.585 716.940 191.650 ;
      LAYER met3 ;
        RECT 709.765 190.255 713.550 190.555 ;
      LAYER met3 ;
        RECT 708.335 189.855 709.365 190.155 ;
        RECT 708.335 189.555 709.100 189.855 ;
        RECT 709.365 189.555 709.830 189.855 ;
        RECT 708.335 189.090 709.830 189.555 ;
      LAYER met3 ;
        RECT 666.210 184.830 708.700 188.690 ;
      LAYER met3 ;
        RECT 709.100 185.230 709.830 189.090 ;
      LAYER met3 ;
        RECT 710.230 187.335 713.550 190.255 ;
      LAYER met3 ;
        RECT 713.950 191.500 715.030 191.585 ;
        RECT 715.095 191.500 716.660 191.585 ;
        RECT 713.950 190.020 716.660 191.500 ;
      LAYER met3 ;
        RECT 718.325 191.465 728.680 196.465 ;
        RECT 717.340 191.185 728.680 191.465 ;
      LAYER met3 ;
        RECT 713.950 187.735 715.095 190.020 ;
      LAYER met3 ;
        RECT 717.060 189.620 728.680 191.185 ;
        RECT 715.495 187.335 728.680 189.620 ;
        RECT 710.230 184.830 728.680 187.335 ;
        RECT 666.210 183.015 728.680 184.830 ;
      LAYER met3 ;
        RECT 729.080 184.215 729.600 200.280 ;
      LAYER met3 ;
        RECT 730.000 184.615 737.035 199.375 ;
        RECT 730.210 184.405 737.035 184.615 ;
      LAYER met3 ;
        RECT 729.080 184.005 729.810 184.215 ;
        RECT 729.080 183.555 730.260 184.005 ;
      LAYER met3 ;
        RECT 730.660 183.955 737.035 184.405 ;
      LAYER met3 ;
        RECT 729.080 183.415 729.670 183.555 ;
        RECT 729.680 183.415 730.710 183.555 ;
      LAYER met3 ;
        RECT 731.110 183.505 737.035 183.955 ;
      LAYER met3 ;
        RECT 729.670 183.105 730.710 183.415 ;
      LAYER met3 ;
        RECT 666.210 182.555 729.270 183.015 ;
      LAYER met3 ;
        RECT 729.670 182.955 731.225 183.105 ;
      LAYER met3 ;
        RECT 666.210 181.980 729.730 182.555 ;
      LAYER met3 ;
        RECT 730.130 182.380 731.225 182.955 ;
      LAYER met3 ;
        RECT 666.210 169.105 730.305 181.980 ;
        RECT 666.210 168.520 729.720 169.105 ;
      LAYER met3 ;
        RECT 730.705 168.705 731.225 182.380 ;
      LAYER met3 ;
        RECT 666.210 167.805 729.005 168.520 ;
      LAYER met3 ;
        RECT 730.120 168.195 731.225 168.705 ;
        RECT 730.120 168.120 730.775 168.195 ;
        RECT 730.850 168.120 731.225 168.195 ;
        RECT 729.405 168.045 730.120 168.120 ;
        RECT 730.135 168.045 730.850 168.120 ;
      LAYER met3 ;
        RECT 666.210 167.220 728.420 167.805 ;
      LAYER met3 ;
        RECT 729.405 167.445 730.850 168.045 ;
      LAYER met3 ;
        RECT 731.625 167.720 737.035 183.505 ;
      LAYER met3 ;
        RECT 729.405 167.405 730.120 167.445 ;
        RECT 730.135 167.405 730.850 167.445 ;
        RECT 728.820 167.295 729.405 167.405 ;
        RECT 729.445 167.295 730.135 167.405 ;
      LAYER met3 ;
        RECT 666.210 167.005 728.205 167.220 ;
        RECT 666.210 165.475 715.325 167.005 ;
      LAYER met3 ;
        RECT 728.820 166.845 730.135 167.295 ;
      LAYER met3 ;
        RECT 731.250 167.005 737.035 167.720 ;
      LAYER met3 ;
        RECT 728.820 166.820 729.425 166.845 ;
        RECT 729.550 166.820 730.135 166.845 ;
        RECT 728.605 166.695 728.820 166.820 ;
        RECT 728.845 166.695 729.550 166.820 ;
        RECT 728.605 166.605 729.550 166.695 ;
        RECT 715.725 166.305 729.550 166.605 ;
      LAYER met3 ;
        RECT 730.535 166.420 737.035 167.005 ;
      LAYER met3 ;
        RECT 715.725 166.300 728.885 166.305 ;
        RECT 729.030 166.300 729.550 166.305 ;
        RECT 715.725 165.875 729.030 166.300 ;
      LAYER met3 ;
        RECT 729.950 165.900 737.035 166.420 ;
        RECT 729.430 165.475 737.035 165.900 ;
        RECT 666.210 135.800 737.035 165.475 ;
      LAYER met3 ;
        RECT 776.000 164.765 794.010 180.085 ;
        RECT 796.000 164.765 814.010 180.085 ;
        RECT 816.000 164.765 834.010 180.085 ;
        RECT 836.000 164.765 854.010 180.085 ;
        RECT 856.000 164.765 874.010 180.085 ;
        RECT 876.000 164.765 894.010 180.085 ;
        RECT 664.075 133.800 667.410 135.400 ;
      LAYER met3 ;
        RECT 667.810 134.200 737.035 135.800 ;
        RECT 663.300 131.800 665.410 133.400 ;
      LAYER met3 ;
        RECT 665.810 132.400 668.810 133.800 ;
      LAYER met3 ;
        RECT 669.210 132.800 737.035 134.200 ;
      LAYER met3 ;
        RECT 665.810 132.250 669.745 132.400 ;
        RECT 665.810 132.200 667.410 132.250 ;
        RECT 667.510 132.200 669.745 132.250 ;
      LAYER met3 ;
        RECT 663.300 130.515 667.010 131.800 ;
      LAYER met3 ;
        RECT 667.410 131.465 669.745 132.200 ;
      LAYER met3 ;
        RECT 670.145 131.865 737.035 132.800 ;
      LAYER met3 ;
        RECT 667.410 131.350 669.710 131.465 ;
        RECT 669.745 131.350 670.610 131.465 ;
        RECT 667.410 131.050 670.610 131.350 ;
        RECT 667.410 130.915 668.695 131.050 ;
        RECT 668.710 130.915 670.610 131.050 ;
      LAYER met3 ;
        RECT 671.010 131.000 737.035 131.865 ;
      LAYER met3 ;
        RECT 668.695 130.600 670.610 130.915 ;
      LAYER met3 ;
        RECT 663.300 129.565 668.295 130.515 ;
      LAYER met3 ;
        RECT 668.695 130.000 671.960 130.600 ;
        RECT 668.695 129.965 669.645 130.000 ;
        RECT 669.760 129.965 671.960 130.000 ;
      LAYER met3 ;
        RECT 663.300 128.600 669.245 129.565 ;
      LAYER met3 ;
        RECT 669.645 129.250 671.960 129.965 ;
      LAYER met3 ;
        RECT 672.360 129.650 737.035 131.000 ;
      LAYER met3 ;
        RECT 669.645 129.100 673.140 129.250 ;
        RECT 669.645 129.000 670.610 129.100 ;
        RECT 670.660 129.000 673.140 129.100 ;
      LAYER met3 ;
        RECT 663.300 127.390 670.210 128.600 ;
      LAYER met3 ;
        RECT 670.610 127.920 673.140 129.000 ;
        RECT 670.610 127.790 671.820 127.920 ;
        RECT 671.840 127.790 673.140 127.920 ;
        RECT 671.820 127.600 673.140 127.790 ;
      LAYER met3 ;
        RECT 663.300 127.200 671.420 127.390 ;
        RECT 663.300 104.955 671.610 127.200 ;
      LAYER met3 ;
        RECT 672.010 105.355 673.140 127.600 ;
      LAYER met3 ;
        RECT 673.540 104.955 737.035 129.650 ;
        RECT 663.300 0.000 737.035 104.955 ;
        RECT 932.430 0.000 1011.690 201.310 ;
      LAYER met3 ;
        RECT 1268.065 198.000 1269.135 210.215 ;
        RECT 1050.000 164.765 1068.010 180.085 ;
        RECT 1070.000 164.765 1088.010 180.085 ;
        RECT 1090.000 164.765 1108.010 180.085 ;
        RECT 1110.000 164.765 1128.010 180.085 ;
        RECT 1130.000 164.765 1148.010 180.085 ;
        RECT 1150.000 164.765 1168.010 180.085 ;
      LAYER met3 ;
        RECT 1194.860 159.805 1205.560 163.270 ;
        RECT 1194.860 153.765 1205.395 158.415 ;
      LAYER met3 ;
        RECT 1206.300 158.400 1230.245 198.000 ;
      LAYER met3 ;
        RECT 1231.745 197.965 1242.620 198.000 ;
        RECT 1244.120 197.965 1255.000 198.000 ;
        RECT 1230.645 158.000 1256.100 197.965 ;
      LAYER met3 ;
        RECT 1256.500 158.400 1280.500 198.000 ;
        RECT 1319.000 164.765 1337.010 180.085 ;
        RECT 1339.000 164.765 1357.010 180.085 ;
        RECT 1359.000 164.765 1377.010 180.085 ;
        RECT 1379.000 164.765 1397.010 180.085 ;
        RECT 1399.000 164.765 1417.010 180.085 ;
        RECT 1419.000 164.765 1437.010 180.085 ;
      LAYER met3 ;
        RECT 1206.000 4.395 1280.500 158.000 ;
        RECT 1475.430 0.000 1554.690 201.310 ;
      LAYER met3 ;
        RECT 1593.000 164.765 1611.010 180.085 ;
        RECT 1613.000 164.765 1631.010 180.085 ;
        RECT 1633.000 164.765 1651.010 180.085 ;
        RECT 1653.000 164.765 1671.010 180.085 ;
        RECT 1673.000 164.765 1691.010 180.085 ;
        RECT 1693.000 164.765 1711.010 180.085 ;
      LAYER met3 ;
        RECT 1749.430 0.000 1828.690 201.310 ;
      LAYER met3 ;
        RECT 1867.000 164.765 1885.010 180.085 ;
        RECT 1887.000 164.765 1905.010 180.085 ;
        RECT 1907.000 164.765 1925.010 180.085 ;
        RECT 1927.000 164.765 1945.010 180.085 ;
        RECT 1947.000 164.765 1965.010 180.085 ;
        RECT 1967.000 164.765 1985.010 180.085 ;
      LAYER met3 ;
        RECT 2023.430 0.000 2102.690 201.310 ;
      LAYER met3 ;
        RECT 2141.000 164.765 2159.010 180.085 ;
        RECT 2161.000 164.765 2179.010 180.085 ;
        RECT 2181.000 164.765 2199.010 180.085 ;
        RECT 2201.000 164.765 2219.010 180.085 ;
        RECT 2221.000 164.765 2239.010 180.085 ;
        RECT 2241.000 164.765 2259.010 180.085 ;
      LAYER met3 ;
        RECT 2297.430 0.000 2376.690 201.310 ;
      LAYER met3 ;
        RECT 2415.000 164.765 2433.010 180.085 ;
        RECT 2435.000 164.765 2453.010 180.085 ;
        RECT 2455.000 164.765 2473.010 180.085 ;
        RECT 2475.000 164.765 2493.010 180.085 ;
        RECT 2495.000 164.765 2513.010 180.085 ;
        RECT 2515.000 164.765 2533.010 180.085 ;
      LAYER met3 ;
        RECT 2571.430 0.000 2650.690 201.310 ;
      LAYER met3 ;
        RECT 2856.965 200.000 2858.460 212.915 ;
        RECT 2689.000 164.765 2707.010 180.085 ;
        RECT 2709.000 164.765 2727.010 180.085 ;
        RECT 2729.000 164.765 2747.010 180.085 ;
        RECT 2749.000 164.765 2767.010 180.085 ;
        RECT 2769.000 164.765 2787.010 180.085 ;
        RECT 2789.000 164.765 2807.010 180.085 ;
        RECT 2845.710 174.150 2869.610 200.000 ;
      LAYER met3 ;
        RECT 2871.110 197.965 2882.110 200.000 ;
        RECT 2883.105 197.965 2894.105 200.000 ;
        RECT 2870.010 173.750 2895.205 197.965 ;
      LAYER met3 ;
        RECT 2895.605 174.150 2919.505 200.000 ;
        RECT 3114.710 185.040 3138.610 200.000 ;
      LAYER met3 ;
        RECT 3140.110 197.965 3151.110 200.000 ;
        RECT 3152.105 197.965 3163.105 200.000 ;
        RECT 3139.010 184.640 3164.205 197.965 ;
      LAYER met3 ;
        RECT 3164.605 185.040 3188.505 200.000 ;
      LAYER met3 ;
        RECT 2845.710 0.000 2919.760 173.750 ;
      LAYER met3 ;
        RECT 2958.000 164.765 2976.010 180.085 ;
        RECT 2978.000 164.765 2996.010 180.085 ;
        RECT 2998.000 164.765 3016.010 180.085 ;
        RECT 3018.000 164.765 3036.010 180.085 ;
        RECT 3038.000 164.765 3056.010 180.085 ;
        RECT 3058.000 164.765 3076.010 180.085 ;
      LAYER met3 ;
        RECT 3114.710 0.000 3188.760 184.640 ;
      LAYER met3 ;
        RECT 3227.000 164.765 3245.010 180.085 ;
        RECT 3247.000 164.765 3265.010 180.085 ;
        RECT 3267.000 164.765 3285.010 180.085 ;
        RECT 3287.000 164.765 3305.010 180.085 ;
        RECT 3307.000 164.765 3325.010 180.085 ;
        RECT 3327.000 164.765 3345.010 180.085 ;
      LAYER via3 ;
        RECT 238.230 175.875 255.720 179.885 ;
        RECT 238.260 164.935 255.910 167.885 ;
        RECT 258.230 175.875 275.720 179.885 ;
        RECT 258.260 164.935 275.910 167.885 ;
        RECT 278.230 175.875 295.720 179.885 ;
        RECT 278.260 164.935 295.910 167.885 ;
        RECT 298.230 175.875 315.720 179.885 ;
        RECT 298.260 164.935 315.910 167.885 ;
        RECT 318.230 175.875 335.720 179.885 ;
        RECT 318.260 164.935 335.910 167.885 ;
        RECT 338.230 175.875 355.720 179.885 ;
        RECT 338.260 164.935 355.910 167.885 ;
        RECT 507.230 175.875 524.720 179.885 ;
        RECT 507.260 164.935 524.910 167.885 ;
        RECT 527.230 175.875 544.720 179.885 ;
        RECT 527.260 164.935 544.910 167.885 ;
        RECT 547.230 175.875 564.720 179.885 ;
        RECT 547.260 164.935 564.910 167.885 ;
        RECT 567.230 175.875 584.720 179.885 ;
        RECT 567.260 164.935 584.910 167.885 ;
        RECT 587.230 175.875 604.720 179.885 ;
        RECT 587.260 164.935 604.910 167.885 ;
        RECT 607.230 175.875 624.720 179.885 ;
        RECT 607.260 164.935 624.910 167.885 ;
        RECT 776.230 175.875 793.720 179.885 ;
        RECT 776.260 164.935 793.910 167.885 ;
        RECT 796.230 175.875 813.720 179.885 ;
        RECT 796.260 164.935 813.910 167.885 ;
        RECT 816.230 175.875 833.720 179.885 ;
        RECT 816.260 164.935 833.910 167.885 ;
        RECT 836.230 175.875 853.720 179.885 ;
        RECT 836.260 164.935 853.910 167.885 ;
        RECT 856.230 175.875 873.720 179.885 ;
        RECT 856.260 164.935 873.910 167.885 ;
        RECT 876.230 175.875 893.720 179.885 ;
        RECT 876.260 164.935 893.910 167.885 ;
        RECT 1050.230 175.875 1067.720 179.885 ;
        RECT 1050.260 164.935 1067.910 167.885 ;
        RECT 1070.230 175.875 1087.720 179.885 ;
        RECT 1070.260 164.935 1087.910 167.885 ;
        RECT 1090.230 175.875 1107.720 179.885 ;
        RECT 1090.260 164.935 1107.910 167.885 ;
        RECT 1110.230 175.875 1127.720 179.885 ;
        RECT 1110.260 164.935 1127.910 167.885 ;
        RECT 1130.230 175.875 1147.720 179.885 ;
        RECT 1130.260 164.935 1147.910 167.885 ;
        RECT 1150.230 175.875 1167.720 179.885 ;
        RECT 1150.260 164.935 1167.910 167.885 ;
        RECT 1319.230 175.875 1336.720 179.885 ;
        RECT 1319.260 164.935 1336.910 167.885 ;
        RECT 1339.230 175.875 1356.720 179.885 ;
        RECT 1339.260 164.935 1356.910 167.885 ;
        RECT 1359.230 175.875 1376.720 179.885 ;
        RECT 1359.260 164.935 1376.910 167.885 ;
        RECT 1379.230 175.875 1396.720 179.885 ;
        RECT 1379.260 164.935 1396.910 167.885 ;
        RECT 1399.230 175.875 1416.720 179.885 ;
        RECT 1399.260 164.935 1416.910 167.885 ;
        RECT 1419.230 175.875 1436.720 179.885 ;
        RECT 1419.260 164.935 1436.910 167.885 ;
        RECT 1593.230 175.875 1610.720 179.885 ;
        RECT 1593.260 164.935 1610.910 167.885 ;
        RECT 1613.230 175.875 1630.720 179.885 ;
        RECT 1613.260 164.935 1630.910 167.885 ;
        RECT 1633.230 175.875 1650.720 179.885 ;
        RECT 1633.260 164.935 1650.910 167.885 ;
        RECT 1653.230 175.875 1670.720 179.885 ;
        RECT 1653.260 164.935 1670.910 167.885 ;
        RECT 1673.230 175.875 1690.720 179.885 ;
        RECT 1673.260 164.935 1690.910 167.885 ;
        RECT 1693.230 175.875 1710.720 179.885 ;
        RECT 1693.260 164.935 1710.910 167.885 ;
        RECT 1867.230 175.875 1884.720 179.885 ;
        RECT 1867.260 164.935 1884.910 167.885 ;
        RECT 1887.230 175.875 1904.720 179.885 ;
        RECT 1887.260 164.935 1904.910 167.885 ;
        RECT 1907.230 175.875 1924.720 179.885 ;
        RECT 1907.260 164.935 1924.910 167.885 ;
        RECT 1927.230 175.875 1944.720 179.885 ;
        RECT 1927.260 164.935 1944.910 167.885 ;
        RECT 1947.230 175.875 1964.720 179.885 ;
        RECT 1947.260 164.935 1964.910 167.885 ;
        RECT 1967.230 175.875 1984.720 179.885 ;
        RECT 1967.260 164.935 1984.910 167.885 ;
        RECT 2141.230 175.875 2158.720 179.885 ;
        RECT 2141.260 164.935 2158.910 167.885 ;
        RECT 2161.230 175.875 2178.720 179.885 ;
        RECT 2161.260 164.935 2178.910 167.885 ;
        RECT 2181.230 175.875 2198.720 179.885 ;
        RECT 2181.260 164.935 2198.910 167.885 ;
        RECT 2201.230 175.875 2218.720 179.885 ;
        RECT 2201.260 164.935 2218.910 167.885 ;
        RECT 2221.230 175.875 2238.720 179.885 ;
        RECT 2221.260 164.935 2238.910 167.885 ;
        RECT 2241.230 175.875 2258.720 179.885 ;
        RECT 2241.260 164.935 2258.910 167.885 ;
        RECT 2415.230 175.875 2432.720 179.885 ;
        RECT 2415.260 164.935 2432.910 167.885 ;
        RECT 2435.230 175.875 2452.720 179.885 ;
        RECT 2435.260 164.935 2452.910 167.885 ;
        RECT 2455.230 175.875 2472.720 179.885 ;
        RECT 2455.260 164.935 2472.910 167.885 ;
        RECT 2475.230 175.875 2492.720 179.885 ;
        RECT 2475.260 164.935 2492.910 167.885 ;
        RECT 2495.230 175.875 2512.720 179.885 ;
        RECT 2495.260 164.935 2512.910 167.885 ;
        RECT 2515.230 175.875 2532.720 179.885 ;
        RECT 2515.260 164.935 2532.910 167.885 ;
        RECT 2689.230 175.875 2706.720 179.885 ;
        RECT 2689.260 164.935 2706.910 167.885 ;
        RECT 2709.230 175.875 2726.720 179.885 ;
        RECT 2709.260 164.935 2726.910 167.885 ;
        RECT 2729.230 175.875 2746.720 179.885 ;
        RECT 2729.260 164.935 2746.910 167.885 ;
        RECT 2749.230 175.875 2766.720 179.885 ;
        RECT 2749.260 164.935 2766.910 167.885 ;
        RECT 2769.230 175.875 2786.720 179.885 ;
        RECT 2769.260 164.935 2786.910 167.885 ;
        RECT 2789.230 175.875 2806.720 179.885 ;
        RECT 2958.230 175.875 2975.720 179.885 ;
        RECT 2789.260 164.935 2806.910 167.885 ;
        RECT 2958.260 164.935 2975.910 167.885 ;
        RECT 2978.230 175.875 2995.720 179.885 ;
        RECT 2978.260 164.935 2995.910 167.885 ;
        RECT 2998.230 175.875 3015.720 179.885 ;
        RECT 2998.260 164.935 3015.910 167.885 ;
        RECT 3018.230 175.875 3035.720 179.885 ;
        RECT 3018.260 164.935 3035.910 167.885 ;
        RECT 3038.230 175.875 3055.720 179.885 ;
        RECT 3038.260 164.935 3055.910 167.885 ;
        RECT 3058.230 175.875 3075.720 179.885 ;
        RECT 3058.260 164.935 3075.910 167.885 ;
        RECT 3227.230 175.875 3244.720 179.885 ;
        RECT 3227.260 164.935 3244.910 167.885 ;
        RECT 3247.230 175.875 3264.720 179.885 ;
        RECT 3247.260 164.935 3264.910 167.885 ;
        RECT 3267.230 175.875 3284.720 179.885 ;
        RECT 3267.260 164.935 3284.910 167.885 ;
        RECT 3287.230 175.875 3304.720 179.885 ;
        RECT 3287.260 164.935 3304.910 167.885 ;
        RECT 3307.230 175.875 3324.720 179.885 ;
        RECT 3307.260 164.935 3324.910 167.885 ;
        RECT 3327.230 175.875 3344.720 179.885 ;
        RECT 3327.260 164.935 3344.910 167.885 ;
      LAYER met4 ;
        RECT 0.000 5163.385 202.330 5188.000 ;
      LAYER met4 ;
        RECT 202.730 5163.785 204.000 5188.000 ;
      LAYER met4 ;
        RECT 0.000 5083.400 202.745 5163.385 ;
        RECT 204.000 5083.400 386.000 5188.000 ;
      LAYER met4 ;
        RECT 386.000 5163.785 387.270 5188.000 ;
      LAYER met4 ;
        RECT 387.670 5163.385 459.330 5188.000 ;
      LAYER met4 ;
        RECT 459.730 5163.785 461.000 5188.000 ;
      LAYER met4 ;
        RECT 386.965 5083.400 460.035 5163.385 ;
        RECT 461.000 5083.400 643.000 5188.000 ;
      LAYER met4 ;
        RECT 643.000 5163.785 644.270 5188.000 ;
      LAYER met4 ;
        RECT 644.670 5163.385 716.330 5188.000 ;
      LAYER met4 ;
        RECT 716.730 5163.785 718.000 5188.000 ;
      LAYER met4 ;
        RECT 643.965 5083.400 717.035 5163.385 ;
        RECT 718.000 5083.400 900.000 5188.000 ;
      LAYER met4 ;
        RECT 900.000 5163.785 901.270 5188.000 ;
      LAYER met4 ;
        RECT 901.670 5163.385 973.330 5188.000 ;
      LAYER met4 ;
        RECT 973.730 5163.785 975.000 5188.000 ;
      LAYER met4 ;
        RECT 900.965 5083.400 974.035 5163.385 ;
        RECT 975.000 5083.400 1105.000 5188.000 ;
      LAYER met4 ;
        RECT 1105.000 5163.785 1153.205 5188.000 ;
      LAYER met4 ;
        RECT 1153.605 5163.385 1232.845 5188.000 ;
      LAYER met4 ;
        RECT 1233.245 5163.785 1274.000 5188.000 ;
      LAYER met4 ;
        RECT 1152.240 5083.400 1233.245 5163.385 ;
        RECT 1274.000 5083.400 1368.000 5188.000 ;
      LAYER met4 ;
        RECT 1368.000 5163.785 1416.205 5188.000 ;
      LAYER met4 ;
        RECT 1416.605 5163.385 1495.845 5188.000 ;
      LAYER met4 ;
        RECT 1496.245 5163.785 1537.000 5188.000 ;
      LAYER met4 ;
        RECT 1415.240 5083.400 1496.245 5163.385 ;
        RECT 1537.000 5083.400 1667.000 5188.000 ;
      LAYER met4 ;
        RECT 1667.000 5163.785 1668.270 5188.000 ;
      LAYER met4 ;
        RECT 1668.670 5163.385 1740.330 5188.000 ;
      LAYER met4 ;
        RECT 1740.730 5163.785 1742.000 5188.000 ;
      LAYER met4 ;
        RECT 1742.000 5163.785 1877.000 5188.000 ;
      LAYER met4 ;
        RECT 1877.000 5163.785 1925.205 5188.000 ;
      LAYER met4 ;
        RECT 1667.965 5083.400 1741.035 5163.385 ;
        RECT 1742.000 5083.400 1862.000 5163.785 ;
        RECT 1867.000 5083.400 1877.000 5163.785 ;
        RECT 1925.605 5163.385 2004.845 5188.000 ;
      LAYER met4 ;
        RECT 2005.245 5163.785 2046.000 5188.000 ;
      LAYER met4 ;
        RECT 1924.240 5083.400 2005.245 5163.385 ;
        RECT 2046.000 5083.400 2369.000 5188.000 ;
      LAYER met4 ;
        RECT 2369.000 5163.785 2370.270 5188.000 ;
      LAYER met4 ;
        RECT 2370.670 5163.385 2442.330 5188.000 ;
      LAYER met4 ;
        RECT 2442.730 5163.785 2444.000 5188.000 ;
      LAYER met4 ;
        RECT 2369.965 5083.400 2443.035 5163.385 ;
        RECT 2444.000 5083.400 2626.000 5188.000 ;
      LAYER met4 ;
        RECT 2626.000 5163.785 2627.270 5188.000 ;
      LAYER met4 ;
        RECT 2627.670 5163.385 2699.330 5188.000 ;
      LAYER met4 ;
        RECT 2699.730 5163.785 2701.000 5188.000 ;
      LAYER met4 ;
        RECT 2626.965 5083.400 2700.035 5163.385 ;
        RECT 2701.000 5083.400 2878.000 5188.000 ;
      LAYER met4 ;
        RECT 2878.000 5163.785 2879.270 5188.000 ;
      LAYER met4 ;
        RECT 2879.670 5163.385 2951.330 5188.000 ;
      LAYER met4 ;
        RECT 2951.730 5163.785 2953.000 5188.000 ;
      LAYER met4 ;
        RECT 2878.965 5083.400 2952.035 5163.385 ;
        RECT 2953.000 5083.400 3135.000 5188.000 ;
      LAYER met4 ;
        RECT 3135.000 5163.785 3136.270 5188.000 ;
      LAYER met4 ;
        RECT 3136.670 5163.385 3208.330 5188.000 ;
      LAYER met4 ;
        RECT 3208.730 5163.785 3210.000 5188.000 ;
      LAYER met4 ;
        RECT 3210.000 5163.385 3388.000 5188.000 ;
      LAYER met4 ;
        RECT 3388.000 5163.785 3389.435 5188.000 ;
      LAYER met4 ;
        RECT 3389.835 5163.385 3588.000 5188.000 ;
        RECT 3135.965 5083.400 3209.035 5163.385 ;
        RECT 3210.000 5083.400 3588.000 5163.385 ;
        RECT 0.000 5057.635 201.745 5083.400 ;
      LAYER met4 ;
        RECT 202.145 5058.035 387.270 5083.000 ;
      LAYER met4 ;
        RECT 387.670 5057.635 459.330 5083.400 ;
      LAYER met4 ;
        RECT 459.730 5058.035 644.270 5083.000 ;
      LAYER met4 ;
        RECT 644.670 5057.635 716.330 5083.400 ;
      LAYER met4 ;
        RECT 716.730 5058.035 901.270 5083.000 ;
      LAYER met4 ;
        RECT 901.670 5057.635 973.330 5083.400 ;
      LAYER met4 ;
        RECT 973.730 5058.035 1152.715 5083.000 ;
      LAYER met4 ;
        RECT 1153.115 5057.635 1230.485 5083.400 ;
      LAYER met4 ;
        RECT 1230.885 5058.035 1415.715 5083.000 ;
      LAYER met4 ;
        RECT 1416.115 5057.635 1493.485 5083.400 ;
      LAYER met4 ;
        RECT 1493.885 5058.035 1668.270 5083.000 ;
      LAYER met4 ;
        RECT 1668.670 5057.635 1740.330 5083.400 ;
      LAYER met4 ;
        RECT 1740.730 5058.035 1924.715 5083.000 ;
      LAYER met4 ;
        RECT 1925.115 5057.635 2002.485 5083.400 ;
      LAYER met4 ;
        RECT 2002.885 5058.035 2370.270 5083.000 ;
      LAYER met4 ;
        RECT 2370.670 5057.635 2442.330 5083.400 ;
      LAYER met4 ;
        RECT 2442.730 5058.035 2627.270 5083.000 ;
      LAYER met4 ;
        RECT 2627.670 5057.635 2699.330 5083.400 ;
      LAYER met4 ;
        RECT 2699.730 5058.035 2879.270 5083.000 ;
      LAYER met4 ;
        RECT 2879.670 5057.635 2951.330 5083.400 ;
      LAYER met4 ;
        RECT 2951.730 5058.035 3136.270 5083.000 ;
      LAYER met4 ;
        RECT 3136.670 5057.635 3208.330 5083.400 ;
      LAYER met4 ;
        RECT 3208.730 5058.035 3390.645 5083.000 ;
      LAYER met4 ;
        RECT 3391.045 5057.635 3588.000 5083.400 ;
        RECT 0.000 5056.935 202.745 5057.635 ;
        RECT 204.000 5056.935 386.000 5057.635 ;
        RECT 386.965 5056.935 460.035 5057.635 ;
        RECT 461.000 5056.935 643.000 5057.635 ;
        RECT 643.965 5056.935 717.035 5057.635 ;
        RECT 718.000 5056.935 900.000 5057.635 ;
        RECT 900.965 5056.935 974.035 5057.635 ;
        RECT 975.000 5056.935 1105.000 5057.635 ;
        RECT 1152.240 5056.935 1233.245 5057.635 ;
        RECT 1274.000 5056.935 1368.000 5057.635 ;
        RECT 1415.240 5056.935 1496.245 5057.635 ;
        RECT 1537.000 5056.935 1667.000 5057.635 ;
        RECT 1667.965 5056.935 1741.035 5057.635 ;
        RECT 1742.000 5056.935 1862.000 5057.635 ;
        RECT 1867.000 5056.935 1877.000 5057.635 ;
        RECT 1924.240 5056.935 2005.245 5057.635 ;
        RECT 2046.000 5056.935 2369.000 5057.635 ;
        RECT 2369.965 5056.935 2443.035 5057.635 ;
        RECT 2444.000 5056.935 2626.000 5057.635 ;
        RECT 2626.965 5056.935 2700.035 5057.635 ;
        RECT 2701.000 5056.935 2878.000 5057.635 ;
        RECT 2878.965 5056.935 2952.035 5057.635 ;
        RECT 2953.000 5056.935 3135.000 5057.635 ;
        RECT 3135.965 5056.935 3209.035 5057.635 ;
        RECT 3210.000 5056.935 3588.000 5057.635 ;
        RECT 0.000 5051.685 202.330 5056.935 ;
      LAYER met4 ;
        RECT 202.730 5052.085 387.270 5056.535 ;
      LAYER met4 ;
        RECT 387.670 5051.685 459.330 5056.935 ;
      LAYER met4 ;
        RECT 459.730 5052.085 644.270 5056.535 ;
      LAYER met4 ;
        RECT 644.670 5051.685 716.330 5056.935 ;
      LAYER met4 ;
        RECT 716.730 5052.085 901.270 5056.535 ;
      LAYER met4 ;
        RECT 901.670 5051.685 973.330 5056.935 ;
      LAYER met4 ;
        RECT 973.730 5052.085 1152.715 5056.535 ;
      LAYER met4 ;
        RECT 1153.115 5051.685 1230.485 5056.935 ;
      LAYER met4 ;
        RECT 1230.885 5052.085 1415.715 5056.535 ;
      LAYER met4 ;
        RECT 1416.115 5051.685 1493.485 5056.935 ;
      LAYER met4 ;
        RECT 1493.885 5052.085 1668.270 5056.535 ;
      LAYER met4 ;
        RECT 1668.670 5051.685 1740.330 5056.935 ;
      LAYER met4 ;
        RECT 1740.730 5052.085 1924.715 5056.535 ;
      LAYER met4 ;
        RECT 1925.115 5051.685 2002.485 5056.935 ;
      LAYER met4 ;
        RECT 2002.885 5052.085 2370.270 5056.535 ;
      LAYER met4 ;
        RECT 2370.670 5051.685 2442.330 5056.935 ;
      LAYER met4 ;
        RECT 2442.730 5052.085 2627.270 5056.535 ;
      LAYER met4 ;
        RECT 2627.670 5051.685 2699.330 5056.935 ;
      LAYER met4 ;
        RECT 2699.730 5052.085 2879.270 5056.535 ;
      LAYER met4 ;
        RECT 2879.670 5051.685 2951.330 5056.935 ;
      LAYER met4 ;
        RECT 2951.730 5052.085 3136.270 5056.535 ;
      LAYER met4 ;
        RECT 3136.670 5051.685 3208.330 5056.935 ;
      LAYER met4 ;
        RECT 3208.730 5052.085 3389.480 5056.535 ;
      LAYER met4 ;
        RECT 3389.880 5051.685 3588.000 5056.935 ;
        RECT 0.000 5051.085 202.745 5051.685 ;
        RECT 204.000 5051.085 386.000 5051.685 ;
        RECT 386.965 5051.085 460.035 5051.685 ;
        RECT 461.000 5051.085 643.000 5051.685 ;
        RECT 643.965 5051.085 717.035 5051.685 ;
        RECT 718.000 5051.085 900.000 5051.685 ;
        RECT 900.965 5051.085 974.035 5051.685 ;
        RECT 975.000 5051.085 1105.000 5051.685 ;
        RECT 1152.240 5051.085 1233.245 5051.685 ;
        RECT 1274.000 5051.085 1368.000 5051.685 ;
        RECT 1415.240 5051.085 1496.245 5051.685 ;
        RECT 1537.000 5051.085 1667.000 5051.685 ;
        RECT 1667.965 5051.085 1741.035 5051.685 ;
        RECT 1742.000 5051.085 1862.000 5051.685 ;
        RECT 1867.000 5051.085 1877.000 5051.685 ;
        RECT 1924.240 5051.085 2005.245 5051.685 ;
        RECT 2046.000 5051.085 2369.000 5051.685 ;
        RECT 2369.965 5051.085 2443.035 5051.685 ;
        RECT 2444.000 5051.085 2626.000 5051.685 ;
        RECT 2626.965 5051.085 2700.035 5051.685 ;
        RECT 2701.000 5051.085 2878.000 5051.685 ;
        RECT 2878.965 5051.085 2952.035 5051.685 ;
        RECT 2953.000 5051.085 3135.000 5051.685 ;
        RECT 3135.965 5051.085 3209.035 5051.685 ;
        RECT 3210.000 5051.085 3588.000 5051.685 ;
        RECT 0.000 5045.835 202.330 5051.085 ;
      LAYER met4 ;
        RECT 202.730 5046.235 387.270 5050.685 ;
      LAYER met4 ;
        RECT 387.670 5045.835 459.330 5051.085 ;
      LAYER met4 ;
        RECT 459.730 5046.235 644.270 5050.685 ;
      LAYER met4 ;
        RECT 644.670 5045.835 716.330 5051.085 ;
      LAYER met4 ;
        RECT 716.730 5046.235 901.270 5050.685 ;
      LAYER met4 ;
        RECT 901.670 5045.835 973.330 5051.085 ;
      LAYER met4 ;
        RECT 973.730 5046.235 1152.715 5050.685 ;
      LAYER met4 ;
        RECT 1153.115 5045.835 1230.485 5051.085 ;
      LAYER met4 ;
        RECT 1230.885 5046.235 1415.715 5050.685 ;
      LAYER met4 ;
        RECT 1416.115 5045.835 1493.485 5051.085 ;
      LAYER met4 ;
        RECT 1493.885 5046.235 1668.270 5050.685 ;
      LAYER met4 ;
        RECT 1668.670 5045.835 1740.330 5051.085 ;
      LAYER met4 ;
        RECT 1740.730 5046.235 1924.715 5050.685 ;
      LAYER met4 ;
        RECT 1925.115 5045.835 2002.485 5051.085 ;
      LAYER met4 ;
        RECT 2002.885 5046.235 2370.270 5050.685 ;
      LAYER met4 ;
        RECT 2370.670 5045.835 2442.330 5051.085 ;
      LAYER met4 ;
        RECT 2442.730 5046.235 2627.270 5050.685 ;
      LAYER met4 ;
        RECT 2627.670 5045.835 2699.330 5051.085 ;
      LAYER met4 ;
        RECT 2699.730 5046.235 2879.270 5050.685 ;
      LAYER met4 ;
        RECT 2879.670 5045.835 2951.330 5051.085 ;
      LAYER met4 ;
        RECT 2951.730 5046.235 3136.270 5050.685 ;
      LAYER met4 ;
        RECT 3136.670 5045.835 3208.330 5051.085 ;
      LAYER met4 ;
        RECT 3208.730 5046.235 3389.625 5050.685 ;
      LAYER met4 ;
        RECT 3390.025 5045.835 3588.000 5051.085 ;
        RECT 0.000 5045.135 202.745 5045.835 ;
        RECT 204.000 5045.135 386.000 5045.835 ;
        RECT 386.965 5045.135 460.035 5045.835 ;
        RECT 461.000 5045.135 643.000 5045.835 ;
        RECT 643.965 5045.135 717.035 5045.835 ;
        RECT 718.000 5045.135 900.000 5045.835 ;
        RECT 900.965 5045.135 974.035 5045.835 ;
        RECT 975.000 5045.135 1105.000 5045.835 ;
        RECT 1152.240 5045.135 1233.245 5045.835 ;
        RECT 1274.000 5045.135 1368.000 5045.835 ;
        RECT 1415.240 5045.135 1496.245 5045.835 ;
        RECT 1537.000 5045.135 1667.000 5045.835 ;
        RECT 1667.965 5045.135 1741.035 5045.835 ;
        RECT 1742.000 5045.135 1862.000 5045.835 ;
        RECT 1867.000 5045.135 1877.000 5045.835 ;
        RECT 1924.240 5045.135 2005.245 5045.835 ;
        RECT 2046.000 5045.135 2369.000 5045.835 ;
        RECT 2369.965 5045.135 2443.035 5045.835 ;
        RECT 2444.000 5045.135 2626.000 5045.835 ;
        RECT 2626.965 5045.135 2700.035 5045.835 ;
        RECT 2701.000 5045.135 2878.000 5045.835 ;
        RECT 2878.965 5045.135 2952.035 5045.835 ;
        RECT 2953.000 5045.135 3135.000 5045.835 ;
        RECT 3135.965 5045.135 3209.035 5045.835 ;
        RECT 3210.000 5045.135 3588.000 5045.835 ;
        RECT 0.000 5044.005 176.425 5045.135 ;
      LAYER met4 ;
        RECT 176.825 5044.405 1862.000 5044.735 ;
        RECT 1867.000 5044.405 2879.270 5044.735 ;
      LAYER met4 ;
        RECT 2879.670 5044.505 2951.330 5045.135 ;
      LAYER met4 ;
        RECT 2951.730 5044.405 3411.175 5044.735 ;
      LAYER met4 ;
        RECT 0.000 5040.725 176.690 5044.005 ;
      LAYER met4 ;
        RECT 177.090 5041.125 3410.910 5044.105 ;
      LAYER met4 ;
        RECT 3411.575 5044.005 3588.000 5045.135 ;
        RECT 0.000 5039.245 182.045 5040.725 ;
      LAYER met4 ;
        RECT 182.445 5039.645 204.000 5040.825 ;
      LAYER met4 ;
        RECT 204.000 5039.645 386.000 5040.825 ;
      LAYER met4 ;
        RECT 386.000 5039.645 387.270 5040.825 ;
      LAYER met4 ;
        RECT 387.670 5039.745 459.330 5040.725 ;
      LAYER met4 ;
        RECT 459.730 5039.645 461.000 5040.825 ;
      LAYER met4 ;
        RECT 461.000 5039.645 643.000 5040.825 ;
      LAYER met4 ;
        RECT 643.000 5039.645 644.270 5040.825 ;
      LAYER met4 ;
        RECT 644.670 5039.745 716.330 5040.725 ;
      LAYER met4 ;
        RECT 716.730 5039.645 718.000 5040.825 ;
      LAYER met4 ;
        RECT 718.000 5039.645 900.000 5040.825 ;
      LAYER met4 ;
        RECT 900.000 5039.645 901.270 5040.825 ;
      LAYER met4 ;
        RECT 901.670 5039.745 973.330 5040.725 ;
      LAYER met4 ;
        RECT 973.730 5039.645 975.000 5040.825 ;
      LAYER met4 ;
        RECT 975.000 5039.645 1105.000 5040.825 ;
      LAYER met4 ;
        RECT 1105.000 5039.645 1152.240 5040.825 ;
      LAYER met4 ;
        RECT 1152.640 5039.745 1230.485 5040.725 ;
      LAYER met4 ;
        RECT 1230.885 5039.645 1274.000 5040.825 ;
      LAYER met4 ;
        RECT 1274.000 5039.645 1368.000 5040.825 ;
      LAYER met4 ;
        RECT 1368.000 5039.645 1415.240 5040.825 ;
      LAYER met4 ;
        RECT 1415.640 5039.745 1493.485 5040.725 ;
      LAYER met4 ;
        RECT 1493.885 5039.645 1537.000 5040.825 ;
      LAYER met4 ;
        RECT 1537.000 5039.645 1667.000 5040.825 ;
      LAYER met4 ;
        RECT 1667.000 5039.645 1668.270 5040.825 ;
      LAYER met4 ;
        RECT 1668.670 5039.745 1740.330 5040.725 ;
      LAYER met4 ;
        RECT 1740.730 5039.645 1742.000 5040.825 ;
      LAYER met4 ;
        RECT 1742.000 5039.645 1862.000 5040.825 ;
        RECT 1867.000 5039.645 1877.000 5040.825 ;
      LAYER met4 ;
        RECT 1877.000 5039.645 1924.240 5040.825 ;
      LAYER met4 ;
        RECT 1924.640 5039.745 2002.485 5040.725 ;
      LAYER met4 ;
        RECT 2002.885 5039.645 2046.000 5040.825 ;
      LAYER met4 ;
        RECT 2046.000 5039.645 2369.000 5040.825 ;
      LAYER met4 ;
        RECT 2369.000 5039.645 2370.270 5040.825 ;
      LAYER met4 ;
        RECT 2370.670 5039.745 2442.330 5040.725 ;
      LAYER met4 ;
        RECT 2442.730 5039.645 2444.000 5040.825 ;
      LAYER met4 ;
        RECT 2444.000 5039.645 2626.000 5040.825 ;
      LAYER met4 ;
        RECT 2626.000 5039.645 2627.270 5040.825 ;
      LAYER met4 ;
        RECT 2627.670 5039.745 2699.330 5040.725 ;
      LAYER met4 ;
        RECT 2699.730 5039.645 2701.000 5040.825 ;
      LAYER met4 ;
        RECT 2701.000 5039.645 2878.000 5040.825 ;
      LAYER met4 ;
        RECT 2878.000 5039.645 2879.270 5040.825 ;
      LAYER met4 ;
        RECT 2879.670 5039.745 2951.330 5040.725 ;
      LAYER met4 ;
        RECT 2951.730 5039.645 2953.000 5040.825 ;
      LAYER met4 ;
        RECT 2953.000 5039.645 3135.000 5040.825 ;
      LAYER met4 ;
        RECT 3135.000 5039.645 3136.270 5040.825 ;
      LAYER met4 ;
        RECT 3136.670 5039.745 3208.330 5040.725 ;
      LAYER met4 ;
        RECT 3208.730 5039.645 3210.000 5040.825 ;
      LAYER met4 ;
        RECT 3210.000 5039.645 3388.000 5040.825 ;
      LAYER met4 ;
        RECT 3388.000 5039.645 3409.550 5040.825 ;
      LAYER met4 ;
        RECT 3411.310 5040.725 3588.000 5044.005 ;
        RECT 0.000 5036.465 182.725 5039.245 ;
        RECT 0.000 5035.335 180.025 5036.465 ;
      LAYER met4 ;
        RECT 183.125 5036.365 3408.935 5039.345 ;
      LAYER met4 ;
        RECT 3409.950 5039.245 3588.000 5040.725 ;
      LAYER met4 ;
        RECT 180.425 5035.735 1862.000 5036.065 ;
        RECT 1867.000 5035.735 2879.270 5036.065 ;
      LAYER met4 ;
        RECT 2879.670 5035.335 2951.330 5035.965 ;
      LAYER met4 ;
        RECT 2951.730 5035.735 3407.575 5036.065 ;
      LAYER met4 ;
        RECT 3409.335 5035.965 3588.000 5039.245 ;
        RECT 3407.975 5035.335 3588.000 5035.965 ;
        RECT 0.000 5034.635 202.745 5035.335 ;
        RECT 386.965 5034.635 460.035 5035.335 ;
        RECT 643.965 5034.635 717.035 5035.335 ;
        RECT 900.965 5034.635 974.035 5035.335 ;
        RECT 1152.240 5034.635 1233.245 5035.335 ;
        RECT 1415.240 5034.635 1496.245 5035.335 ;
        RECT 1667.965 5034.635 1741.035 5035.335 ;
        RECT 1924.240 5034.635 2005.245 5035.335 ;
        RECT 2369.965 5034.635 2443.035 5035.335 ;
        RECT 2626.965 5034.635 2700.035 5035.335 ;
        RECT 2878.965 5034.635 2952.035 5035.335 ;
        RECT 3135.965 5034.635 3209.035 5035.335 ;
        RECT 3388.000 5034.635 3588.000 5035.335 ;
        RECT 0.000 5029.185 202.330 5034.635 ;
      LAYER met4 ;
        RECT 202.730 5029.585 387.270 5034.235 ;
      LAYER met4 ;
        RECT 387.670 5029.185 459.330 5034.635 ;
      LAYER met4 ;
        RECT 459.730 5029.585 644.270 5034.235 ;
      LAYER met4 ;
        RECT 644.670 5029.185 716.330 5034.635 ;
      LAYER met4 ;
        RECT 716.730 5029.585 901.270 5034.235 ;
      LAYER met4 ;
        RECT 901.670 5029.185 973.330 5034.635 ;
      LAYER met4 ;
        RECT 973.730 5029.585 1152.250 5034.235 ;
      LAYER met4 ;
        RECT 1152.650 5029.185 1230.485 5034.635 ;
      LAYER met4 ;
        RECT 1230.885 5029.585 1415.250 5034.235 ;
      LAYER met4 ;
        RECT 1415.650 5029.185 1493.485 5034.635 ;
      LAYER met4 ;
        RECT 1493.885 5029.585 1668.270 5034.235 ;
      LAYER met4 ;
        RECT 1668.670 5029.185 1740.330 5034.635 ;
      LAYER met4 ;
        RECT 1740.730 5029.585 1924.250 5034.235 ;
      LAYER met4 ;
        RECT 1924.650 5029.185 2002.485 5034.635 ;
      LAYER met4 ;
        RECT 2002.885 5029.585 2370.270 5034.235 ;
      LAYER met4 ;
        RECT 2370.670 5029.185 2442.330 5034.635 ;
      LAYER met4 ;
        RECT 2442.730 5029.585 2627.270 5034.235 ;
      LAYER met4 ;
        RECT 2627.670 5029.185 2699.330 5034.635 ;
      LAYER met4 ;
        RECT 2699.730 5029.585 2879.270 5034.235 ;
      LAYER met4 ;
        RECT 2879.670 5029.185 2951.330 5034.635 ;
      LAYER met4 ;
        RECT 2951.730 5029.585 3136.270 5034.235 ;
      LAYER met4 ;
        RECT 3136.670 5029.185 3208.330 5034.635 ;
      LAYER met4 ;
        RECT 3208.730 5029.585 3389.475 5034.235 ;
      LAYER met4 ;
        RECT 3389.875 5029.185 3588.000 5034.635 ;
        RECT 0.000 5028.585 202.745 5029.185 ;
        RECT 386.965 5028.585 460.035 5029.185 ;
        RECT 643.965 5028.585 717.035 5029.185 ;
        RECT 900.965 5028.585 974.035 5029.185 ;
        RECT 1152.240 5028.585 1233.245 5029.185 ;
        RECT 1415.240 5028.585 1496.245 5029.185 ;
        RECT 1667.965 5028.585 1741.035 5029.185 ;
        RECT 1924.240 5028.585 2005.245 5029.185 ;
        RECT 2369.965 5028.585 2443.035 5029.185 ;
        RECT 2626.965 5028.585 2700.035 5029.185 ;
        RECT 2878.965 5028.585 2952.035 5029.185 ;
        RECT 3135.965 5028.585 3209.035 5029.185 ;
        RECT 3388.000 5028.585 3588.000 5029.185 ;
        RECT 0.000 5024.335 202.330 5028.585 ;
      LAYER met4 ;
        RECT 202.730 5024.735 387.270 5028.185 ;
      LAYER met4 ;
        RECT 387.670 5024.335 459.330 5028.585 ;
      LAYER met4 ;
        RECT 459.730 5024.735 644.270 5028.185 ;
      LAYER met4 ;
        RECT 644.670 5024.335 716.330 5028.585 ;
      LAYER met4 ;
        RECT 716.730 5024.735 901.270 5028.185 ;
      LAYER met4 ;
        RECT 901.670 5024.335 973.330 5028.585 ;
      LAYER met4 ;
        RECT 973.730 5024.735 1152.715 5028.185 ;
      LAYER met4 ;
        RECT 1153.115 5024.335 1230.485 5028.585 ;
      LAYER met4 ;
        RECT 1230.885 5024.735 1415.715 5028.185 ;
      LAYER met4 ;
        RECT 1416.115 5024.335 1493.485 5028.585 ;
      LAYER met4 ;
        RECT 1493.885 5024.735 1668.270 5028.185 ;
      LAYER met4 ;
        RECT 1668.670 5024.335 1740.330 5028.585 ;
      LAYER met4 ;
        RECT 1740.730 5024.735 1862.000 5028.185 ;
        RECT 1867.000 5024.735 1924.715 5028.185 ;
      LAYER met4 ;
        RECT 1925.115 5024.335 2002.485 5028.585 ;
      LAYER met4 ;
        RECT 2002.885 5024.735 2370.270 5028.185 ;
      LAYER met4 ;
        RECT 2370.670 5024.335 2442.330 5028.585 ;
      LAYER met4 ;
        RECT 2442.730 5024.735 2627.270 5028.185 ;
      LAYER met4 ;
        RECT 2627.670 5024.335 2699.330 5028.585 ;
      LAYER met4 ;
        RECT 2699.730 5024.735 2879.270 5028.185 ;
      LAYER met4 ;
        RECT 2879.670 5024.335 2951.330 5028.585 ;
      LAYER met4 ;
        RECT 2951.730 5024.735 3136.270 5028.185 ;
      LAYER met4 ;
        RECT 3136.670 5024.335 3208.330 5028.585 ;
      LAYER met4 ;
        RECT 3208.730 5024.735 3389.335 5028.185 ;
      LAYER met4 ;
        RECT 3389.735 5024.335 3588.000 5028.585 ;
        RECT 0.000 5023.735 202.745 5024.335 ;
        RECT 386.965 5023.735 460.035 5024.335 ;
        RECT 643.965 5023.735 717.035 5024.335 ;
        RECT 900.965 5023.735 974.035 5024.335 ;
        RECT 1152.240 5023.735 1233.245 5024.335 ;
        RECT 1415.240 5023.735 1496.245 5024.335 ;
        RECT 1667.965 5023.735 1741.035 5024.335 ;
        RECT 1924.240 5023.735 2005.245 5024.335 ;
        RECT 2369.965 5023.735 2443.035 5024.335 ;
        RECT 2626.965 5023.735 2700.035 5024.335 ;
        RECT 2878.965 5023.735 2952.035 5024.335 ;
        RECT 3135.965 5023.735 3209.035 5024.335 ;
        RECT 3388.000 5023.735 3588.000 5024.335 ;
        RECT 0.000 5019.485 202.330 5023.735 ;
      LAYER met4 ;
        RECT 202.730 5019.885 387.270 5023.335 ;
      LAYER met4 ;
        RECT 387.670 5019.485 459.330 5023.735 ;
      LAYER met4 ;
        RECT 459.730 5019.885 644.270 5023.335 ;
      LAYER met4 ;
        RECT 644.670 5019.485 716.330 5023.735 ;
      LAYER met4 ;
        RECT 716.730 5019.885 901.270 5023.335 ;
      LAYER met4 ;
        RECT 901.670 5019.485 973.330 5023.735 ;
      LAYER met4 ;
        RECT 973.730 5019.885 1152.715 5023.335 ;
      LAYER met4 ;
        RECT 1153.115 5019.485 1230.485 5023.735 ;
      LAYER met4 ;
        RECT 1230.885 5019.885 1415.715 5023.335 ;
      LAYER met4 ;
        RECT 1416.115 5019.485 1493.485 5023.735 ;
      LAYER met4 ;
        RECT 1493.885 5019.885 1668.270 5023.335 ;
      LAYER met4 ;
        RECT 1668.670 5019.485 1740.330 5023.735 ;
      LAYER met4 ;
        RECT 1740.730 5019.885 1924.715 5023.335 ;
      LAYER met4 ;
        RECT 1925.115 5019.485 2002.485 5023.735 ;
      LAYER met4 ;
        RECT 2002.885 5019.885 2370.270 5023.335 ;
      LAYER met4 ;
        RECT 2370.670 5019.485 2442.330 5023.735 ;
      LAYER met4 ;
        RECT 2442.730 5019.885 2627.270 5023.335 ;
      LAYER met4 ;
        RECT 2627.670 5019.485 2699.330 5023.735 ;
      LAYER met4 ;
        RECT 2699.730 5019.885 2879.270 5023.335 ;
      LAYER met4 ;
        RECT 2879.670 5019.485 2951.330 5023.735 ;
      LAYER met4 ;
        RECT 2951.730 5019.885 3136.270 5023.335 ;
      LAYER met4 ;
        RECT 3136.670 5019.485 3208.330 5023.735 ;
      LAYER met4 ;
        RECT 3208.730 5019.885 3389.385 5023.335 ;
      LAYER met4 ;
        RECT 3389.785 5019.485 3588.000 5023.735 ;
        RECT 0.000 5018.885 202.745 5019.485 ;
        RECT 386.965 5018.885 460.035 5019.485 ;
        RECT 643.965 5018.885 717.035 5019.485 ;
        RECT 900.965 5018.885 974.035 5019.485 ;
        RECT 1152.240 5018.885 1233.245 5019.485 ;
        RECT 1415.240 5018.885 1496.245 5019.485 ;
        RECT 1667.965 5018.885 1741.035 5019.485 ;
        RECT 1924.240 5018.885 2005.245 5019.485 ;
        RECT 2369.965 5018.885 2443.035 5019.485 ;
        RECT 2626.965 5018.885 2700.035 5019.485 ;
        RECT 2878.965 5018.885 2952.035 5019.485 ;
        RECT 3135.965 5018.885 3209.035 5019.485 ;
        RECT 3388.000 5018.885 3588.000 5019.485 ;
        RECT 0.000 5013.435 202.330 5018.885 ;
      LAYER met4 ;
        RECT 202.730 5013.835 387.270 5018.485 ;
      LAYER met4 ;
        RECT 387.670 5013.435 459.330 5018.885 ;
      LAYER met4 ;
        RECT 459.730 5013.835 644.270 5018.485 ;
      LAYER met4 ;
        RECT 644.670 5013.435 716.330 5018.885 ;
      LAYER met4 ;
        RECT 716.730 5013.835 901.270 5018.485 ;
      LAYER met4 ;
        RECT 901.670 5013.435 973.330 5018.885 ;
      LAYER met4 ;
        RECT 973.730 5013.835 1152.715 5018.485 ;
      LAYER met4 ;
        RECT 1153.115 5013.435 1230.485 5018.885 ;
      LAYER met4 ;
        RECT 1230.885 5013.835 1415.715 5018.485 ;
      LAYER met4 ;
        RECT 1416.115 5013.435 1493.485 5018.885 ;
      LAYER met4 ;
        RECT 1493.885 5013.835 1668.270 5018.485 ;
      LAYER met4 ;
        RECT 1668.670 5013.435 1740.330 5018.885 ;
      LAYER met4 ;
        RECT 1740.730 5013.835 1924.715 5018.485 ;
      LAYER met4 ;
        RECT 1925.115 5013.435 2002.485 5018.885 ;
      LAYER met4 ;
        RECT 2002.885 5013.835 2370.270 5018.485 ;
      LAYER met4 ;
        RECT 2370.670 5013.435 2442.330 5018.885 ;
      LAYER met4 ;
        RECT 2442.730 5013.835 2627.270 5018.485 ;
      LAYER met4 ;
        RECT 2627.670 5013.435 2699.330 5018.885 ;
      LAYER met4 ;
        RECT 2699.730 5013.835 2879.270 5018.485 ;
      LAYER met4 ;
        RECT 2879.670 5013.435 2951.330 5018.885 ;
      LAYER met4 ;
        RECT 2951.730 5013.835 3136.270 5018.485 ;
      LAYER met4 ;
        RECT 3136.670 5013.435 3208.330 5018.885 ;
      LAYER met4 ;
        RECT 3208.730 5013.835 3389.600 5018.485 ;
      LAYER met4 ;
        RECT 3390.000 5013.435 3588.000 5018.885 ;
        RECT 0.000 5012.835 202.745 5013.435 ;
        RECT 386.965 5012.835 460.035 5013.435 ;
        RECT 643.965 5012.835 717.035 5013.435 ;
        RECT 900.965 5012.835 974.035 5013.435 ;
        RECT 1152.240 5012.835 1233.245 5013.435 ;
        RECT 1415.240 5012.835 1496.245 5013.435 ;
        RECT 1667.965 5012.835 1741.035 5013.435 ;
        RECT 1924.240 5012.835 2005.245 5013.435 ;
        RECT 2369.965 5012.835 2443.035 5013.435 ;
        RECT 2626.965 5012.835 2700.035 5013.435 ;
        RECT 2878.965 5012.835 2952.035 5013.435 ;
        RECT 3135.965 5012.835 3209.035 5013.435 ;
        RECT 3388.000 5012.835 3588.000 5013.435 ;
        RECT 0.000 5011.575 202.330 5012.835 ;
        RECT 0.000 4991.045 142.865 5011.575 ;
        RECT 143.995 5011.310 202.330 5011.575 ;
        RECT 0.000 4989.835 104.600 4991.045 ;
      LAYER met4 ;
        RECT 0.000 4988.000 24.215 4989.435 ;
      LAYER met4 ;
        RECT 24.615 4988.000 104.600 4989.835 ;
        RECT 0.000 4851.000 104.600 4988.000 ;
      LAYER met4 ;
        RECT 0.000 4849.730 24.215 4851.000 ;
      LAYER met4 ;
        RECT 24.615 4849.330 104.600 4850.035 ;
      LAYER met4 ;
        RECT 105.000 4849.730 129.965 4990.645 ;
      LAYER met4 ;
        RECT 130.365 4990.025 142.865 4991.045 ;
        RECT 130.365 4989.880 136.915 4990.025 ;
        RECT 130.365 4851.000 131.065 4989.880 ;
        RECT 130.365 4849.330 131.065 4850.035 ;
      LAYER met4 ;
        RECT 131.465 4849.730 135.915 4989.480 ;
      LAYER met4 ;
        RECT 136.315 4851.000 136.915 4989.880 ;
        RECT 136.315 4849.330 136.915 4850.035 ;
      LAYER met4 ;
        RECT 137.315 4849.730 141.765 4989.625 ;
      LAYER met4 ;
        RECT 142.165 4851.000 142.865 4990.025 ;
        RECT 142.165 4849.330 142.865 4850.035 ;
        RECT 0.000 4777.670 142.865 4849.330 ;
      LAYER met4 ;
        RECT 0.000 4776.000 24.215 4777.270 ;
      LAYER met4 ;
        RECT 24.615 4776.965 104.600 4777.670 ;
        RECT 0.000 4635.000 104.600 4776.000 ;
      LAYER met4 ;
        RECT 105.000 4635.000 129.965 4777.270 ;
      LAYER met4 ;
        RECT 130.365 4776.965 131.065 4777.670 ;
        RECT 130.365 4635.000 131.065 4776.000 ;
      LAYER met4 ;
        RECT 131.465 4635.000 135.915 4777.270 ;
      LAYER met4 ;
        RECT 136.315 4776.965 136.915 4777.670 ;
        RECT 136.315 4635.000 136.915 4776.000 ;
      LAYER met4 ;
        RECT 137.315 4635.000 141.765 4777.270 ;
      LAYER met4 ;
        RECT 142.165 4776.965 142.865 4777.670 ;
        RECT 142.165 4635.000 142.865 4776.000 ;
      LAYER met4 ;
        RECT 143.265 4635.000 143.595 5011.175 ;
        RECT 143.895 4635.000 146.875 5010.910 ;
      LAYER met4 ;
        RECT 147.275 5009.950 202.330 5011.310 ;
      LAYER met4 ;
        RECT 147.175 4988.000 148.355 5009.550 ;
      LAYER met4 ;
        RECT 148.755 5009.335 202.330 5009.950 ;
        RECT 147.175 4851.000 148.355 4988.000 ;
      LAYER met4 ;
        RECT 147.175 4849.730 148.355 4851.000 ;
      LAYER met4 ;
        RECT 147.275 4777.670 148.255 4849.330 ;
      LAYER met4 ;
        RECT 147.175 4776.000 148.355 4777.270 ;
      LAYER met4 ;
        RECT 147.175 4635.000 148.355 4776.000 ;
      LAYER met4 ;
        RECT 148.655 4635.000 151.635 5008.935 ;
      LAYER met4 ;
        RECT 152.035 5007.975 202.330 5009.335 ;
      LAYER met4 ;
        RECT 151.935 4635.000 152.265 5007.575 ;
      LAYER met4 ;
        RECT 152.665 5007.385 202.330 5007.975 ;
      LAYER met4 ;
        RECT 202.730 5007.785 387.270 5012.435 ;
      LAYER met4 ;
        RECT 387.670 5007.385 459.330 5012.835 ;
      LAYER met4 ;
        RECT 459.730 5007.785 644.270 5012.435 ;
      LAYER met4 ;
        RECT 644.670 5007.385 716.330 5012.835 ;
      LAYER met4 ;
        RECT 716.730 5007.785 901.270 5012.435 ;
      LAYER met4 ;
        RECT 901.670 5007.385 973.330 5012.835 ;
      LAYER met4 ;
        RECT 973.730 5007.785 1152.715 5012.435 ;
      LAYER met4 ;
        RECT 1153.115 5007.385 1225.805 5012.835 ;
      LAYER met4 ;
        RECT 1226.205 5007.785 1415.715 5012.435 ;
      LAYER met4 ;
        RECT 1416.115 5007.385 1488.805 5012.835 ;
      LAYER met4 ;
        RECT 1489.205 5007.785 1668.270 5012.435 ;
      LAYER met4 ;
        RECT 1668.670 5007.385 1740.330 5012.835 ;
      LAYER met4 ;
        RECT 1740.730 5007.785 1924.715 5012.435 ;
      LAYER met4 ;
        RECT 1925.115 5007.385 1997.805 5012.835 ;
      LAYER met4 ;
        RECT 1998.205 5007.785 2370.270 5012.435 ;
      LAYER met4 ;
        RECT 2370.670 5007.385 2442.330 5012.835 ;
      LAYER met4 ;
        RECT 2442.730 5007.785 2627.270 5012.435 ;
      LAYER met4 ;
        RECT 2627.670 5007.385 2699.330 5012.835 ;
      LAYER met4 ;
        RECT 2699.730 5007.785 2879.270 5012.435 ;
      LAYER met4 ;
        RECT 2879.670 5007.385 2951.330 5012.835 ;
      LAYER met4 ;
        RECT 2951.730 5007.785 3136.270 5012.435 ;
      LAYER met4 ;
        RECT 3136.670 5007.385 3208.330 5012.835 ;
      LAYER met4 ;
        RECT 3208.730 5007.785 3389.525 5012.435 ;
      LAYER met4 ;
        RECT 3389.925 5011.575 3588.000 5012.835 ;
        RECT 3389.925 5011.310 3444.005 5011.575 ;
        RECT 3389.925 5007.975 3440.725 5011.310 ;
        RECT 3389.925 5007.385 3435.335 5007.975 ;
        RECT 152.665 5006.785 202.745 5007.385 ;
        RECT 386.965 5006.785 460.035 5007.385 ;
        RECT 643.965 5006.785 717.035 5007.385 ;
        RECT 900.965 5006.785 974.035 5007.385 ;
        RECT 1152.240 5006.785 1233.245 5007.385 ;
        RECT 1415.240 5006.785 1496.245 5007.385 ;
        RECT 1667.965 5006.785 1741.035 5007.385 ;
        RECT 1924.240 5006.785 2005.245 5007.385 ;
        RECT 2369.965 5006.785 2443.035 5007.385 ;
        RECT 2626.965 5006.785 2700.035 5007.385 ;
        RECT 2878.965 5006.785 2952.035 5007.385 ;
        RECT 3135.965 5006.785 3209.035 5007.385 ;
        RECT 3388.000 5006.785 3435.335 5007.385 ;
        RECT 152.665 5002.535 202.345 5006.785 ;
      LAYER met4 ;
        RECT 202.745 5002.935 386.965 5006.385 ;
      LAYER met4 ;
        RECT 387.365 5002.535 459.635 5006.785 ;
      LAYER met4 ;
        RECT 460.035 5002.935 643.965 5006.385 ;
      LAYER met4 ;
        RECT 644.365 5002.535 716.635 5006.785 ;
      LAYER met4 ;
        RECT 717.035 5002.935 900.965 5006.385 ;
      LAYER met4 ;
        RECT 901.365 5002.535 973.635 5006.785 ;
      LAYER met4 ;
        RECT 974.035 5002.935 1152.715 5006.385 ;
      LAYER met4 ;
        RECT 1153.115 5002.535 1225.805 5006.785 ;
      LAYER met4 ;
        RECT 1226.205 5002.935 1415.715 5006.385 ;
      LAYER met4 ;
        RECT 1416.115 5002.535 1488.805 5006.785 ;
      LAYER met4 ;
        RECT 1489.205 5002.935 1667.965 5006.385 ;
      LAYER met4 ;
        RECT 1668.365 5002.535 1740.635 5006.785 ;
      LAYER met4 ;
        RECT 1741.035 5002.935 1862.000 5006.385 ;
        RECT 1867.000 5002.935 1924.715 5006.385 ;
      LAYER met4 ;
        RECT 1925.115 5002.535 1997.805 5006.785 ;
      LAYER met4 ;
        RECT 1998.205 5002.935 2369.965 5006.385 ;
      LAYER met4 ;
        RECT 2370.365 5002.535 2442.635 5006.785 ;
      LAYER met4 ;
        RECT 2443.035 5002.935 2626.965 5006.385 ;
      LAYER met4 ;
        RECT 2627.365 5002.535 2699.635 5006.785 ;
      LAYER met4 ;
        RECT 2700.035 5002.935 2878.965 5006.385 ;
      LAYER met4 ;
        RECT 2879.365 5002.535 2951.635 5006.785 ;
      LAYER met4 ;
        RECT 2952.035 5002.935 3135.965 5006.385 ;
      LAYER met4 ;
        RECT 3136.365 5002.535 3208.635 5006.785 ;
      LAYER met4 ;
        RECT 3209.035 5002.935 3389.470 5006.385 ;
      LAYER met4 ;
        RECT 3389.870 5002.535 3435.335 5006.785 ;
        RECT 152.665 5001.935 202.745 5002.535 ;
        RECT 386.965 5001.935 460.035 5002.535 ;
        RECT 643.965 5001.935 717.035 5002.535 ;
        RECT 900.965 5001.935 974.035 5002.535 ;
        RECT 1152.240 5001.935 1233.245 5002.535 ;
        RECT 1415.240 5001.935 1496.245 5002.535 ;
        RECT 1667.965 5001.935 1741.035 5002.535 ;
        RECT 1924.240 5001.935 2005.245 5002.535 ;
        RECT 2369.965 5001.935 2443.035 5002.535 ;
        RECT 2626.965 5001.935 2700.035 5002.535 ;
        RECT 2878.965 5001.935 2952.035 5002.535 ;
        RECT 3135.965 5001.935 3209.035 5002.535 ;
        RECT 3388.000 5001.935 3435.335 5002.535 ;
        RECT 152.665 4996.485 202.330 5001.935 ;
      LAYER met4 ;
        RECT 202.730 4996.885 387.270 5001.535 ;
      LAYER met4 ;
        RECT 387.670 4996.485 459.330 5001.935 ;
      LAYER met4 ;
        RECT 459.730 4996.885 644.270 5001.535 ;
      LAYER met4 ;
        RECT 644.670 4996.485 716.330 5001.935 ;
      LAYER met4 ;
        RECT 716.730 4996.885 901.270 5001.535 ;
      LAYER met4 ;
        RECT 901.670 4996.485 973.330 5001.935 ;
      LAYER met4 ;
        RECT 973.730 4996.885 1152.715 5001.535 ;
      LAYER met4 ;
        RECT 1153.115 4996.485 1230.485 5001.935 ;
      LAYER met4 ;
        RECT 1230.885 4996.885 1415.715 5001.535 ;
      LAYER met4 ;
        RECT 1416.115 4996.485 1493.485 5001.935 ;
      LAYER met4 ;
        RECT 1493.885 4996.885 1668.270 5001.535 ;
      LAYER met4 ;
        RECT 1668.670 4996.485 1740.330 5001.935 ;
      LAYER met4 ;
        RECT 1740.730 4996.885 1924.715 5001.535 ;
      LAYER met4 ;
        RECT 1925.115 4996.485 2002.485 5001.935 ;
      LAYER met4 ;
        RECT 2002.885 4996.885 2370.270 5001.535 ;
      LAYER met4 ;
        RECT 2370.670 4996.485 2442.330 5001.935 ;
      LAYER met4 ;
        RECT 2442.730 4996.885 2627.270 5001.535 ;
      LAYER met4 ;
        RECT 2627.670 4996.485 2699.330 5001.935 ;
      LAYER met4 ;
        RECT 2699.730 4996.885 2879.270 5001.535 ;
      LAYER met4 ;
        RECT 2879.670 4996.485 2951.330 5001.935 ;
      LAYER met4 ;
        RECT 2951.730 4996.885 3136.270 5001.535 ;
      LAYER met4 ;
        RECT 3136.670 4996.485 3208.330 5001.935 ;
      LAYER met4 ;
        RECT 3208.730 4996.885 3391.785 5001.535 ;
      LAYER met4 ;
        RECT 3392.185 4996.485 3435.335 5001.935 ;
        RECT 152.665 4995.885 202.745 4996.485 ;
        RECT 386.965 4995.885 460.035 4996.485 ;
        RECT 643.965 4995.885 717.035 4996.485 ;
        RECT 900.965 4995.885 974.035 4996.485 ;
        RECT 1152.240 4995.885 1233.245 4996.485 ;
        RECT 1415.240 4995.885 1496.245 4996.485 ;
        RECT 1667.965 4995.885 1741.035 4996.485 ;
        RECT 1924.240 4995.885 2005.245 4996.485 ;
        RECT 2369.965 4995.885 2443.035 4996.485 ;
        RECT 2626.965 4995.885 2700.035 4996.485 ;
        RECT 2878.965 4995.885 2952.035 4996.485 ;
        RECT 3135.965 4995.885 3209.035 4996.485 ;
        RECT 3388.000 4995.885 3435.335 4996.485 ;
        RECT 152.665 4992.185 202.330 4995.885 ;
        RECT 152.665 4990.000 186.065 4992.185 ;
        RECT 152.665 4989.875 169.115 4990.000 ;
        RECT 152.665 4988.000 153.365 4989.875 ;
        RECT 158.815 4989.785 169.115 4989.875 ;
        RECT 158.815 4989.735 164.265 4989.785 ;
        RECT 152.665 4849.330 153.365 4850.035 ;
      LAYER met4 ;
        RECT 153.765 4849.730 158.415 4989.475 ;
      LAYER met4 ;
        RECT 158.815 4988.000 159.415 4989.735 ;
        RECT 158.815 4849.330 159.415 4850.035 ;
      LAYER met4 ;
        RECT 159.815 4849.730 163.265 4989.335 ;
      LAYER met4 ;
        RECT 163.665 4988.000 164.265 4989.735 ;
        RECT 163.665 4849.330 164.265 4850.035 ;
      LAYER met4 ;
        RECT 164.665 4849.730 168.115 4989.385 ;
      LAYER met4 ;
        RECT 168.515 4988.000 169.115 4989.785 ;
        RECT 174.565 4989.925 186.065 4990.000 ;
        RECT 168.515 4849.330 169.115 4850.035 ;
      LAYER met4 ;
        RECT 169.515 4849.730 174.165 4989.600 ;
      LAYER met4 ;
        RECT 174.565 4988.000 175.165 4989.925 ;
        RECT 180.615 4989.870 186.065 4989.925 ;
        RECT 174.565 4849.330 175.165 4850.035 ;
      LAYER met4 ;
        RECT 175.565 4849.730 180.215 4989.525 ;
      LAYER met4 ;
        RECT 180.615 4988.000 181.215 4989.870 ;
      LAYER met4 ;
        RECT 181.615 4850.035 185.065 4989.470 ;
      LAYER met4 ;
        RECT 185.465 4988.000 186.065 4989.870 ;
        RECT 180.615 4849.635 181.215 4850.035 ;
        RECT 185.465 4849.635 186.065 4850.035 ;
      LAYER met4 ;
        RECT 186.465 4849.730 191.115 4991.785 ;
      LAYER met4 ;
        RECT 191.515 4990.750 202.330 4992.185 ;
        RECT 191.515 4988.000 192.115 4990.750 ;
        RECT 180.615 4849.330 186.065 4849.635 ;
        RECT 191.515 4849.330 192.115 4850.035 ;
      LAYER met4 ;
        RECT 192.515 4849.730 197.965 4990.350 ;
      LAYER met4 ;
        RECT 198.365 4990.035 202.330 4990.750 ;
      LAYER met4 ;
        RECT 202.730 4990.035 387.270 4995.485 ;
      LAYER met4 ;
        RECT 387.670 4990.035 459.330 4995.885 ;
      LAYER met4 ;
        RECT 459.730 4990.035 644.270 4995.485 ;
      LAYER met4 ;
        RECT 644.670 4990.035 716.330 4995.885 ;
      LAYER met4 ;
        RECT 716.730 4990.035 901.270 4995.485 ;
      LAYER met4 ;
        RECT 901.670 4990.035 973.330 4995.885 ;
      LAYER met4 ;
        RECT 973.730 4990.035 1152.715 4995.485 ;
      LAYER met4 ;
        RECT 1153.115 4990.035 1230.485 4995.885 ;
      LAYER met4 ;
        RECT 1230.885 4990.035 1415.715 4995.485 ;
      LAYER met4 ;
        RECT 1416.115 4990.035 1493.485 4995.885 ;
      LAYER met4 ;
        RECT 1493.885 4990.035 1668.270 4995.485 ;
      LAYER met4 ;
        RECT 1668.670 4990.035 1740.330 4995.885 ;
      LAYER met4 ;
        RECT 1740.730 4990.035 1924.715 4995.485 ;
      LAYER met4 ;
        RECT 1925.115 4990.035 2002.485 4995.885 ;
      LAYER met4 ;
        RECT 2002.885 4990.035 2370.270 4995.485 ;
      LAYER met4 ;
        RECT 2370.670 4990.035 2442.330 4995.885 ;
      LAYER met4 ;
        RECT 2442.730 4990.035 2627.270 4995.485 ;
      LAYER met4 ;
        RECT 2627.670 4990.035 2699.330 4995.885 ;
      LAYER met4 ;
        RECT 2699.730 4990.035 2879.270 4995.485 ;
      LAYER met4 ;
        RECT 2879.670 4990.035 2951.330 4995.885 ;
      LAYER met4 ;
        RECT 2951.730 4990.035 3136.270 4995.485 ;
      LAYER met4 ;
        RECT 3136.670 4990.035 3208.330 4995.885 ;
      LAYER met4 ;
        RECT 3208.730 4990.035 3390.350 4995.485 ;
      LAYER met4 ;
        RECT 197.965 4989.635 202.330 4990.035 ;
        POLYGON 3388.000 4990.035 3388.400 4990.035 3388.400 4989.635 ;
        RECT 3388.400 4989.635 3390.035 4990.035 ;
        RECT 3390.750 4989.635 3435.335 4995.885 ;
        RECT 197.965 4988.400 202.745 4989.635 ;
        POLYGON 197.965 4988.400 198.365 4988.400 197.965 4988.000 ;
        RECT 198.365 4988.000 202.745 4988.400 ;
        RECT 3388.000 4985.670 3435.335 4989.635 ;
        RECT 3388.000 4985.255 3389.635 4985.670 ;
        RECT 152.665 4777.670 197.965 4849.330 ;
      LAYER met4 ;
        RECT 3390.035 4831.730 3395.485 4985.270 ;
      LAYER met4 ;
        RECT 3395.885 4985.255 3396.485 4985.670 ;
        RECT 3401.935 4985.655 3407.385 4985.670 ;
        RECT 3395.885 4831.330 3396.485 4832.035 ;
      LAYER met4 ;
        RECT 3396.885 4831.730 3401.535 4985.270 ;
      LAYER met4 ;
        RECT 3401.935 4985.255 3402.535 4985.655 ;
        RECT 3406.785 4985.255 3407.385 4985.655 ;
      LAYER met4 ;
        RECT 3402.935 4832.035 3406.385 4985.255 ;
      LAYER met4 ;
        RECT 3401.935 4831.635 3402.535 4832.035 ;
        RECT 3406.785 4831.635 3407.385 4832.035 ;
      LAYER met4 ;
        RECT 3407.785 4831.730 3412.435 4985.270 ;
      LAYER met4 ;
        RECT 3412.835 4985.255 3413.435 4985.670 ;
        RECT 3401.935 4831.330 3407.385 4831.635 ;
        RECT 3412.835 4831.330 3413.435 4832.035 ;
      LAYER met4 ;
        RECT 3413.835 4831.730 3418.485 4985.270 ;
      LAYER met4 ;
        RECT 3418.885 4985.255 3419.485 4985.670 ;
        RECT 3418.885 4831.330 3419.485 4832.035 ;
      LAYER met4 ;
        RECT 3419.885 4831.730 3423.335 4985.270 ;
      LAYER met4 ;
        RECT 3423.735 4985.255 3424.335 4985.670 ;
        RECT 3423.735 4831.330 3424.335 4832.035 ;
      LAYER met4 ;
        RECT 3424.735 4831.730 3428.185 4985.270 ;
      LAYER met4 ;
        RECT 3428.585 4985.255 3429.185 4985.670 ;
        RECT 3428.585 4831.330 3429.185 4832.035 ;
      LAYER met4 ;
        RECT 3429.585 4831.730 3434.235 4985.270 ;
      LAYER met4 ;
        RECT 3434.635 4985.255 3435.335 4985.670 ;
        RECT 3434.635 4831.330 3435.335 4832.035 ;
        RECT 152.665 4776.965 153.365 4777.670 ;
      LAYER met4 ;
        RECT 153.765 4635.000 158.415 4777.270 ;
      LAYER met4 ;
        RECT 158.815 4776.965 159.415 4777.670 ;
      LAYER met4 ;
        RECT 159.815 4635.000 163.265 4777.270 ;
      LAYER met4 ;
        RECT 163.665 4776.965 164.265 4777.670 ;
      LAYER met4 ;
        RECT 164.665 4635.000 168.115 4777.270 ;
      LAYER met4 ;
        RECT 168.515 4776.965 169.115 4777.670 ;
      LAYER met4 ;
        RECT 169.515 4635.000 174.165 4777.270 ;
      LAYER met4 ;
        RECT 174.565 4776.965 175.165 4777.670 ;
        RECT 180.615 4777.365 186.065 4777.670 ;
      LAYER met4 ;
        RECT 175.565 4635.000 180.215 4777.270 ;
      LAYER met4 ;
        RECT 180.615 4776.965 181.215 4777.365 ;
        RECT 185.465 4776.965 186.065 4777.365 ;
      LAYER met4 ;
        RECT 181.615 4635.000 185.065 4776.965 ;
        RECT 186.465 4635.000 191.115 4777.270 ;
      LAYER met4 ;
        RECT 191.515 4776.965 192.115 4777.670 ;
      LAYER met4 ;
        RECT 192.515 4635.000 197.965 4777.270 ;
      LAYER met4 ;
        RECT 3390.035 4759.670 3435.335 4831.330 ;
      LAYER met4 ;
        RECT 3390.035 4613.000 3395.485 4759.270 ;
      LAYER met4 ;
        RECT 3395.885 4758.965 3396.485 4759.670 ;
        RECT 3401.935 4759.365 3407.385 4759.670 ;
      LAYER met4 ;
        RECT 3396.885 4613.000 3401.535 4759.270 ;
      LAYER met4 ;
        RECT 3401.935 4758.965 3402.535 4759.365 ;
        RECT 3406.785 4758.965 3407.385 4759.365 ;
      LAYER met4 ;
        RECT 3402.935 4613.000 3406.385 4758.965 ;
        RECT 3407.785 4613.000 3412.435 4759.270 ;
      LAYER met4 ;
        RECT 3412.835 4758.965 3413.435 4759.670 ;
      LAYER met4 ;
        RECT 3413.835 4613.000 3418.485 4759.270 ;
      LAYER met4 ;
        RECT 3418.885 4758.965 3419.485 4759.670 ;
      LAYER met4 ;
        RECT 3419.885 4613.000 3423.335 4759.270 ;
      LAYER met4 ;
        RECT 3423.735 4758.965 3424.335 4759.670 ;
      LAYER met4 ;
        RECT 3424.735 4613.000 3428.185 4759.270 ;
      LAYER met4 ;
        RECT 3428.585 4758.965 3429.185 4759.670 ;
      LAYER met4 ;
        RECT 3429.585 4613.000 3434.235 4759.270 ;
      LAYER met4 ;
        RECT 3434.635 4758.965 3435.335 4759.670 ;
      LAYER met4 ;
        RECT 3435.735 4613.000 3436.065 5007.575 ;
      LAYER met4 ;
        RECT 3436.465 5005.955 3440.725 5007.975 ;
        RECT 3436.465 5005.275 3439.245 5005.955 ;
      LAYER met4 ;
        RECT 3436.365 4613.000 3439.345 5004.875 ;
        RECT 3439.645 4984.000 3440.825 5005.555 ;
      LAYER met4 ;
        RECT 3439.645 4833.000 3440.825 4984.000 ;
      LAYER met4 ;
        RECT 3439.645 4831.730 3440.825 4833.000 ;
      LAYER met4 ;
        RECT 3439.745 4759.670 3440.725 4831.330 ;
      LAYER met4 ;
        RECT 3439.645 4758.000 3440.825 4759.270 ;
      LAYER met4 ;
        RECT 3439.645 4613.000 3440.825 4758.000 ;
      LAYER met4 ;
        RECT 3441.125 4613.000 3444.105 5010.910 ;
        RECT 3444.405 4613.000 3444.735 5011.175 ;
      LAYER met4 ;
        RECT 3445.135 4986.255 3588.000 5011.575 ;
        RECT 3445.135 4985.670 3457.635 4986.255 ;
        RECT 3445.135 4985.255 3445.835 4985.670 ;
        RECT 3445.135 4833.000 3445.835 4984.000 ;
        RECT 3445.135 4831.330 3445.835 4832.035 ;
      LAYER met4 ;
        RECT 3446.235 4831.730 3450.685 4985.270 ;
      LAYER met4 ;
        RECT 3451.085 4985.255 3451.685 4985.670 ;
        RECT 3451.085 4833.000 3451.685 4984.000 ;
        RECT 3451.085 4831.330 3451.685 4832.035 ;
      LAYER met4 ;
        RECT 3452.085 4831.730 3456.535 4985.270 ;
      LAYER met4 ;
        RECT 3456.935 4985.255 3457.635 4985.670 ;
        RECT 3456.935 4833.000 3457.635 4984.000 ;
        RECT 3456.935 4831.330 3457.635 4832.035 ;
      LAYER met4 ;
        RECT 3458.035 4831.730 3483.000 4985.855 ;
      LAYER met4 ;
        RECT 3483.400 4985.670 3588.000 4986.255 ;
        RECT 3483.400 4985.255 3563.385 4985.670 ;
      LAYER met4 ;
        RECT 3563.785 4984.000 3588.000 4985.270 ;
      LAYER met4 ;
        RECT 3483.400 4833.000 3588.000 4984.000 ;
        RECT 3483.400 4831.330 3563.385 4832.035 ;
      LAYER met4 ;
        RECT 3563.785 4831.730 3588.000 4833.000 ;
      LAYER met4 ;
        RECT 3445.135 4759.670 3588.000 4831.330 ;
        RECT 3445.135 4758.965 3445.835 4759.670 ;
        RECT 3445.135 4613.000 3445.835 4758.000 ;
      LAYER met4 ;
        RECT 3446.235 4613.000 3450.685 4759.270 ;
      LAYER met4 ;
        RECT 3451.085 4758.965 3451.685 4759.670 ;
        RECT 3451.085 4613.000 3451.685 4758.000 ;
      LAYER met4 ;
        RECT 3452.085 4613.000 3456.535 4759.270 ;
      LAYER met4 ;
        RECT 3456.935 4758.965 3457.635 4759.670 ;
        RECT 3456.935 4613.000 3457.635 4758.000 ;
      LAYER met4 ;
        RECT 3458.035 4613.000 3483.000 4759.270 ;
      LAYER met4 ;
        RECT 3483.400 4758.965 3563.385 4759.670 ;
      LAYER met4 ;
        RECT 3563.785 4758.000 3588.000 4759.270 ;
      LAYER met4 ;
        RECT 3483.400 4613.000 3588.000 4758.000 ;
        RECT 0.000 4424.000 104.600 4560.000 ;
      LAYER met4 ;
        RECT 0.000 4422.730 24.215 4424.000 ;
      LAYER met4 ;
        RECT 24.615 4422.330 104.600 4423.035 ;
      LAYER met4 ;
        RECT 105.000 4422.730 129.965 4560.000 ;
      LAYER met4 ;
        RECT 130.365 4424.000 131.065 4560.000 ;
        RECT 130.365 4422.330 131.065 4423.035 ;
      LAYER met4 ;
        RECT 131.465 4422.730 135.915 4560.000 ;
      LAYER met4 ;
        RECT 136.315 4424.000 136.915 4560.000 ;
        RECT 136.315 4422.330 136.915 4423.035 ;
      LAYER met4 ;
        RECT 137.315 4422.730 141.765 4560.000 ;
      LAYER met4 ;
        RECT 142.165 4424.000 142.865 4560.000 ;
        RECT 142.165 4422.330 142.865 4423.035 ;
        RECT 0.000 4350.670 142.865 4422.330 ;
      LAYER met4 ;
        RECT 0.000 4349.000 24.215 4350.270 ;
      LAYER met4 ;
        RECT 24.615 4349.965 104.600 4350.670 ;
        RECT 0.000 4213.000 104.600 4349.000 ;
      LAYER met4 ;
        RECT 0.000 4211.730 24.215 4213.000 ;
      LAYER met4 ;
        RECT 24.615 4211.330 104.600 4212.035 ;
      LAYER met4 ;
        RECT 105.000 4211.730 129.965 4350.270 ;
      LAYER met4 ;
        RECT 130.365 4349.965 131.065 4350.670 ;
        RECT 130.365 4213.000 131.065 4349.000 ;
        RECT 130.365 4211.330 131.065 4212.035 ;
      LAYER met4 ;
        RECT 131.465 4211.730 135.915 4350.270 ;
      LAYER met4 ;
        RECT 136.315 4349.965 136.915 4350.670 ;
        RECT 136.315 4213.000 136.915 4349.000 ;
        RECT 136.315 4211.330 136.915 4212.035 ;
      LAYER met4 ;
        RECT 137.315 4211.730 141.765 4350.270 ;
      LAYER met4 ;
        RECT 142.165 4349.965 142.865 4350.670 ;
        RECT 142.165 4213.000 142.865 4349.000 ;
        RECT 142.165 4211.330 142.865 4212.035 ;
      LAYER met4 ;
        RECT 143.265 4211.730 143.595 4560.000 ;
      LAYER met4 ;
        RECT 0.000 4139.670 143.495 4211.330 ;
      LAYER met4 ;
        RECT 0.000 4138.000 24.215 4139.270 ;
      LAYER met4 ;
        RECT 24.615 4138.965 104.600 4139.670 ;
        RECT 0.000 4002.000 104.600 4138.000 ;
      LAYER met4 ;
        RECT 0.000 4000.730 24.215 4002.000 ;
      LAYER met4 ;
        RECT 24.615 4000.330 104.600 4000.970 ;
      LAYER met4 ;
        RECT 105.000 4000.730 129.965 4139.270 ;
      LAYER met4 ;
        RECT 130.365 4138.965 131.065 4139.670 ;
        RECT 130.365 4002.000 131.065 4138.000 ;
        RECT 130.365 4000.330 131.065 4000.970 ;
      LAYER met4 ;
        RECT 131.465 4000.730 135.915 4139.270 ;
      LAYER met4 ;
        RECT 136.315 4138.965 136.915 4139.670 ;
        RECT 136.315 4002.000 136.915 4138.000 ;
        RECT 136.315 4000.330 136.915 4000.970 ;
      LAYER met4 ;
        RECT 137.315 4000.730 141.765 4139.270 ;
      LAYER met4 ;
        RECT 142.165 4138.965 142.865 4139.670 ;
        RECT 142.165 4002.000 142.865 4138.000 ;
        RECT 142.165 4000.330 142.865 4000.970 ;
        RECT 0.000 3968.690 142.865 4000.330 ;
      LAYER met4 ;
        RECT 143.265 3969.090 143.595 4139.270 ;
      LAYER met4 ;
        RECT 0.000 3960.360 143.495 3968.690 ;
      LAYER met4 ;
        RECT 143.895 3960.760 146.875 4560.000 ;
      LAYER met4 ;
        RECT 147.175 4424.000 148.355 4560.000 ;
      LAYER met4 ;
        RECT 147.175 4422.730 148.355 4424.000 ;
      LAYER met4 ;
        RECT 147.275 4350.670 148.255 4422.330 ;
      LAYER met4 ;
        RECT 147.175 4349.000 148.355 4350.270 ;
      LAYER met4 ;
        RECT 147.175 4213.000 148.355 4349.000 ;
      LAYER met4 ;
        RECT 147.175 4211.730 148.355 4213.000 ;
      LAYER met4 ;
        RECT 147.275 4139.670 148.255 4211.330 ;
      LAYER met4 ;
        RECT 147.175 4138.000 148.355 4139.270 ;
      LAYER met4 ;
        RECT 147.175 4002.000 148.355 4138.000 ;
      LAYER met4 ;
        RECT 147.175 4000.730 148.355 4002.000 ;
      LAYER met4 ;
        RECT 147.275 3976.065 148.255 4000.330 ;
      LAYER met4 ;
        RECT 148.655 3976.465 151.635 4560.000 ;
        RECT 151.935 4211.730 152.265 4560.000 ;
      LAYER met4 ;
        RECT 152.665 4422.330 153.365 4423.035 ;
      LAYER met4 ;
        RECT 153.765 4422.730 158.415 4560.000 ;
      LAYER met4 ;
        RECT 158.815 4422.330 159.415 4423.035 ;
      LAYER met4 ;
        RECT 159.815 4422.730 163.265 4560.000 ;
      LAYER met4 ;
        RECT 163.665 4422.330 164.265 4423.035 ;
      LAYER met4 ;
        RECT 164.665 4422.730 168.115 4560.000 ;
      LAYER met4 ;
        RECT 168.515 4422.330 169.115 4423.035 ;
      LAYER met4 ;
        RECT 169.515 4422.730 174.165 4560.000 ;
      LAYER met4 ;
        RECT 174.565 4422.330 175.165 4423.035 ;
      LAYER met4 ;
        RECT 175.565 4422.730 180.215 4560.000 ;
        RECT 181.615 4423.035 185.065 4560.000 ;
      LAYER met4 ;
        RECT 180.615 4422.635 181.215 4423.035 ;
        RECT 185.465 4422.635 186.065 4423.035 ;
      LAYER met4 ;
        RECT 186.465 4422.730 191.115 4560.000 ;
      LAYER met4 ;
        RECT 180.615 4422.330 186.065 4422.635 ;
        RECT 191.515 4422.330 192.115 4423.035 ;
      LAYER met4 ;
        RECT 192.515 4422.730 197.965 4560.000 ;
      LAYER met4 ;
        RECT 152.665 4350.670 197.965 4422.330 ;
        RECT 3388.535 4390.330 3389.635 4391.035 ;
      LAYER met4 ;
        RECT 3390.035 4390.730 3395.485 4538.000 ;
      LAYER met4 ;
        RECT 3395.885 4390.330 3396.485 4391.035 ;
      LAYER met4 ;
        RECT 3396.885 4390.730 3401.535 4538.000 ;
        RECT 3402.935 4391.035 3406.385 4538.000 ;
      LAYER met4 ;
        RECT 3401.935 4390.635 3402.535 4391.035 ;
        RECT 3406.785 4390.635 3407.385 4391.035 ;
      LAYER met4 ;
        RECT 3407.785 4390.730 3412.435 4538.000 ;
      LAYER met4 ;
        RECT 3401.935 4390.330 3407.385 4390.635 ;
        RECT 3412.835 4390.330 3413.435 4391.035 ;
      LAYER met4 ;
        RECT 3413.835 4390.730 3418.485 4538.000 ;
      LAYER met4 ;
        RECT 3418.885 4390.330 3419.485 4391.035 ;
      LAYER met4 ;
        RECT 3419.885 4390.730 3423.335 4538.000 ;
      LAYER met4 ;
        RECT 3423.735 4390.330 3424.335 4391.035 ;
      LAYER met4 ;
        RECT 3424.735 4390.730 3428.185 4538.000 ;
      LAYER met4 ;
        RECT 3428.585 4390.330 3429.185 4391.035 ;
      LAYER met4 ;
        RECT 3429.585 4390.730 3434.235 4538.000 ;
      LAYER met4 ;
        RECT 3434.635 4390.330 3435.335 4391.035 ;
        RECT 3388.535 4388.990 3435.335 4390.330 ;
      LAYER met4 ;
        RECT 3435.735 4389.390 3436.065 4538.000 ;
      LAYER met4 ;
        RECT 152.665 4349.965 153.365 4350.670 ;
        RECT 152.665 4211.330 153.365 4212.035 ;
      LAYER met4 ;
        RECT 153.765 4211.730 158.415 4350.270 ;
      LAYER met4 ;
        RECT 158.815 4349.965 159.415 4350.670 ;
        RECT 158.815 4211.330 159.415 4212.035 ;
      LAYER met4 ;
        RECT 159.815 4211.730 163.265 4350.270 ;
      LAYER met4 ;
        RECT 163.665 4349.965 164.265 4350.670 ;
        RECT 163.665 4211.330 164.265 4212.035 ;
      LAYER met4 ;
        RECT 164.665 4211.730 168.115 4350.270 ;
      LAYER met4 ;
        RECT 168.515 4349.965 169.115 4350.670 ;
        RECT 168.515 4211.330 169.115 4212.035 ;
      LAYER met4 ;
        RECT 169.515 4211.730 174.165 4350.270 ;
      LAYER met4 ;
        RECT 174.565 4349.965 175.165 4350.670 ;
        RECT 180.615 4350.365 186.065 4350.670 ;
        RECT 174.565 4211.330 175.165 4212.035 ;
      LAYER met4 ;
        RECT 175.565 4211.730 180.215 4350.270 ;
      LAYER met4 ;
        RECT 180.615 4349.965 181.215 4350.365 ;
        RECT 185.465 4349.965 186.065 4350.365 ;
      LAYER met4 ;
        RECT 181.615 4212.035 185.065 4349.965 ;
      LAYER met4 ;
        RECT 180.615 4211.635 181.215 4212.035 ;
        RECT 185.465 4211.635 186.065 4212.035 ;
      LAYER met4 ;
        RECT 186.465 4211.730 191.115 4350.270 ;
      LAYER met4 ;
        RECT 191.515 4349.965 192.115 4350.670 ;
        RECT 180.615 4211.330 186.065 4211.635 ;
        RECT 191.515 4211.330 192.115 4212.035 ;
      LAYER met4 ;
        RECT 192.515 4211.730 197.965 4350.270 ;
      LAYER met4 ;
        RECT 3388.535 4345.310 3435.965 4388.990 ;
        RECT 3388.535 4313.670 3435.335 4345.310 ;
        RECT 3388.535 4313.030 3389.635 4313.670 ;
        RECT 152.035 4139.670 197.965 4211.330 ;
      LAYER met4 ;
        RECT 3390.035 4165.730 3395.485 4313.270 ;
      LAYER met4 ;
        RECT 3395.885 4313.030 3396.485 4313.670 ;
        RECT 3401.935 4313.430 3407.385 4313.670 ;
        RECT 3395.885 4165.330 3396.485 4166.035 ;
      LAYER met4 ;
        RECT 3396.885 4165.730 3401.535 4313.270 ;
      LAYER met4 ;
        RECT 3401.935 4313.030 3402.535 4313.430 ;
        RECT 3406.785 4313.030 3407.385 4313.430 ;
      LAYER met4 ;
        RECT 3402.935 4166.035 3406.385 4313.030 ;
      LAYER met4 ;
        RECT 3401.935 4165.635 3402.535 4166.035 ;
        RECT 3406.785 4165.635 3407.385 4166.035 ;
      LAYER met4 ;
        RECT 3407.785 4165.730 3412.435 4313.270 ;
      LAYER met4 ;
        RECT 3412.835 4313.030 3413.435 4313.670 ;
        RECT 3401.935 4165.330 3407.385 4165.635 ;
        RECT 3412.835 4165.330 3413.435 4166.035 ;
      LAYER met4 ;
        RECT 3413.835 4165.730 3418.485 4313.270 ;
      LAYER met4 ;
        RECT 3418.885 4313.030 3419.485 4313.670 ;
        RECT 3418.885 4165.330 3419.485 4166.035 ;
      LAYER met4 ;
        RECT 3419.885 4165.730 3423.335 4313.270 ;
      LAYER met4 ;
        RECT 3423.735 4313.030 3424.335 4313.670 ;
        RECT 3423.735 4165.330 3424.335 4166.035 ;
      LAYER met4 ;
        RECT 3424.735 4165.730 3428.185 4313.270 ;
      LAYER met4 ;
        RECT 3428.585 4313.030 3429.185 4313.670 ;
        RECT 3428.585 4165.330 3429.185 4166.035 ;
      LAYER met4 ;
        RECT 3429.585 4165.730 3434.235 4313.270 ;
      LAYER met4 ;
        RECT 3434.635 4313.030 3435.335 4313.670 ;
        RECT 3434.635 4165.330 3435.335 4166.035 ;
        RECT 147.275 3974.545 151.535 3976.065 ;
        RECT 147.275 3960.360 148.255 3974.545 ;
        RECT 0.000 3958.840 148.255 3960.360 ;
        RECT 0.000 3925.010 143.495 3958.840 ;
        RECT 0.000 3923.670 142.865 3925.010 ;
      LAYER met4 ;
        RECT 0.000 3922.000 24.215 3923.270 ;
      LAYER met4 ;
        RECT 24.615 3922.965 104.600 3923.670 ;
        RECT 0.000 3786.000 104.600 3922.000 ;
      LAYER met4 ;
        RECT 0.000 3784.730 24.215 3786.000 ;
      LAYER met4 ;
        RECT 24.615 3784.330 104.600 3784.970 ;
      LAYER met4 ;
        RECT 105.000 3784.730 129.965 3923.270 ;
      LAYER met4 ;
        RECT 130.365 3922.965 131.065 3923.670 ;
        RECT 130.365 3786.000 131.065 3922.000 ;
        RECT 130.365 3784.330 131.065 3784.970 ;
      LAYER met4 ;
        RECT 131.465 3784.730 135.915 3923.270 ;
      LAYER met4 ;
        RECT 136.315 3922.965 136.915 3923.670 ;
        RECT 136.315 3786.000 136.915 3922.000 ;
        RECT 136.315 3784.330 136.915 3784.970 ;
      LAYER met4 ;
        RECT 137.315 3784.730 141.765 3923.270 ;
      LAYER met4 ;
        RECT 142.165 3922.965 142.865 3923.670 ;
        RECT 142.165 3786.000 142.865 3922.000 ;
        RECT 142.165 3784.330 142.865 3784.970 ;
        RECT 0.000 3752.690 142.865 3784.330 ;
      LAYER met4 ;
        RECT 143.265 3753.090 143.595 3924.610 ;
      LAYER met4 ;
        RECT 0.000 3744.360 143.495 3752.690 ;
      LAYER met4 ;
        RECT 143.895 3744.760 146.875 3958.440 ;
      LAYER met4 ;
        RECT 147.275 3923.670 148.255 3958.840 ;
      LAYER met4 ;
        RECT 147.175 3922.000 148.355 3923.270 ;
      LAYER met4 ;
        RECT 147.175 3786.000 148.355 3922.000 ;
      LAYER met4 ;
        RECT 147.175 3784.730 148.355 3786.000 ;
      LAYER met4 ;
        RECT 147.275 3760.065 148.255 3784.330 ;
      LAYER met4 ;
        RECT 148.655 3760.465 151.635 3974.145 ;
        RECT 151.935 3969.090 152.265 4139.270 ;
      LAYER met4 ;
        RECT 152.665 4138.965 153.365 4139.670 ;
        RECT 152.665 4000.330 153.365 4000.970 ;
      LAYER met4 ;
        RECT 153.765 4000.730 158.415 4139.270 ;
      LAYER met4 ;
        RECT 158.815 4138.965 159.415 4139.670 ;
        RECT 158.815 4000.330 159.415 4000.970 ;
      LAYER met4 ;
        RECT 159.815 4000.730 163.265 4139.270 ;
      LAYER met4 ;
        RECT 163.665 4138.965 164.265 4139.670 ;
        RECT 163.665 4000.330 164.265 4000.970 ;
      LAYER met4 ;
        RECT 164.665 4000.730 168.115 4139.270 ;
      LAYER met4 ;
        RECT 168.515 4138.965 169.115 4139.670 ;
        RECT 168.515 4000.330 169.115 4000.970 ;
      LAYER met4 ;
        RECT 169.515 4000.730 174.165 4139.270 ;
      LAYER met4 ;
        RECT 174.565 4138.965 175.165 4139.670 ;
        RECT 180.615 4139.365 186.065 4139.670 ;
        RECT 174.565 4000.330 175.165 4000.970 ;
      LAYER met4 ;
        RECT 175.565 4000.730 180.215 4139.270 ;
      LAYER met4 ;
        RECT 180.615 4138.965 181.215 4139.365 ;
        RECT 185.465 4138.965 186.065 4139.365 ;
      LAYER met4 ;
        RECT 181.615 4000.970 185.065 4138.965 ;
      LAYER met4 ;
        RECT 180.615 4000.570 181.215 4000.970 ;
        RECT 185.465 4000.570 186.065 4000.970 ;
      LAYER met4 ;
        RECT 186.465 4000.730 191.115 4139.270 ;
      LAYER met4 ;
        RECT 191.515 4138.965 192.115 4139.670 ;
        RECT 180.615 4000.330 186.065 4000.570 ;
        RECT 191.515 4000.330 192.115 4000.970 ;
      LAYER met4 ;
        RECT 192.515 4000.730 197.965 4139.270 ;
      LAYER met4 ;
        RECT 3390.035 4093.670 3435.335 4165.330 ;
        RECT 198.365 4000.330 199.465 4000.970 ;
        RECT 152.665 3968.690 199.465 4000.330 ;
        RECT 152.035 3925.010 199.465 3968.690 ;
        RECT 147.275 3758.545 151.535 3760.065 ;
        RECT 147.275 3744.360 148.255 3758.545 ;
        RECT 0.000 3742.840 148.255 3744.360 ;
        RECT 0.000 3709.010 143.495 3742.840 ;
        RECT 0.000 3707.670 142.865 3709.010 ;
      LAYER met4 ;
        RECT 0.000 3706.000 24.215 3707.270 ;
      LAYER met4 ;
        RECT 24.615 3706.965 104.600 3707.670 ;
        RECT 0.000 3570.000 104.600 3706.000 ;
      LAYER met4 ;
        RECT 0.000 3568.730 24.215 3570.000 ;
      LAYER met4 ;
        RECT 24.615 3568.330 104.600 3568.970 ;
      LAYER met4 ;
        RECT 105.000 3568.730 129.965 3707.270 ;
      LAYER met4 ;
        RECT 130.365 3706.965 131.065 3707.670 ;
        RECT 130.365 3570.000 131.065 3706.000 ;
        RECT 130.365 3568.330 131.065 3568.970 ;
      LAYER met4 ;
        RECT 131.465 3568.730 135.915 3707.270 ;
      LAYER met4 ;
        RECT 136.315 3706.965 136.915 3707.670 ;
        RECT 136.315 3570.000 136.915 3706.000 ;
        RECT 136.315 3568.330 136.915 3568.970 ;
      LAYER met4 ;
        RECT 137.315 3568.730 141.765 3707.270 ;
      LAYER met4 ;
        RECT 142.165 3706.965 142.865 3707.670 ;
        RECT 142.165 3570.000 142.865 3706.000 ;
        RECT 142.165 3568.330 142.865 3568.970 ;
        RECT 0.000 3536.690 142.865 3568.330 ;
      LAYER met4 ;
        RECT 143.265 3537.090 143.595 3708.610 ;
      LAYER met4 ;
        RECT 0.000 3528.360 143.495 3536.690 ;
      LAYER met4 ;
        RECT 143.895 3528.760 146.875 3742.440 ;
      LAYER met4 ;
        RECT 147.275 3707.670 148.255 3742.840 ;
      LAYER met4 ;
        RECT 147.175 3706.000 148.355 3707.270 ;
      LAYER met4 ;
        RECT 147.175 3570.000 148.355 3706.000 ;
      LAYER met4 ;
        RECT 147.175 3568.730 148.355 3570.000 ;
      LAYER met4 ;
        RECT 147.275 3544.065 148.255 3568.330 ;
      LAYER met4 ;
        RECT 148.655 3544.465 151.635 3758.145 ;
        RECT 151.935 3753.090 152.265 3924.610 ;
      LAYER met4 ;
        RECT 152.665 3923.670 199.465 3925.010 ;
        RECT 152.665 3922.965 153.365 3923.670 ;
        RECT 152.665 3784.330 153.365 3784.970 ;
      LAYER met4 ;
        RECT 153.765 3784.730 158.415 3923.270 ;
      LAYER met4 ;
        RECT 158.815 3922.965 159.415 3923.670 ;
        RECT 158.815 3784.330 159.415 3784.970 ;
      LAYER met4 ;
        RECT 159.815 3784.730 163.265 3923.270 ;
      LAYER met4 ;
        RECT 163.665 3922.965 164.265 3923.670 ;
        RECT 163.665 3784.330 164.265 3784.970 ;
      LAYER met4 ;
        RECT 164.665 3784.730 168.115 3923.270 ;
      LAYER met4 ;
        RECT 168.515 3922.965 169.115 3923.670 ;
        RECT 168.515 3784.330 169.115 3784.970 ;
      LAYER met4 ;
        RECT 169.515 3784.730 174.165 3923.270 ;
      LAYER met4 ;
        RECT 174.565 3922.965 175.165 3923.670 ;
        RECT 180.615 3923.365 186.065 3923.670 ;
        RECT 174.565 3784.330 175.165 3784.970 ;
      LAYER met4 ;
        RECT 175.565 3784.730 180.215 3923.270 ;
      LAYER met4 ;
        RECT 180.615 3922.965 181.215 3923.365 ;
        RECT 185.465 3922.965 186.065 3923.365 ;
      LAYER met4 ;
        RECT 181.615 3784.970 185.065 3922.965 ;
      LAYER met4 ;
        RECT 180.615 3784.570 181.215 3784.970 ;
        RECT 185.465 3784.570 186.065 3784.970 ;
      LAYER met4 ;
        RECT 186.465 3784.730 191.115 3923.270 ;
      LAYER met4 ;
        RECT 191.515 3922.965 192.115 3923.670 ;
        RECT 180.615 3784.330 186.065 3784.570 ;
        RECT 191.515 3784.330 192.115 3784.970 ;
      LAYER met4 ;
        RECT 192.515 3784.730 197.965 3923.270 ;
      LAYER met4 ;
        RECT 198.365 3922.965 199.465 3923.670 ;
        RECT 3388.535 3944.330 3389.635 3945.035 ;
      LAYER met4 ;
        RECT 3390.035 3944.730 3395.485 4093.270 ;
      LAYER met4 ;
        RECT 3395.885 4092.965 3396.485 4093.670 ;
        RECT 3401.935 4093.365 3407.385 4093.670 ;
        RECT 3395.885 3944.330 3396.485 3945.035 ;
      LAYER met4 ;
        RECT 3396.885 3944.730 3401.535 4093.270 ;
      LAYER met4 ;
        RECT 3401.935 4092.965 3402.535 4093.365 ;
        RECT 3406.785 4092.965 3407.385 4093.365 ;
      LAYER met4 ;
        RECT 3402.935 3945.035 3406.385 4092.965 ;
      LAYER met4 ;
        RECT 3401.935 3944.635 3402.535 3945.035 ;
        RECT 3406.785 3944.635 3407.385 3945.035 ;
      LAYER met4 ;
        RECT 3407.785 3944.730 3412.435 4093.270 ;
      LAYER met4 ;
        RECT 3412.835 4092.965 3413.435 4093.670 ;
        RECT 3401.935 3944.330 3407.385 3944.635 ;
        RECT 3412.835 3944.330 3413.435 3945.035 ;
      LAYER met4 ;
        RECT 3413.835 3944.730 3418.485 4093.270 ;
      LAYER met4 ;
        RECT 3418.885 4092.965 3419.485 4093.670 ;
        RECT 3418.885 3944.330 3419.485 3945.035 ;
      LAYER met4 ;
        RECT 3419.885 3944.730 3423.335 4093.270 ;
      LAYER met4 ;
        RECT 3423.735 4092.965 3424.335 4093.670 ;
        RECT 3423.735 3944.330 3424.335 3945.035 ;
      LAYER met4 ;
        RECT 3424.735 3944.730 3428.185 4093.270 ;
      LAYER met4 ;
        RECT 3428.585 4092.965 3429.185 4093.670 ;
        RECT 3428.585 3944.330 3429.185 3945.035 ;
      LAYER met4 ;
        RECT 3429.585 3944.730 3434.235 4093.270 ;
      LAYER met4 ;
        RECT 3434.635 4092.965 3435.335 4093.670 ;
        RECT 3434.635 3944.330 3435.335 3945.035 ;
        RECT 3388.535 3942.990 3435.335 3944.330 ;
      LAYER met4 ;
        RECT 3435.735 3943.390 3436.065 4344.910 ;
        RECT 3436.365 4339.855 3439.345 4538.000 ;
      LAYER met4 ;
        RECT 3439.645 4392.000 3440.825 4538.000 ;
      LAYER met4 ;
        RECT 3439.645 4390.730 3440.825 4392.000 ;
      LAYER met4 ;
        RECT 3439.745 4355.160 3440.725 4390.330 ;
      LAYER met4 ;
        RECT 3441.125 4355.560 3444.105 4538.000 ;
        RECT 3444.405 4389.390 3444.735 4538.000 ;
      LAYER met4 ;
        RECT 3445.135 4392.000 3445.835 4538.000 ;
        RECT 3445.135 4390.330 3445.835 4391.035 ;
      LAYER met4 ;
        RECT 3446.235 4390.730 3450.685 4538.000 ;
      LAYER met4 ;
        RECT 3451.085 4392.000 3451.685 4538.000 ;
        RECT 3451.085 4390.330 3451.685 4391.035 ;
      LAYER met4 ;
        RECT 3452.085 4390.730 3456.535 4538.000 ;
      LAYER met4 ;
        RECT 3456.935 4392.000 3457.635 4538.000 ;
        RECT 3456.935 4390.330 3457.635 4391.035 ;
      LAYER met4 ;
        RECT 3458.035 4390.730 3483.000 4538.000 ;
      LAYER met4 ;
        RECT 3483.400 4392.000 3588.000 4538.000 ;
        RECT 3483.400 4390.330 3563.385 4391.035 ;
      LAYER met4 ;
        RECT 3563.785 4390.730 3588.000 4392.000 ;
      LAYER met4 ;
        RECT 3445.135 4388.990 3588.000 4390.330 ;
        RECT 3444.505 4355.160 3588.000 4388.990 ;
        RECT 3439.745 4353.640 3588.000 4355.160 ;
        RECT 3439.745 4339.455 3440.725 4353.640 ;
        RECT 3436.465 4337.935 3440.725 4339.455 ;
        RECT 3388.535 3899.310 3435.965 3942.990 ;
        RECT 3388.535 3867.670 3435.335 3899.310 ;
        RECT 3388.535 3867.030 3389.635 3867.670 ;
        RECT 198.365 3784.330 199.465 3784.970 ;
        RECT 152.665 3752.690 199.465 3784.330 ;
        RECT 152.035 3709.010 199.465 3752.690 ;
        RECT 147.275 3542.545 151.535 3544.065 ;
        RECT 147.275 3528.360 148.255 3542.545 ;
        RECT 0.000 3526.840 148.255 3528.360 ;
        RECT 0.000 3493.010 143.495 3526.840 ;
        RECT 0.000 3491.670 142.865 3493.010 ;
      LAYER met4 ;
        RECT 0.000 3490.000 24.215 3491.270 ;
      LAYER met4 ;
        RECT 24.615 3490.965 104.600 3491.670 ;
        RECT 0.000 3354.000 104.600 3490.000 ;
      LAYER met4 ;
        RECT 0.000 3352.730 24.215 3354.000 ;
      LAYER met4 ;
        RECT 24.615 3352.330 104.600 3352.970 ;
      LAYER met4 ;
        RECT 105.000 3352.730 129.965 3491.270 ;
      LAYER met4 ;
        RECT 130.365 3490.965 131.065 3491.670 ;
        RECT 130.365 3354.000 131.065 3490.000 ;
        RECT 130.365 3352.330 131.065 3352.970 ;
      LAYER met4 ;
        RECT 131.465 3352.730 135.915 3491.270 ;
      LAYER met4 ;
        RECT 136.315 3490.965 136.915 3491.670 ;
        RECT 136.315 3354.000 136.915 3490.000 ;
        RECT 136.315 3352.330 136.915 3352.970 ;
      LAYER met4 ;
        RECT 137.315 3352.730 141.765 3491.270 ;
      LAYER met4 ;
        RECT 142.165 3490.965 142.865 3491.670 ;
        RECT 142.165 3354.000 142.865 3490.000 ;
        RECT 142.165 3352.330 142.865 3352.970 ;
        RECT 0.000 3320.690 142.865 3352.330 ;
      LAYER met4 ;
        RECT 143.265 3321.090 143.595 3492.610 ;
      LAYER met4 ;
        RECT 0.000 3312.360 143.495 3320.690 ;
      LAYER met4 ;
        RECT 143.895 3312.760 146.875 3526.440 ;
      LAYER met4 ;
        RECT 147.275 3491.670 148.255 3526.840 ;
      LAYER met4 ;
        RECT 147.175 3490.000 148.355 3491.270 ;
      LAYER met4 ;
        RECT 147.175 3354.000 148.355 3490.000 ;
      LAYER met4 ;
        RECT 147.175 3352.730 148.355 3354.000 ;
      LAYER met4 ;
        RECT 147.275 3328.065 148.255 3352.330 ;
      LAYER met4 ;
        RECT 148.655 3328.465 151.635 3542.145 ;
        RECT 151.935 3537.090 152.265 3708.610 ;
      LAYER met4 ;
        RECT 152.665 3707.670 199.465 3709.010 ;
        RECT 152.665 3706.965 153.365 3707.670 ;
        RECT 152.665 3568.330 153.365 3568.970 ;
      LAYER met4 ;
        RECT 153.765 3568.730 158.415 3707.270 ;
      LAYER met4 ;
        RECT 158.815 3706.965 159.415 3707.670 ;
        RECT 158.815 3568.330 159.415 3568.970 ;
      LAYER met4 ;
        RECT 159.815 3568.730 163.265 3707.270 ;
      LAYER met4 ;
        RECT 163.665 3706.965 164.265 3707.670 ;
        RECT 163.665 3568.330 164.265 3568.970 ;
      LAYER met4 ;
        RECT 164.665 3568.730 168.115 3707.270 ;
      LAYER met4 ;
        RECT 168.515 3706.965 169.115 3707.670 ;
        RECT 168.515 3568.330 169.115 3568.970 ;
      LAYER met4 ;
        RECT 169.515 3568.730 174.165 3707.270 ;
      LAYER met4 ;
        RECT 174.565 3706.965 175.165 3707.670 ;
        RECT 180.615 3707.365 186.065 3707.670 ;
        RECT 174.565 3568.330 175.165 3568.970 ;
      LAYER met4 ;
        RECT 175.565 3568.730 180.215 3707.270 ;
      LAYER met4 ;
        RECT 180.615 3706.965 181.215 3707.365 ;
        RECT 185.465 3706.965 186.065 3707.365 ;
      LAYER met4 ;
        RECT 181.615 3568.970 185.065 3706.965 ;
      LAYER met4 ;
        RECT 180.615 3568.570 181.215 3568.970 ;
        RECT 185.465 3568.570 186.065 3568.970 ;
      LAYER met4 ;
        RECT 186.465 3568.730 191.115 3707.270 ;
      LAYER met4 ;
        RECT 191.515 3706.965 192.115 3707.670 ;
        RECT 180.615 3568.330 186.065 3568.570 ;
        RECT 191.515 3568.330 192.115 3568.970 ;
      LAYER met4 ;
        RECT 192.515 3568.730 197.965 3707.270 ;
      LAYER met4 ;
        RECT 198.365 3706.965 199.465 3707.670 ;
        RECT 3388.535 3719.330 3389.635 3720.035 ;
      LAYER met4 ;
        RECT 3390.035 3719.730 3395.485 3867.270 ;
      LAYER met4 ;
        RECT 3395.885 3867.030 3396.485 3867.670 ;
        RECT 3401.935 3867.430 3407.385 3867.670 ;
        RECT 3395.885 3719.330 3396.485 3720.035 ;
      LAYER met4 ;
        RECT 3396.885 3719.730 3401.535 3867.270 ;
      LAYER met4 ;
        RECT 3401.935 3867.030 3402.535 3867.430 ;
        RECT 3406.785 3867.030 3407.385 3867.430 ;
      LAYER met4 ;
        RECT 3402.935 3720.035 3406.385 3867.030 ;
      LAYER met4 ;
        RECT 3401.935 3719.635 3402.535 3720.035 ;
        RECT 3406.785 3719.635 3407.385 3720.035 ;
      LAYER met4 ;
        RECT 3407.785 3719.730 3412.435 3867.270 ;
      LAYER met4 ;
        RECT 3412.835 3867.030 3413.435 3867.670 ;
        RECT 3401.935 3719.330 3407.385 3719.635 ;
        RECT 3412.835 3719.330 3413.435 3720.035 ;
      LAYER met4 ;
        RECT 3413.835 3719.730 3418.485 3867.270 ;
      LAYER met4 ;
        RECT 3418.885 3867.030 3419.485 3867.670 ;
        RECT 3418.885 3719.330 3419.485 3720.035 ;
      LAYER met4 ;
        RECT 3419.885 3719.730 3423.335 3867.270 ;
      LAYER met4 ;
        RECT 3423.735 3867.030 3424.335 3867.670 ;
        RECT 3423.735 3719.330 3424.335 3720.035 ;
      LAYER met4 ;
        RECT 3424.735 3719.730 3428.185 3867.270 ;
      LAYER met4 ;
        RECT 3428.585 3867.030 3429.185 3867.670 ;
        RECT 3428.585 3719.330 3429.185 3720.035 ;
      LAYER met4 ;
        RECT 3429.585 3719.730 3434.235 3867.270 ;
      LAYER met4 ;
        RECT 3434.635 3867.030 3435.335 3867.670 ;
        RECT 3434.635 3719.330 3435.335 3720.035 ;
        RECT 3388.535 3717.990 3435.335 3719.330 ;
      LAYER met4 ;
        RECT 3435.735 3718.390 3436.065 3898.910 ;
        RECT 3436.365 3893.855 3439.345 4337.535 ;
      LAYER met4 ;
        RECT 3439.745 4313.670 3440.725 4337.935 ;
      LAYER met4 ;
        RECT 3439.645 4312.000 3440.825 4313.270 ;
      LAYER met4 ;
        RECT 3439.645 4167.000 3440.825 4312.000 ;
      LAYER met4 ;
        RECT 3439.645 4165.730 3440.825 4167.000 ;
      LAYER met4 ;
        RECT 3439.745 4093.670 3440.725 4165.330 ;
      LAYER met4 ;
        RECT 3439.645 4092.000 3440.825 4093.270 ;
      LAYER met4 ;
        RECT 3439.645 3946.000 3440.825 4092.000 ;
      LAYER met4 ;
        RECT 3439.645 3944.730 3440.825 3946.000 ;
      LAYER met4 ;
        RECT 3439.745 3909.160 3440.725 3944.330 ;
      LAYER met4 ;
        RECT 3441.125 3909.560 3444.105 4353.240 ;
      LAYER met4 ;
        RECT 3444.505 4345.310 3588.000 4353.640 ;
      LAYER met4 ;
        RECT 3444.405 3943.390 3444.735 4344.910 ;
      LAYER met4 ;
        RECT 3445.135 4313.670 3588.000 4345.310 ;
        RECT 3445.135 4313.030 3445.835 4313.670 ;
        RECT 3445.135 4167.000 3445.835 4312.000 ;
        RECT 3445.135 4165.330 3445.835 4166.035 ;
      LAYER met4 ;
        RECT 3446.235 4165.730 3450.685 4313.270 ;
      LAYER met4 ;
        RECT 3451.085 4313.030 3451.685 4313.670 ;
        RECT 3451.085 4167.000 3451.685 4312.000 ;
        RECT 3451.085 4165.330 3451.685 4166.035 ;
      LAYER met4 ;
        RECT 3452.085 4165.730 3456.535 4313.270 ;
      LAYER met4 ;
        RECT 3456.935 4313.030 3457.635 4313.670 ;
        RECT 3456.935 4167.000 3457.635 4312.000 ;
        RECT 3456.935 4165.330 3457.635 4166.035 ;
      LAYER met4 ;
        RECT 3458.035 4165.730 3483.000 4313.270 ;
      LAYER met4 ;
        RECT 3483.400 4313.030 3563.385 4313.670 ;
      LAYER met4 ;
        RECT 3563.785 4312.000 3588.000 4313.270 ;
      LAYER met4 ;
        RECT 3483.400 4167.000 3588.000 4312.000 ;
        RECT 3483.400 4165.330 3563.385 4166.035 ;
      LAYER met4 ;
        RECT 3563.785 4165.730 3588.000 4167.000 ;
      LAYER met4 ;
        RECT 3445.135 4093.670 3588.000 4165.330 ;
        RECT 3445.135 4092.965 3445.835 4093.670 ;
        RECT 3445.135 3946.000 3445.835 4092.000 ;
        RECT 3445.135 3944.330 3445.835 3945.035 ;
      LAYER met4 ;
        RECT 3446.235 3944.730 3450.685 4093.270 ;
      LAYER met4 ;
        RECT 3451.085 4092.965 3451.685 4093.670 ;
        RECT 3451.085 3946.000 3451.685 4092.000 ;
        RECT 3451.085 3944.330 3451.685 3945.035 ;
      LAYER met4 ;
        RECT 3452.085 3944.730 3456.535 4093.270 ;
      LAYER met4 ;
        RECT 3456.935 4092.965 3457.635 4093.670 ;
        RECT 3456.935 3946.000 3457.635 4092.000 ;
        RECT 3456.935 3944.330 3457.635 3945.035 ;
      LAYER met4 ;
        RECT 3458.035 3944.730 3483.000 4093.270 ;
      LAYER met4 ;
        RECT 3483.400 4092.965 3563.385 4093.670 ;
      LAYER met4 ;
        RECT 3563.785 4092.000 3588.000 4093.270 ;
      LAYER met4 ;
        RECT 3483.400 3946.000 3588.000 4092.000 ;
        RECT 3483.400 3944.330 3563.385 3945.035 ;
      LAYER met4 ;
        RECT 3563.785 3944.730 3588.000 3946.000 ;
      LAYER met4 ;
        RECT 3445.135 3942.990 3588.000 3944.330 ;
        RECT 3444.505 3909.160 3588.000 3942.990 ;
        RECT 3439.745 3907.640 3588.000 3909.160 ;
        RECT 3439.745 3893.455 3440.725 3907.640 ;
        RECT 3436.465 3891.935 3440.725 3893.455 ;
        RECT 3388.535 3674.310 3435.965 3717.990 ;
        RECT 3388.535 3642.670 3435.335 3674.310 ;
        RECT 3388.535 3642.030 3389.635 3642.670 ;
        RECT 198.365 3568.330 199.465 3568.970 ;
        RECT 152.665 3536.690 199.465 3568.330 ;
        RECT 152.035 3493.010 199.465 3536.690 ;
        RECT 147.275 3326.545 151.535 3328.065 ;
        RECT 147.275 3312.360 148.255 3326.545 ;
        RECT 0.000 3310.840 148.255 3312.360 ;
        RECT 0.000 3277.010 143.495 3310.840 ;
        RECT 0.000 3275.670 142.865 3277.010 ;
      LAYER met4 ;
        RECT 0.000 3274.000 24.215 3275.270 ;
      LAYER met4 ;
        RECT 24.615 3274.965 104.600 3275.670 ;
        RECT 0.000 3138.000 104.600 3274.000 ;
      LAYER met4 ;
        RECT 0.000 3136.730 24.215 3138.000 ;
      LAYER met4 ;
        RECT 24.615 3136.330 104.600 3136.970 ;
      LAYER met4 ;
        RECT 105.000 3136.730 129.965 3275.270 ;
      LAYER met4 ;
        RECT 130.365 3274.965 131.065 3275.670 ;
        RECT 130.365 3138.000 131.065 3274.000 ;
        RECT 130.365 3136.330 131.065 3136.970 ;
      LAYER met4 ;
        RECT 131.465 3136.730 135.915 3275.270 ;
      LAYER met4 ;
        RECT 136.315 3274.965 136.915 3275.670 ;
        RECT 136.315 3138.000 136.915 3274.000 ;
        RECT 136.315 3136.330 136.915 3136.970 ;
      LAYER met4 ;
        RECT 137.315 3136.730 141.765 3275.270 ;
      LAYER met4 ;
        RECT 142.165 3274.965 142.865 3275.670 ;
        RECT 142.165 3138.000 142.865 3274.000 ;
        RECT 142.165 3136.330 142.865 3136.970 ;
        RECT 0.000 3104.690 142.865 3136.330 ;
      LAYER met4 ;
        RECT 143.265 3105.090 143.595 3276.610 ;
      LAYER met4 ;
        RECT 0.000 3096.360 143.495 3104.690 ;
      LAYER met4 ;
        RECT 143.895 3096.760 146.875 3310.440 ;
      LAYER met4 ;
        RECT 147.275 3275.670 148.255 3310.840 ;
      LAYER met4 ;
        RECT 147.175 3274.000 148.355 3275.270 ;
      LAYER met4 ;
        RECT 147.175 3138.000 148.355 3274.000 ;
      LAYER met4 ;
        RECT 147.175 3136.730 148.355 3138.000 ;
      LAYER met4 ;
        RECT 147.275 3112.065 148.255 3136.330 ;
      LAYER met4 ;
        RECT 148.655 3112.465 151.635 3326.145 ;
        RECT 151.935 3321.090 152.265 3492.610 ;
      LAYER met4 ;
        RECT 152.665 3491.670 199.465 3493.010 ;
        RECT 152.665 3490.965 153.365 3491.670 ;
        RECT 152.665 3352.330 153.365 3352.970 ;
      LAYER met4 ;
        RECT 153.765 3352.730 158.415 3491.270 ;
      LAYER met4 ;
        RECT 158.815 3490.965 159.415 3491.670 ;
        RECT 158.815 3352.330 159.415 3352.970 ;
      LAYER met4 ;
        RECT 159.815 3352.730 163.265 3491.270 ;
      LAYER met4 ;
        RECT 163.665 3490.965 164.265 3491.670 ;
        RECT 163.665 3352.330 164.265 3352.970 ;
      LAYER met4 ;
        RECT 164.665 3352.730 168.115 3491.270 ;
      LAYER met4 ;
        RECT 168.515 3490.965 169.115 3491.670 ;
        RECT 168.515 3352.330 169.115 3352.970 ;
      LAYER met4 ;
        RECT 169.515 3352.730 174.165 3491.270 ;
      LAYER met4 ;
        RECT 174.565 3490.965 175.165 3491.670 ;
        RECT 180.615 3491.365 186.065 3491.670 ;
        RECT 174.565 3352.330 175.165 3352.970 ;
      LAYER met4 ;
        RECT 175.565 3352.730 180.215 3491.270 ;
      LAYER met4 ;
        RECT 180.615 3490.965 181.215 3491.365 ;
        RECT 185.465 3490.965 186.065 3491.365 ;
      LAYER met4 ;
        RECT 181.615 3352.970 185.065 3490.965 ;
      LAYER met4 ;
        RECT 180.615 3352.570 181.215 3352.970 ;
        RECT 185.465 3352.570 186.065 3352.970 ;
      LAYER met4 ;
        RECT 186.465 3352.730 191.115 3491.270 ;
      LAYER met4 ;
        RECT 191.515 3490.965 192.115 3491.670 ;
        RECT 180.615 3352.330 186.065 3352.570 ;
        RECT 191.515 3352.330 192.115 3352.970 ;
      LAYER met4 ;
        RECT 192.515 3352.730 197.965 3491.270 ;
      LAYER met4 ;
        RECT 198.365 3490.965 199.465 3491.670 ;
        RECT 3388.535 3494.330 3389.635 3495.035 ;
      LAYER met4 ;
        RECT 3390.035 3494.730 3395.485 3642.270 ;
      LAYER met4 ;
        RECT 3395.885 3642.030 3396.485 3642.670 ;
        RECT 3401.935 3642.430 3407.385 3642.670 ;
        RECT 3395.885 3494.330 3396.485 3495.035 ;
      LAYER met4 ;
        RECT 3396.885 3494.730 3401.535 3642.270 ;
      LAYER met4 ;
        RECT 3401.935 3642.030 3402.535 3642.430 ;
        RECT 3406.785 3642.030 3407.385 3642.430 ;
      LAYER met4 ;
        RECT 3402.935 3495.035 3406.385 3642.030 ;
      LAYER met4 ;
        RECT 3401.935 3494.635 3402.535 3495.035 ;
        RECT 3406.785 3494.635 3407.385 3495.035 ;
      LAYER met4 ;
        RECT 3407.785 3494.730 3412.435 3642.270 ;
      LAYER met4 ;
        RECT 3412.835 3642.030 3413.435 3642.670 ;
        RECT 3401.935 3494.330 3407.385 3494.635 ;
        RECT 3412.835 3494.330 3413.435 3495.035 ;
      LAYER met4 ;
        RECT 3413.835 3494.730 3418.485 3642.270 ;
      LAYER met4 ;
        RECT 3418.885 3642.030 3419.485 3642.670 ;
        RECT 3418.885 3494.330 3419.485 3495.035 ;
      LAYER met4 ;
        RECT 3419.885 3494.730 3423.335 3642.270 ;
      LAYER met4 ;
        RECT 3423.735 3642.030 3424.335 3642.670 ;
        RECT 3423.735 3494.330 3424.335 3495.035 ;
      LAYER met4 ;
        RECT 3424.735 3494.730 3428.185 3642.270 ;
      LAYER met4 ;
        RECT 3428.585 3642.030 3429.185 3642.670 ;
        RECT 3428.585 3494.330 3429.185 3495.035 ;
      LAYER met4 ;
        RECT 3429.585 3494.730 3434.235 3642.270 ;
      LAYER met4 ;
        RECT 3434.635 3642.030 3435.335 3642.670 ;
        RECT 3434.635 3494.330 3435.335 3495.035 ;
        RECT 3388.535 3492.990 3435.335 3494.330 ;
      LAYER met4 ;
        RECT 3435.735 3493.390 3436.065 3673.910 ;
        RECT 3436.365 3668.855 3439.345 3891.535 ;
      LAYER met4 ;
        RECT 3439.745 3867.670 3440.725 3891.935 ;
      LAYER met4 ;
        RECT 3439.645 3866.000 3440.825 3867.270 ;
      LAYER met4 ;
        RECT 3439.645 3721.000 3440.825 3866.000 ;
      LAYER met4 ;
        RECT 3439.645 3719.730 3440.825 3721.000 ;
      LAYER met4 ;
        RECT 3439.745 3684.160 3440.725 3719.330 ;
      LAYER met4 ;
        RECT 3441.125 3684.560 3444.105 3907.240 ;
      LAYER met4 ;
        RECT 3444.505 3899.310 3588.000 3907.640 ;
      LAYER met4 ;
        RECT 3444.405 3718.390 3444.735 3898.910 ;
      LAYER met4 ;
        RECT 3445.135 3867.670 3588.000 3899.310 ;
        RECT 3445.135 3867.030 3445.835 3867.670 ;
        RECT 3445.135 3721.000 3445.835 3866.000 ;
        RECT 3445.135 3719.330 3445.835 3720.035 ;
      LAYER met4 ;
        RECT 3446.235 3719.730 3450.685 3867.270 ;
      LAYER met4 ;
        RECT 3451.085 3867.030 3451.685 3867.670 ;
        RECT 3451.085 3721.000 3451.685 3866.000 ;
        RECT 3451.085 3719.330 3451.685 3720.035 ;
      LAYER met4 ;
        RECT 3452.085 3719.730 3456.535 3867.270 ;
      LAYER met4 ;
        RECT 3456.935 3867.030 3457.635 3867.670 ;
        RECT 3456.935 3721.000 3457.635 3866.000 ;
        RECT 3456.935 3719.330 3457.635 3720.035 ;
      LAYER met4 ;
        RECT 3458.035 3719.730 3483.000 3867.270 ;
      LAYER met4 ;
        RECT 3483.400 3867.030 3563.385 3867.670 ;
      LAYER met4 ;
        RECT 3563.785 3866.000 3588.000 3867.270 ;
      LAYER met4 ;
        RECT 3483.400 3721.000 3588.000 3866.000 ;
        RECT 3483.400 3719.330 3563.385 3720.035 ;
      LAYER met4 ;
        RECT 3563.785 3719.730 3588.000 3721.000 ;
      LAYER met4 ;
        RECT 3445.135 3717.990 3588.000 3719.330 ;
        RECT 3444.505 3684.160 3588.000 3717.990 ;
        RECT 3439.745 3682.640 3588.000 3684.160 ;
        RECT 3439.745 3668.455 3440.725 3682.640 ;
        RECT 3436.465 3666.935 3440.725 3668.455 ;
        RECT 3388.535 3449.310 3435.965 3492.990 ;
        RECT 3388.535 3417.670 3435.335 3449.310 ;
        RECT 3388.535 3417.030 3389.635 3417.670 ;
        RECT 198.365 3352.330 199.465 3352.970 ;
        RECT 152.665 3320.690 199.465 3352.330 ;
        RECT 152.035 3277.010 199.465 3320.690 ;
        RECT 147.275 3110.545 151.535 3112.065 ;
        RECT 147.275 3096.360 148.255 3110.545 ;
        RECT 0.000 3094.840 148.255 3096.360 ;
        RECT 0.000 3061.010 143.495 3094.840 ;
        RECT 0.000 3059.670 142.865 3061.010 ;
      LAYER met4 ;
        RECT 0.000 3058.000 24.215 3059.270 ;
      LAYER met4 ;
        RECT 24.615 3058.965 104.600 3059.670 ;
        RECT 0.000 2922.000 104.600 3058.000 ;
      LAYER met4 ;
        RECT 0.000 2920.730 24.215 2922.000 ;
      LAYER met4 ;
        RECT 24.615 2920.330 104.600 2920.970 ;
      LAYER met4 ;
        RECT 105.000 2920.730 129.965 3059.270 ;
      LAYER met4 ;
        RECT 130.365 3058.965 131.065 3059.670 ;
        RECT 130.365 2922.000 131.065 3058.000 ;
        RECT 130.365 2920.330 131.065 2920.970 ;
      LAYER met4 ;
        RECT 131.465 2920.730 135.915 3059.270 ;
      LAYER met4 ;
        RECT 136.315 3058.965 136.915 3059.670 ;
        RECT 136.315 2922.000 136.915 3058.000 ;
        RECT 136.315 2920.330 136.915 2920.970 ;
      LAYER met4 ;
        RECT 137.315 2920.730 141.765 3059.270 ;
      LAYER met4 ;
        RECT 142.165 3058.965 142.865 3059.670 ;
        RECT 142.165 2922.000 142.865 3058.000 ;
        RECT 142.165 2920.330 142.865 2920.970 ;
        RECT 0.000 2888.690 142.865 2920.330 ;
      LAYER met4 ;
        RECT 143.265 2889.090 143.595 3060.610 ;
      LAYER met4 ;
        RECT 0.000 2880.360 143.495 2888.690 ;
      LAYER met4 ;
        RECT 143.895 2880.760 146.875 3094.440 ;
      LAYER met4 ;
        RECT 147.275 3059.670 148.255 3094.840 ;
      LAYER met4 ;
        RECT 147.175 3058.000 148.355 3059.270 ;
      LAYER met4 ;
        RECT 147.175 2922.000 148.355 3058.000 ;
      LAYER met4 ;
        RECT 147.175 2920.730 148.355 2922.000 ;
      LAYER met4 ;
        RECT 147.275 2896.065 148.255 2920.330 ;
      LAYER met4 ;
        RECT 148.655 2896.465 151.635 3110.145 ;
        RECT 151.935 3105.090 152.265 3276.610 ;
      LAYER met4 ;
        RECT 152.665 3275.670 199.465 3277.010 ;
        RECT 152.665 3274.965 153.365 3275.670 ;
        RECT 152.665 3136.330 153.365 3136.970 ;
      LAYER met4 ;
        RECT 153.765 3136.730 158.415 3275.270 ;
      LAYER met4 ;
        RECT 158.815 3274.965 159.415 3275.670 ;
        RECT 158.815 3136.330 159.415 3136.970 ;
      LAYER met4 ;
        RECT 159.815 3136.730 163.265 3275.270 ;
      LAYER met4 ;
        RECT 163.665 3274.965 164.265 3275.670 ;
        RECT 163.665 3136.330 164.265 3136.970 ;
      LAYER met4 ;
        RECT 164.665 3136.730 168.115 3275.270 ;
      LAYER met4 ;
        RECT 168.515 3274.965 169.115 3275.670 ;
        RECT 168.515 3136.330 169.115 3136.970 ;
      LAYER met4 ;
        RECT 169.515 3136.730 174.165 3275.270 ;
      LAYER met4 ;
        RECT 174.565 3274.965 175.165 3275.670 ;
        RECT 180.615 3275.365 186.065 3275.670 ;
        RECT 174.565 3136.330 175.165 3136.970 ;
      LAYER met4 ;
        RECT 175.565 3136.730 180.215 3275.270 ;
      LAYER met4 ;
        RECT 180.615 3274.965 181.215 3275.365 ;
        RECT 185.465 3274.965 186.065 3275.365 ;
      LAYER met4 ;
        RECT 181.615 3136.970 185.065 3274.965 ;
      LAYER met4 ;
        RECT 180.615 3136.570 181.215 3136.970 ;
        RECT 185.465 3136.570 186.065 3136.970 ;
      LAYER met4 ;
        RECT 186.465 3136.730 191.115 3275.270 ;
      LAYER met4 ;
        RECT 191.515 3274.965 192.115 3275.670 ;
        RECT 180.615 3136.330 186.065 3136.570 ;
        RECT 191.515 3136.330 192.115 3136.970 ;
      LAYER met4 ;
        RECT 192.515 3136.730 197.965 3275.270 ;
      LAYER met4 ;
        RECT 198.365 3274.965 199.465 3275.670 ;
        RECT 3388.535 3268.330 3389.635 3269.035 ;
      LAYER met4 ;
        RECT 3390.035 3268.730 3395.485 3417.270 ;
      LAYER met4 ;
        RECT 3395.885 3417.030 3396.485 3417.670 ;
        RECT 3401.935 3417.430 3407.385 3417.670 ;
        RECT 3395.885 3268.330 3396.485 3269.035 ;
      LAYER met4 ;
        RECT 3396.885 3268.730 3401.535 3417.270 ;
      LAYER met4 ;
        RECT 3401.935 3417.030 3402.535 3417.430 ;
        RECT 3406.785 3417.030 3407.385 3417.430 ;
      LAYER met4 ;
        RECT 3402.935 3269.035 3406.385 3417.030 ;
      LAYER met4 ;
        RECT 3401.935 3268.635 3402.535 3269.035 ;
        RECT 3406.785 3268.635 3407.385 3269.035 ;
      LAYER met4 ;
        RECT 3407.785 3268.730 3412.435 3417.270 ;
      LAYER met4 ;
        RECT 3412.835 3417.030 3413.435 3417.670 ;
        RECT 3401.935 3268.330 3407.385 3268.635 ;
        RECT 3412.835 3268.330 3413.435 3269.035 ;
      LAYER met4 ;
        RECT 3413.835 3268.730 3418.485 3417.270 ;
      LAYER met4 ;
        RECT 3418.885 3417.030 3419.485 3417.670 ;
        RECT 3418.885 3268.330 3419.485 3269.035 ;
      LAYER met4 ;
        RECT 3419.885 3268.730 3423.335 3417.270 ;
      LAYER met4 ;
        RECT 3423.735 3417.030 3424.335 3417.670 ;
        RECT 3423.735 3268.330 3424.335 3269.035 ;
      LAYER met4 ;
        RECT 3424.735 3268.730 3428.185 3417.270 ;
      LAYER met4 ;
        RECT 3428.585 3417.030 3429.185 3417.670 ;
        RECT 3428.585 3268.330 3429.185 3269.035 ;
      LAYER met4 ;
        RECT 3429.585 3268.730 3434.235 3417.270 ;
      LAYER met4 ;
        RECT 3434.635 3417.030 3435.335 3417.670 ;
        RECT 3434.635 3268.330 3435.335 3269.035 ;
        RECT 3388.535 3266.990 3435.335 3268.330 ;
      LAYER met4 ;
        RECT 3435.735 3267.390 3436.065 3448.910 ;
        RECT 3436.365 3443.855 3439.345 3666.535 ;
      LAYER met4 ;
        RECT 3439.745 3642.670 3440.725 3666.935 ;
      LAYER met4 ;
        RECT 3439.645 3641.000 3440.825 3642.270 ;
      LAYER met4 ;
        RECT 3439.645 3496.000 3440.825 3641.000 ;
      LAYER met4 ;
        RECT 3439.645 3494.730 3440.825 3496.000 ;
      LAYER met4 ;
        RECT 3439.745 3459.160 3440.725 3494.330 ;
      LAYER met4 ;
        RECT 3441.125 3459.560 3444.105 3682.240 ;
      LAYER met4 ;
        RECT 3444.505 3674.310 3588.000 3682.640 ;
      LAYER met4 ;
        RECT 3444.405 3493.390 3444.735 3673.910 ;
      LAYER met4 ;
        RECT 3445.135 3642.670 3588.000 3674.310 ;
        RECT 3445.135 3642.030 3445.835 3642.670 ;
        RECT 3445.135 3496.000 3445.835 3641.000 ;
        RECT 3445.135 3494.330 3445.835 3495.035 ;
      LAYER met4 ;
        RECT 3446.235 3494.730 3450.685 3642.270 ;
      LAYER met4 ;
        RECT 3451.085 3642.030 3451.685 3642.670 ;
        RECT 3451.085 3496.000 3451.685 3641.000 ;
        RECT 3451.085 3494.330 3451.685 3495.035 ;
      LAYER met4 ;
        RECT 3452.085 3494.730 3456.535 3642.270 ;
      LAYER met4 ;
        RECT 3456.935 3642.030 3457.635 3642.670 ;
        RECT 3456.935 3496.000 3457.635 3641.000 ;
        RECT 3456.935 3494.330 3457.635 3495.035 ;
      LAYER met4 ;
        RECT 3458.035 3494.730 3483.000 3642.270 ;
      LAYER met4 ;
        RECT 3483.400 3642.030 3563.385 3642.670 ;
      LAYER met4 ;
        RECT 3563.785 3641.000 3588.000 3642.270 ;
      LAYER met4 ;
        RECT 3483.400 3496.000 3588.000 3641.000 ;
        RECT 3483.400 3494.330 3563.385 3495.035 ;
      LAYER met4 ;
        RECT 3563.785 3494.730 3588.000 3496.000 ;
      LAYER met4 ;
        RECT 3445.135 3492.990 3588.000 3494.330 ;
        RECT 3444.505 3459.160 3588.000 3492.990 ;
        RECT 3439.745 3457.640 3588.000 3459.160 ;
        RECT 3439.745 3443.455 3440.725 3457.640 ;
        RECT 3436.465 3441.935 3440.725 3443.455 ;
        RECT 3388.535 3223.310 3435.965 3266.990 ;
        RECT 3388.535 3191.670 3435.335 3223.310 ;
        RECT 3388.535 3191.030 3389.635 3191.670 ;
        RECT 198.365 3136.330 199.465 3136.970 ;
        RECT 152.665 3104.690 199.465 3136.330 ;
        RECT 152.035 3061.010 199.465 3104.690 ;
        RECT 147.275 2894.545 151.535 2896.065 ;
        RECT 147.275 2880.360 148.255 2894.545 ;
        RECT 0.000 2878.840 148.255 2880.360 ;
        RECT 0.000 2845.010 143.495 2878.840 ;
        RECT 0.000 2843.670 142.865 2845.010 ;
      LAYER met4 ;
        RECT 0.000 2842.000 24.215 2843.270 ;
      LAYER met4 ;
        RECT 24.615 2842.965 104.600 2843.670 ;
        RECT 0.000 2706.000 104.600 2842.000 ;
      LAYER met4 ;
        RECT 0.000 2704.730 24.215 2706.000 ;
      LAYER met4 ;
        RECT 24.615 2704.330 104.600 2704.970 ;
      LAYER met4 ;
        RECT 105.000 2704.730 129.965 2843.270 ;
      LAYER met4 ;
        RECT 130.365 2842.965 131.065 2843.670 ;
        RECT 130.365 2706.000 131.065 2842.000 ;
        RECT 130.365 2704.330 131.065 2704.970 ;
      LAYER met4 ;
        RECT 131.465 2704.730 135.915 2843.270 ;
      LAYER met4 ;
        RECT 136.315 2842.965 136.915 2843.670 ;
        RECT 136.315 2706.000 136.915 2842.000 ;
        RECT 136.315 2704.330 136.915 2704.970 ;
      LAYER met4 ;
        RECT 137.315 2704.730 141.765 2843.270 ;
      LAYER met4 ;
        RECT 142.165 2842.965 142.865 2843.670 ;
        RECT 142.165 2706.000 142.865 2842.000 ;
        RECT 142.165 2704.330 142.865 2704.970 ;
        RECT 0.000 2672.690 142.865 2704.330 ;
      LAYER met4 ;
        RECT 143.265 2673.090 143.595 2844.610 ;
      LAYER met4 ;
        RECT 0.000 2664.360 143.495 2672.690 ;
      LAYER met4 ;
        RECT 143.895 2664.760 146.875 2878.440 ;
      LAYER met4 ;
        RECT 147.275 2843.670 148.255 2878.840 ;
      LAYER met4 ;
        RECT 147.175 2842.000 148.355 2843.270 ;
      LAYER met4 ;
        RECT 147.175 2706.000 148.355 2842.000 ;
      LAYER met4 ;
        RECT 147.175 2704.730 148.355 2706.000 ;
      LAYER met4 ;
        RECT 147.275 2680.065 148.255 2704.330 ;
      LAYER met4 ;
        RECT 148.655 2680.465 151.635 2894.145 ;
        RECT 151.935 2889.090 152.265 3060.610 ;
      LAYER met4 ;
        RECT 152.665 3059.670 199.465 3061.010 ;
        RECT 152.665 3058.965 153.365 3059.670 ;
        RECT 152.665 2920.330 153.365 2920.970 ;
      LAYER met4 ;
        RECT 153.765 2920.730 158.415 3059.270 ;
      LAYER met4 ;
        RECT 158.815 3058.965 159.415 3059.670 ;
        RECT 158.815 2920.330 159.415 2920.970 ;
      LAYER met4 ;
        RECT 159.815 2920.730 163.265 3059.270 ;
      LAYER met4 ;
        RECT 163.665 3058.965 164.265 3059.670 ;
        RECT 163.665 2920.330 164.265 2920.970 ;
      LAYER met4 ;
        RECT 164.665 2920.730 168.115 3059.270 ;
      LAYER met4 ;
        RECT 168.515 3058.965 169.115 3059.670 ;
        RECT 168.515 2920.330 169.115 2920.970 ;
      LAYER met4 ;
        RECT 169.515 2920.730 174.165 3059.270 ;
      LAYER met4 ;
        RECT 174.565 3058.965 175.165 3059.670 ;
        RECT 180.615 3059.365 186.065 3059.670 ;
        RECT 174.565 2920.330 175.165 2920.970 ;
      LAYER met4 ;
        RECT 175.565 2920.730 180.215 3059.270 ;
      LAYER met4 ;
        RECT 180.615 3058.965 181.215 3059.365 ;
        RECT 185.465 3058.965 186.065 3059.365 ;
      LAYER met4 ;
        RECT 181.615 2920.970 185.065 3058.965 ;
      LAYER met4 ;
        RECT 180.615 2920.570 181.215 2920.970 ;
        RECT 185.465 2920.570 186.065 2920.970 ;
      LAYER met4 ;
        RECT 186.465 2920.730 191.115 3059.270 ;
      LAYER met4 ;
        RECT 191.515 3058.965 192.115 3059.670 ;
        RECT 180.615 2920.330 186.065 2920.570 ;
        RECT 191.515 2920.330 192.115 2920.970 ;
      LAYER met4 ;
        RECT 192.515 2920.730 197.965 3059.270 ;
      LAYER met4 ;
        RECT 198.365 3058.965 199.465 3059.670 ;
        RECT 3388.535 3043.330 3389.635 3044.035 ;
      LAYER met4 ;
        RECT 3390.035 3043.730 3395.485 3191.270 ;
      LAYER met4 ;
        RECT 3395.885 3191.030 3396.485 3191.670 ;
        RECT 3401.935 3191.430 3407.385 3191.670 ;
        RECT 3395.885 3043.330 3396.485 3044.035 ;
      LAYER met4 ;
        RECT 3396.885 3043.730 3401.535 3191.270 ;
      LAYER met4 ;
        RECT 3401.935 3191.030 3402.535 3191.430 ;
        RECT 3406.785 3191.030 3407.385 3191.430 ;
      LAYER met4 ;
        RECT 3402.935 3044.035 3406.385 3191.030 ;
      LAYER met4 ;
        RECT 3401.935 3043.635 3402.535 3044.035 ;
        RECT 3406.785 3043.635 3407.385 3044.035 ;
      LAYER met4 ;
        RECT 3407.785 3043.730 3412.435 3191.270 ;
      LAYER met4 ;
        RECT 3412.835 3191.030 3413.435 3191.670 ;
        RECT 3401.935 3043.330 3407.385 3043.635 ;
        RECT 3412.835 3043.330 3413.435 3044.035 ;
      LAYER met4 ;
        RECT 3413.835 3043.730 3418.485 3191.270 ;
      LAYER met4 ;
        RECT 3418.885 3191.030 3419.485 3191.670 ;
        RECT 3418.885 3043.330 3419.485 3044.035 ;
      LAYER met4 ;
        RECT 3419.885 3043.730 3423.335 3191.270 ;
      LAYER met4 ;
        RECT 3423.735 3191.030 3424.335 3191.670 ;
        RECT 3423.735 3043.330 3424.335 3044.035 ;
      LAYER met4 ;
        RECT 3424.735 3043.730 3428.185 3191.270 ;
      LAYER met4 ;
        RECT 3428.585 3191.030 3429.185 3191.670 ;
        RECT 3428.585 3043.330 3429.185 3044.035 ;
      LAYER met4 ;
        RECT 3429.585 3043.730 3434.235 3191.270 ;
      LAYER met4 ;
        RECT 3434.635 3191.030 3435.335 3191.670 ;
        RECT 3434.635 3043.330 3435.335 3044.035 ;
        RECT 3388.535 3041.990 3435.335 3043.330 ;
      LAYER met4 ;
        RECT 3435.735 3042.390 3436.065 3222.910 ;
        RECT 3436.365 3217.855 3439.345 3441.535 ;
      LAYER met4 ;
        RECT 3439.745 3417.670 3440.725 3441.935 ;
      LAYER met4 ;
        RECT 3439.645 3416.000 3440.825 3417.270 ;
      LAYER met4 ;
        RECT 3439.645 3270.000 3440.825 3416.000 ;
      LAYER met4 ;
        RECT 3439.645 3268.730 3440.825 3270.000 ;
      LAYER met4 ;
        RECT 3439.745 3233.160 3440.725 3268.330 ;
      LAYER met4 ;
        RECT 3441.125 3233.560 3444.105 3457.240 ;
      LAYER met4 ;
        RECT 3444.505 3449.310 3588.000 3457.640 ;
      LAYER met4 ;
        RECT 3444.405 3267.390 3444.735 3448.910 ;
      LAYER met4 ;
        RECT 3445.135 3417.670 3588.000 3449.310 ;
        RECT 3445.135 3417.030 3445.835 3417.670 ;
        RECT 3445.135 3270.000 3445.835 3416.000 ;
        RECT 3445.135 3268.330 3445.835 3269.035 ;
      LAYER met4 ;
        RECT 3446.235 3268.730 3450.685 3417.270 ;
      LAYER met4 ;
        RECT 3451.085 3417.030 3451.685 3417.670 ;
        RECT 3451.085 3270.000 3451.685 3416.000 ;
        RECT 3451.085 3268.330 3451.685 3269.035 ;
      LAYER met4 ;
        RECT 3452.085 3268.730 3456.535 3417.270 ;
      LAYER met4 ;
        RECT 3456.935 3417.030 3457.635 3417.670 ;
        RECT 3456.935 3270.000 3457.635 3416.000 ;
        RECT 3456.935 3268.330 3457.635 3269.035 ;
      LAYER met4 ;
        RECT 3458.035 3268.730 3483.000 3417.270 ;
      LAYER met4 ;
        RECT 3483.400 3417.030 3563.385 3417.670 ;
      LAYER met4 ;
        RECT 3563.785 3416.000 3588.000 3417.270 ;
      LAYER met4 ;
        RECT 3483.400 3270.000 3588.000 3416.000 ;
        RECT 3483.400 3268.330 3563.385 3269.035 ;
      LAYER met4 ;
        RECT 3563.785 3268.730 3588.000 3270.000 ;
      LAYER met4 ;
        RECT 3445.135 3266.990 3588.000 3268.330 ;
        RECT 3444.505 3233.160 3588.000 3266.990 ;
        RECT 3439.745 3231.640 3588.000 3233.160 ;
        RECT 3439.745 3217.455 3440.725 3231.640 ;
        RECT 3436.465 3215.935 3440.725 3217.455 ;
        RECT 3388.535 2998.310 3435.965 3041.990 ;
        RECT 3388.535 2966.670 3435.335 2998.310 ;
        RECT 3388.535 2966.030 3389.635 2966.670 ;
        RECT 198.365 2920.330 199.465 2920.970 ;
        RECT 152.665 2888.690 199.465 2920.330 ;
        RECT 152.035 2845.010 199.465 2888.690 ;
        RECT 147.275 2678.545 151.535 2680.065 ;
        RECT 147.275 2664.360 148.255 2678.545 ;
        RECT 0.000 2662.840 148.255 2664.360 ;
        RECT 0.000 2629.010 143.495 2662.840 ;
        RECT 0.000 2627.670 142.865 2629.010 ;
      LAYER met4 ;
        RECT 0.000 2626.000 24.215 2627.270 ;
      LAYER met4 ;
        RECT 24.615 2626.965 104.600 2627.670 ;
        RECT 0.000 2490.000 104.600 2626.000 ;
      LAYER met4 ;
        RECT 0.000 2488.730 24.215 2490.000 ;
      LAYER met4 ;
        RECT 24.615 2488.330 104.600 2489.035 ;
      LAYER met4 ;
        RECT 105.000 2488.730 129.965 2627.270 ;
      LAYER met4 ;
        RECT 130.365 2626.965 131.065 2627.670 ;
        RECT 130.365 2490.000 131.065 2626.000 ;
        RECT 130.365 2488.330 131.065 2489.035 ;
      LAYER met4 ;
        RECT 131.465 2488.730 135.915 2627.270 ;
      LAYER met4 ;
        RECT 136.315 2626.965 136.915 2627.670 ;
        RECT 136.315 2490.000 136.915 2626.000 ;
        RECT 136.315 2488.330 136.915 2489.035 ;
      LAYER met4 ;
        RECT 137.315 2488.730 141.765 2627.270 ;
      LAYER met4 ;
        RECT 142.165 2626.965 142.865 2627.670 ;
        RECT 142.165 2490.000 142.865 2626.000 ;
        RECT 142.165 2488.330 142.865 2489.035 ;
        RECT 0.000 2416.670 142.865 2488.330 ;
      LAYER met4 ;
        RECT 0.000 2415.000 24.215 2416.270 ;
      LAYER met4 ;
        RECT 24.615 2415.965 104.600 2416.670 ;
        RECT 0.000 2280.465 104.600 2415.000 ;
        RECT 0.000 2279.000 0.035 2280.465 ;
        RECT 24.215 2279.000 104.600 2280.465 ;
      LAYER met4 ;
        RECT 105.000 2279.000 129.965 2416.270 ;
      LAYER met4 ;
        RECT 130.365 2415.965 131.065 2416.670 ;
        RECT 130.365 2279.000 131.065 2415.000 ;
      LAYER met4 ;
        RECT 131.465 2279.000 135.915 2416.270 ;
      LAYER met4 ;
        RECT 136.315 2415.965 136.915 2416.670 ;
        RECT 136.315 2279.000 136.915 2415.000 ;
      LAYER met4 ;
        RECT 137.315 2279.000 141.765 2416.270 ;
      LAYER met4 ;
        RECT 142.165 2415.965 142.865 2416.670 ;
        RECT 142.165 2279.000 142.865 2415.000 ;
      LAYER met4 ;
        RECT 143.895 2279.000 146.875 2662.440 ;
      LAYER met4 ;
        RECT 147.275 2627.670 148.255 2662.840 ;
      LAYER met4 ;
        RECT 147.175 2626.000 148.355 2627.270 ;
      LAYER met4 ;
        RECT 147.175 2490.000 148.355 2626.000 ;
      LAYER met4 ;
        RECT 147.175 2488.730 148.355 2490.000 ;
      LAYER met4 ;
        RECT 147.275 2416.670 148.255 2488.330 ;
      LAYER met4 ;
        RECT 147.175 2415.000 148.355 2416.270 ;
      LAYER met4 ;
        RECT 147.175 2279.000 148.355 2415.000 ;
      LAYER met4 ;
        RECT 148.655 2279.000 151.635 2678.145 ;
        RECT 151.935 2673.090 152.265 2844.610 ;
      LAYER met4 ;
        RECT 152.665 2843.670 199.465 2845.010 ;
        RECT 152.665 2842.965 153.365 2843.670 ;
        RECT 152.665 2704.330 153.365 2704.970 ;
      LAYER met4 ;
        RECT 153.765 2704.730 158.415 2843.270 ;
      LAYER met4 ;
        RECT 158.815 2842.965 159.415 2843.670 ;
        RECT 158.815 2704.330 159.415 2704.970 ;
      LAYER met4 ;
        RECT 159.815 2704.730 163.265 2843.270 ;
      LAYER met4 ;
        RECT 163.665 2842.965 164.265 2843.670 ;
        RECT 163.665 2704.330 164.265 2704.970 ;
      LAYER met4 ;
        RECT 164.665 2704.730 168.115 2843.270 ;
      LAYER met4 ;
        RECT 168.515 2842.965 169.115 2843.670 ;
        RECT 168.515 2704.330 169.115 2704.970 ;
      LAYER met4 ;
        RECT 169.515 2704.730 174.165 2843.270 ;
      LAYER met4 ;
        RECT 174.565 2842.965 175.165 2843.670 ;
        RECT 180.615 2843.365 186.065 2843.670 ;
        RECT 174.565 2704.330 175.165 2704.970 ;
      LAYER met4 ;
        RECT 175.565 2704.730 180.215 2843.270 ;
      LAYER met4 ;
        RECT 180.615 2842.965 181.215 2843.365 ;
        RECT 185.465 2842.965 186.065 2843.365 ;
      LAYER met4 ;
        RECT 181.615 2704.970 185.065 2842.965 ;
      LAYER met4 ;
        RECT 180.615 2704.570 181.215 2704.970 ;
        RECT 185.465 2704.570 186.065 2704.970 ;
      LAYER met4 ;
        RECT 186.465 2704.730 191.115 2843.270 ;
      LAYER met4 ;
        RECT 191.515 2842.965 192.115 2843.670 ;
        RECT 180.615 2704.330 186.065 2704.570 ;
        RECT 191.515 2704.330 192.115 2704.970 ;
      LAYER met4 ;
        RECT 192.515 2704.730 197.965 2843.270 ;
      LAYER met4 ;
        RECT 198.365 2842.965 199.465 2843.670 ;
        RECT 3388.535 2817.330 3389.635 2818.035 ;
      LAYER met4 ;
        RECT 3390.035 2817.730 3395.485 2966.270 ;
      LAYER met4 ;
        RECT 3395.885 2966.030 3396.485 2966.670 ;
        RECT 3401.935 2966.430 3407.385 2966.670 ;
        RECT 3395.885 2817.330 3396.485 2818.035 ;
      LAYER met4 ;
        RECT 3396.885 2817.730 3401.535 2966.270 ;
      LAYER met4 ;
        RECT 3401.935 2966.030 3402.535 2966.430 ;
        RECT 3406.785 2966.030 3407.385 2966.430 ;
      LAYER met4 ;
        RECT 3402.935 2818.035 3406.385 2966.030 ;
      LAYER met4 ;
        RECT 3401.935 2817.635 3402.535 2818.035 ;
        RECT 3406.785 2817.635 3407.385 2818.035 ;
      LAYER met4 ;
        RECT 3407.785 2817.730 3412.435 2966.270 ;
      LAYER met4 ;
        RECT 3412.835 2966.030 3413.435 2966.670 ;
        RECT 3401.935 2817.330 3407.385 2817.635 ;
        RECT 3412.835 2817.330 3413.435 2818.035 ;
      LAYER met4 ;
        RECT 3413.835 2817.730 3418.485 2966.270 ;
      LAYER met4 ;
        RECT 3418.885 2966.030 3419.485 2966.670 ;
        RECT 3418.885 2817.330 3419.485 2818.035 ;
      LAYER met4 ;
        RECT 3419.885 2817.730 3423.335 2966.270 ;
      LAYER met4 ;
        RECT 3423.735 2966.030 3424.335 2966.670 ;
        RECT 3423.735 2817.330 3424.335 2818.035 ;
      LAYER met4 ;
        RECT 3424.735 2817.730 3428.185 2966.270 ;
      LAYER met4 ;
        RECT 3428.585 2966.030 3429.185 2966.670 ;
        RECT 3428.585 2817.330 3429.185 2818.035 ;
      LAYER met4 ;
        RECT 3429.585 2817.730 3434.235 2966.270 ;
      LAYER met4 ;
        RECT 3434.635 2966.030 3435.335 2966.670 ;
        RECT 3434.635 2817.330 3435.335 2818.035 ;
        RECT 3388.535 2815.990 3435.335 2817.330 ;
      LAYER met4 ;
        RECT 3435.735 2816.390 3436.065 2997.910 ;
        RECT 3436.365 2992.855 3439.345 3215.535 ;
      LAYER met4 ;
        RECT 3439.745 3191.670 3440.725 3215.935 ;
      LAYER met4 ;
        RECT 3439.645 3190.000 3440.825 3191.270 ;
      LAYER met4 ;
        RECT 3439.645 3045.000 3440.825 3190.000 ;
      LAYER met4 ;
        RECT 3439.645 3043.730 3440.825 3045.000 ;
      LAYER met4 ;
        RECT 3439.745 3008.160 3440.725 3043.330 ;
      LAYER met4 ;
        RECT 3441.125 3008.560 3444.105 3231.240 ;
      LAYER met4 ;
        RECT 3444.505 3223.310 3588.000 3231.640 ;
      LAYER met4 ;
        RECT 3444.405 3042.390 3444.735 3222.910 ;
      LAYER met4 ;
        RECT 3445.135 3191.670 3588.000 3223.310 ;
        RECT 3445.135 3191.030 3445.835 3191.670 ;
        RECT 3445.135 3045.000 3445.835 3190.000 ;
        RECT 3445.135 3043.330 3445.835 3044.035 ;
      LAYER met4 ;
        RECT 3446.235 3043.730 3450.685 3191.270 ;
      LAYER met4 ;
        RECT 3451.085 3191.030 3451.685 3191.670 ;
        RECT 3451.085 3045.000 3451.685 3190.000 ;
        RECT 3451.085 3043.330 3451.685 3044.035 ;
      LAYER met4 ;
        RECT 3452.085 3043.730 3456.535 3191.270 ;
      LAYER met4 ;
        RECT 3456.935 3191.030 3457.635 3191.670 ;
        RECT 3456.935 3045.000 3457.635 3190.000 ;
        RECT 3456.935 3043.330 3457.635 3044.035 ;
      LAYER met4 ;
        RECT 3458.035 3043.730 3483.000 3191.270 ;
      LAYER met4 ;
        RECT 3483.400 3191.030 3563.385 3191.670 ;
      LAYER met4 ;
        RECT 3563.785 3190.000 3588.000 3191.270 ;
      LAYER met4 ;
        RECT 3483.400 3045.000 3588.000 3190.000 ;
        RECT 3483.400 3043.330 3563.385 3044.035 ;
      LAYER met4 ;
        RECT 3563.785 3043.730 3588.000 3045.000 ;
      LAYER met4 ;
        RECT 3445.135 3041.990 3588.000 3043.330 ;
        RECT 3444.505 3008.160 3588.000 3041.990 ;
        RECT 3439.745 3006.640 3588.000 3008.160 ;
        RECT 3439.745 2992.455 3440.725 3006.640 ;
        RECT 3436.465 2990.935 3440.725 2992.455 ;
        RECT 3388.535 2772.310 3435.965 2815.990 ;
        RECT 3388.535 2740.670 3435.335 2772.310 ;
        RECT 3388.535 2740.030 3389.635 2740.670 ;
        RECT 198.365 2704.330 199.465 2704.970 ;
        RECT 152.665 2672.690 199.465 2704.330 ;
        RECT 152.035 2629.010 199.465 2672.690 ;
      LAYER met4 ;
        RECT 151.935 2279.000 152.265 2628.610 ;
      LAYER met4 ;
        RECT 152.665 2627.670 199.465 2629.010 ;
        RECT 152.665 2626.965 153.365 2627.670 ;
        RECT 152.665 2488.330 153.365 2489.035 ;
      LAYER met4 ;
        RECT 153.765 2488.730 158.415 2627.270 ;
      LAYER met4 ;
        RECT 158.815 2626.965 159.415 2627.670 ;
        RECT 158.815 2488.330 159.415 2489.035 ;
      LAYER met4 ;
        RECT 159.815 2488.730 163.265 2627.270 ;
      LAYER met4 ;
        RECT 163.665 2626.965 164.265 2627.670 ;
        RECT 163.665 2488.330 164.265 2489.035 ;
      LAYER met4 ;
        RECT 164.665 2488.730 168.115 2627.270 ;
      LAYER met4 ;
        RECT 168.515 2626.965 169.115 2627.670 ;
        RECT 168.515 2488.330 169.115 2489.035 ;
      LAYER met4 ;
        RECT 169.515 2488.730 174.165 2627.270 ;
      LAYER met4 ;
        RECT 174.565 2626.965 175.165 2627.670 ;
        RECT 180.615 2627.365 186.065 2627.670 ;
        RECT 174.565 2488.330 175.165 2489.035 ;
      LAYER met4 ;
        RECT 175.565 2488.730 180.215 2627.270 ;
      LAYER met4 ;
        RECT 180.615 2626.965 181.215 2627.365 ;
        RECT 185.465 2626.965 186.065 2627.365 ;
      LAYER met4 ;
        RECT 181.615 2489.035 185.065 2626.965 ;
      LAYER met4 ;
        RECT 180.615 2488.635 181.215 2489.035 ;
        RECT 185.465 2488.635 186.065 2489.035 ;
      LAYER met4 ;
        RECT 186.465 2488.730 191.115 2627.270 ;
      LAYER met4 ;
        RECT 191.515 2626.965 192.115 2627.670 ;
        RECT 180.615 2488.330 186.065 2488.635 ;
        RECT 191.515 2488.330 192.115 2489.035 ;
      LAYER met4 ;
        RECT 192.515 2488.730 197.965 2627.270 ;
      LAYER met4 ;
        RECT 198.365 2626.965 199.465 2627.670 ;
      LAYER met4 ;
        RECT 3390.035 2592.730 3395.485 2740.270 ;
      LAYER met4 ;
        RECT 3395.885 2740.030 3396.485 2740.670 ;
        RECT 3401.935 2740.430 3407.385 2740.670 ;
        RECT 3395.885 2592.330 3396.485 2593.035 ;
      LAYER met4 ;
        RECT 3396.885 2592.730 3401.535 2740.270 ;
      LAYER met4 ;
        RECT 3401.935 2740.030 3402.535 2740.430 ;
        RECT 3406.785 2740.030 3407.385 2740.430 ;
      LAYER met4 ;
        RECT 3402.935 2593.035 3406.385 2740.030 ;
      LAYER met4 ;
        RECT 3401.935 2592.635 3402.535 2593.035 ;
        RECT 3406.785 2592.635 3407.385 2593.035 ;
      LAYER met4 ;
        RECT 3407.785 2592.730 3412.435 2740.270 ;
      LAYER met4 ;
        RECT 3412.835 2740.030 3413.435 2740.670 ;
        RECT 3401.935 2592.330 3407.385 2592.635 ;
        RECT 3412.835 2592.330 3413.435 2593.035 ;
      LAYER met4 ;
        RECT 3413.835 2592.730 3418.485 2740.270 ;
      LAYER met4 ;
        RECT 3418.885 2740.030 3419.485 2740.670 ;
        RECT 3418.885 2592.330 3419.485 2593.035 ;
      LAYER met4 ;
        RECT 3419.885 2592.730 3423.335 2740.270 ;
      LAYER met4 ;
        RECT 3423.735 2740.030 3424.335 2740.670 ;
        RECT 3423.735 2592.330 3424.335 2593.035 ;
      LAYER met4 ;
        RECT 3424.735 2592.730 3428.185 2740.270 ;
      LAYER met4 ;
        RECT 3428.585 2740.030 3429.185 2740.670 ;
        RECT 3428.585 2592.330 3429.185 2593.035 ;
      LAYER met4 ;
        RECT 3429.585 2592.730 3434.235 2740.270 ;
      LAYER met4 ;
        RECT 3434.635 2740.030 3435.335 2740.670 ;
        RECT 3434.635 2592.330 3435.335 2593.035 ;
        RECT 3390.035 2520.670 3435.335 2592.330 ;
        RECT 152.665 2416.670 197.965 2488.330 ;
        RECT 152.665 2415.965 153.365 2416.670 ;
      LAYER met4 ;
        RECT 153.765 2279.000 158.415 2416.270 ;
      LAYER met4 ;
        RECT 158.815 2415.965 159.415 2416.670 ;
      LAYER met4 ;
        RECT 159.815 2279.000 163.265 2416.270 ;
      LAYER met4 ;
        RECT 163.665 2415.965 164.265 2416.670 ;
        RECT 168.515 2415.965 169.115 2416.670 ;
      LAYER met4 ;
        RECT 169.515 2279.000 174.165 2416.270 ;
      LAYER met4 ;
        RECT 174.565 2415.965 175.165 2416.670 ;
        RECT 180.615 2416.365 186.065 2416.670 ;
      LAYER met4 ;
        RECT 175.565 2279.000 180.215 2416.270 ;
      LAYER met4 ;
        RECT 180.615 2415.965 181.215 2416.365 ;
        RECT 185.465 2415.965 186.065 2416.365 ;
      LAYER met4 ;
        RECT 181.615 2279.000 185.065 2415.965 ;
        RECT 186.465 2277.730 191.115 2416.270 ;
      LAYER met4 ;
        RECT 191.515 2415.965 192.115 2416.670 ;
      LAYER met4 ;
        RECT 3390.035 2374.000 3395.485 2520.270 ;
      LAYER met4 ;
        RECT 3395.885 2519.965 3396.485 2520.670 ;
        RECT 3401.935 2520.365 3407.385 2520.670 ;
      LAYER met4 ;
        RECT 3396.885 2374.000 3401.535 2520.270 ;
      LAYER met4 ;
        RECT 3401.935 2519.965 3402.535 2520.365 ;
        RECT 3406.785 2519.965 3407.385 2520.365 ;
      LAYER met4 ;
        RECT 3402.935 2374.000 3406.385 2519.965 ;
        RECT 3407.785 2374.000 3412.435 2520.270 ;
      LAYER met4 ;
        RECT 3412.835 2519.965 3413.435 2520.670 ;
      LAYER met4 ;
        RECT 3413.835 2374.000 3418.485 2520.270 ;
      LAYER met4 ;
        RECT 3418.885 2519.965 3419.485 2520.670 ;
      LAYER met4 ;
        RECT 3419.885 2374.000 3423.335 2520.270 ;
      LAYER met4 ;
        RECT 3423.735 2519.965 3424.335 2520.670 ;
      LAYER met4 ;
        RECT 3424.735 2374.000 3428.185 2520.270 ;
      LAYER met4 ;
        RECT 3428.585 2519.965 3429.185 2520.670 ;
      LAYER met4 ;
        RECT 3429.585 2374.000 3434.235 2520.270 ;
      LAYER met4 ;
        RECT 3434.635 2519.965 3435.335 2520.670 ;
      LAYER met4 ;
        RECT 3435.735 2374.000 3436.065 2771.910 ;
        RECT 3436.365 2766.855 3439.345 2990.535 ;
      LAYER met4 ;
        RECT 3439.745 2966.670 3440.725 2990.935 ;
      LAYER met4 ;
        RECT 3439.645 2965.000 3440.825 2966.270 ;
      LAYER met4 ;
        RECT 3439.645 2819.000 3440.825 2965.000 ;
      LAYER met4 ;
        RECT 3439.645 2817.730 3440.825 2819.000 ;
      LAYER met4 ;
        RECT 3439.745 2782.160 3440.725 2817.330 ;
      LAYER met4 ;
        RECT 3441.125 2782.560 3444.105 3006.240 ;
      LAYER met4 ;
        RECT 3444.505 2998.310 3588.000 3006.640 ;
      LAYER met4 ;
        RECT 3444.405 2816.390 3444.735 2997.910 ;
      LAYER met4 ;
        RECT 3445.135 2966.670 3588.000 2998.310 ;
        RECT 3445.135 2966.030 3445.835 2966.670 ;
        RECT 3445.135 2819.000 3445.835 2965.000 ;
        RECT 3445.135 2817.330 3445.835 2818.035 ;
      LAYER met4 ;
        RECT 3446.235 2817.730 3450.685 2966.270 ;
      LAYER met4 ;
        RECT 3451.085 2966.030 3451.685 2966.670 ;
        RECT 3451.085 2819.000 3451.685 2965.000 ;
        RECT 3451.085 2817.330 3451.685 2818.035 ;
      LAYER met4 ;
        RECT 3452.085 2817.730 3456.535 2966.270 ;
      LAYER met4 ;
        RECT 3456.935 2966.030 3457.635 2966.670 ;
        RECT 3456.935 2819.000 3457.635 2965.000 ;
        RECT 3456.935 2817.330 3457.635 2818.035 ;
      LAYER met4 ;
        RECT 3458.035 2817.730 3483.000 2966.270 ;
      LAYER met4 ;
        RECT 3483.400 2966.030 3563.385 2966.670 ;
      LAYER met4 ;
        RECT 3563.785 2965.000 3588.000 2966.270 ;
      LAYER met4 ;
        RECT 3483.400 2819.000 3588.000 2965.000 ;
        RECT 3483.400 2817.330 3563.385 2818.035 ;
      LAYER met4 ;
        RECT 3563.785 2817.730 3588.000 2819.000 ;
      LAYER met4 ;
        RECT 3445.135 2815.990 3588.000 2817.330 ;
        RECT 3444.505 2782.160 3588.000 2815.990 ;
        RECT 3439.745 2780.640 3588.000 2782.160 ;
        RECT 3439.745 2766.455 3440.725 2780.640 ;
        RECT 3436.465 2764.935 3440.725 2766.455 ;
      LAYER met4 ;
        RECT 3436.365 2374.000 3439.345 2764.535 ;
      LAYER met4 ;
        RECT 3439.745 2740.670 3440.725 2764.935 ;
      LAYER met4 ;
        RECT 3439.645 2739.000 3440.825 2740.270 ;
      LAYER met4 ;
        RECT 3439.645 2594.000 3440.825 2739.000 ;
      LAYER met4 ;
        RECT 3439.645 2592.730 3440.825 2594.000 ;
      LAYER met4 ;
        RECT 3439.745 2520.670 3440.725 2592.330 ;
      LAYER met4 ;
        RECT 3439.645 2519.000 3440.825 2520.270 ;
      LAYER met4 ;
        RECT 3439.645 2374.000 3440.825 2519.000 ;
      LAYER met4 ;
        RECT 3441.125 2374.000 3444.105 2780.240 ;
      LAYER met4 ;
        RECT 3444.505 2772.310 3588.000 2780.640 ;
        RECT 3445.135 2740.670 3588.000 2772.310 ;
        RECT 3445.135 2740.030 3445.835 2740.670 ;
        RECT 3445.135 2594.000 3445.835 2739.000 ;
        RECT 3445.135 2592.330 3445.835 2593.035 ;
      LAYER met4 ;
        RECT 3446.235 2592.730 3450.685 2740.270 ;
      LAYER met4 ;
        RECT 3451.085 2740.030 3451.685 2740.670 ;
        RECT 3451.085 2594.000 3451.685 2739.000 ;
        RECT 3451.085 2592.330 3451.685 2593.035 ;
      LAYER met4 ;
        RECT 3452.085 2592.730 3456.535 2740.270 ;
      LAYER met4 ;
        RECT 3456.935 2740.030 3457.635 2740.670 ;
        RECT 3456.935 2594.000 3457.635 2739.000 ;
        RECT 3456.935 2592.330 3457.635 2593.035 ;
      LAYER met4 ;
        RECT 3458.035 2592.730 3483.000 2740.270 ;
      LAYER met4 ;
        RECT 3483.400 2740.030 3563.385 2740.670 ;
      LAYER met4 ;
        RECT 3563.785 2739.000 3588.000 2740.270 ;
      LAYER met4 ;
        RECT 3483.400 2594.000 3588.000 2739.000 ;
        RECT 3483.400 2592.330 3563.385 2593.035 ;
      LAYER met4 ;
        RECT 3563.785 2592.730 3588.000 2594.000 ;
      LAYER met4 ;
        RECT 3445.135 2520.670 3588.000 2592.330 ;
        RECT 3445.135 2519.965 3445.835 2520.670 ;
        RECT 3445.135 2374.000 3445.835 2519.000 ;
      LAYER met4 ;
        RECT 3446.235 2374.000 3450.685 2520.270 ;
      LAYER met4 ;
        RECT 3451.085 2519.965 3451.685 2520.670 ;
        RECT 3451.085 2374.000 3451.685 2519.000 ;
      LAYER met4 ;
        RECT 3452.085 2374.000 3456.535 2520.270 ;
      LAYER met4 ;
        RECT 3456.935 2519.965 3457.635 2520.670 ;
        RECT 3456.935 2374.000 3457.635 2519.000 ;
      LAYER met4 ;
        RECT 3458.035 2374.000 3483.000 2520.270 ;
      LAYER met4 ;
        RECT 3483.400 2519.965 3563.385 2520.670 ;
      LAYER met4 ;
        RECT 3563.785 2519.000 3588.000 2520.270 ;
      LAYER met4 ;
        RECT 3483.400 2374.000 3588.000 2519.000 ;
        RECT 0.000 2068.000 104.600 2204.000 ;
      LAYER met4 ;
        RECT 0.000 2066.730 24.215 2068.000 ;
      LAYER met4 ;
        RECT 24.615 2066.330 104.600 2066.970 ;
      LAYER met4 ;
        RECT 105.000 2066.730 129.965 2204.000 ;
      LAYER met4 ;
        RECT 130.365 2068.000 131.065 2204.000 ;
        RECT 130.365 2066.330 131.065 2066.970 ;
      LAYER met4 ;
        RECT 131.465 2066.730 135.915 2204.000 ;
      LAYER met4 ;
        RECT 136.315 2068.000 136.915 2204.000 ;
        RECT 136.315 2066.330 136.915 2066.970 ;
      LAYER met4 ;
        RECT 137.315 2066.730 141.765 2204.000 ;
      LAYER met4 ;
        RECT 142.165 2068.000 142.865 2204.000 ;
        RECT 142.165 2066.330 142.865 2066.970 ;
        RECT 0.000 2034.690 142.865 2066.330 ;
        RECT 0.000 2026.360 143.495 2034.690 ;
      LAYER met4 ;
        RECT 143.895 2026.760 146.875 2204.000 ;
      LAYER met4 ;
        RECT 147.175 2068.000 148.355 2204.000 ;
      LAYER met4 ;
        RECT 147.175 2066.730 148.355 2068.000 ;
      LAYER met4 ;
        RECT 147.275 2042.065 148.255 2066.330 ;
      LAYER met4 ;
        RECT 148.655 2042.465 151.635 2204.000 ;
      LAYER met4 ;
        RECT 147.275 2040.545 151.535 2042.065 ;
        RECT 147.275 2026.360 148.255 2040.545 ;
        RECT 0.000 2024.840 148.255 2026.360 ;
        RECT 0.000 1991.010 143.495 2024.840 ;
        RECT 0.000 1989.670 142.865 1991.010 ;
      LAYER met4 ;
        RECT 0.000 1988.000 24.215 1989.270 ;
      LAYER met4 ;
        RECT 24.615 1988.965 104.600 1989.670 ;
        RECT 0.000 1852.000 104.600 1988.000 ;
      LAYER met4 ;
        RECT 0.000 1850.730 24.215 1852.000 ;
      LAYER met4 ;
        RECT 24.615 1850.330 104.600 1850.970 ;
      LAYER met4 ;
        RECT 105.000 1850.730 129.965 1989.270 ;
      LAYER met4 ;
        RECT 130.365 1988.965 131.065 1989.670 ;
        RECT 130.365 1852.000 131.065 1988.000 ;
        RECT 130.365 1850.330 131.065 1850.970 ;
      LAYER met4 ;
        RECT 131.465 1850.730 135.915 1989.270 ;
      LAYER met4 ;
        RECT 136.315 1988.965 136.915 1989.670 ;
        RECT 136.315 1852.000 136.915 1988.000 ;
        RECT 136.315 1850.330 136.915 1850.970 ;
      LAYER met4 ;
        RECT 137.315 1850.730 141.765 1989.270 ;
      LAYER met4 ;
        RECT 142.165 1988.965 142.865 1989.670 ;
        RECT 142.165 1852.000 142.865 1988.000 ;
        RECT 142.165 1850.330 142.865 1850.970 ;
        RECT 0.000 1818.690 142.865 1850.330 ;
      LAYER met4 ;
        RECT 143.265 1819.090 143.595 1990.610 ;
      LAYER met4 ;
        RECT 0.000 1810.360 143.495 1818.690 ;
      LAYER met4 ;
        RECT 143.895 1810.760 146.875 2024.440 ;
      LAYER met4 ;
        RECT 147.275 1989.670 148.255 2024.840 ;
      LAYER met4 ;
        RECT 147.175 1988.000 148.355 1989.270 ;
      LAYER met4 ;
        RECT 147.175 1852.000 148.355 1988.000 ;
      LAYER met4 ;
        RECT 147.175 1850.730 148.355 1852.000 ;
      LAYER met4 ;
        RECT 147.275 1826.065 148.255 1850.330 ;
      LAYER met4 ;
        RECT 148.655 1826.465 151.635 2040.145 ;
        RECT 151.935 2035.090 152.265 2204.000 ;
      LAYER met4 ;
        RECT 152.665 2066.330 153.365 2066.970 ;
      LAYER met4 ;
        RECT 153.765 2066.730 158.415 2204.000 ;
      LAYER met4 ;
        RECT 158.815 2066.330 159.415 2066.970 ;
      LAYER met4 ;
        RECT 159.815 2066.730 163.265 2204.000 ;
      LAYER met4 ;
        RECT 163.665 2066.330 164.265 2066.970 ;
      LAYER met4 ;
        RECT 164.665 2066.730 168.115 2204.000 ;
      LAYER met4 ;
        RECT 168.515 2066.330 169.115 2066.970 ;
      LAYER met4 ;
        RECT 169.515 2066.730 174.165 2204.000 ;
      LAYER met4 ;
        RECT 174.565 2066.330 175.165 2066.970 ;
      LAYER met4 ;
        RECT 175.565 2066.730 180.215 2204.000 ;
        RECT 181.615 2066.970 185.065 2204.000 ;
      LAYER met4 ;
        RECT 180.615 2066.570 181.215 2066.970 ;
        RECT 185.465 2066.570 186.065 2066.970 ;
      LAYER met4 ;
        RECT 186.465 2066.730 191.115 2204.000 ;
      LAYER met4 ;
        RECT 180.615 2066.330 186.065 2066.570 ;
        RECT 191.515 2066.330 192.115 2066.970 ;
      LAYER met4 ;
        RECT 192.515 2066.730 197.965 2204.000 ;
        RECT 3390.035 2151.730 3395.485 2299.000 ;
      LAYER met4 ;
        RECT 3395.885 2151.330 3396.485 2152.035 ;
      LAYER met4 ;
        RECT 3396.885 2151.730 3401.535 2300.270 ;
      LAYER met4 ;
        RECT 3401.935 2151.635 3402.535 2152.035 ;
        RECT 3406.785 2151.635 3407.385 2152.035 ;
      LAYER met4 ;
        RECT 3407.785 2151.730 3412.435 2299.000 ;
      LAYER met4 ;
        RECT 3401.935 2151.330 3407.385 2151.635 ;
        RECT 3412.835 2151.330 3413.435 2152.035 ;
      LAYER met4 ;
        RECT 3413.835 2151.730 3418.485 2299.000 ;
      LAYER met4 ;
        RECT 3418.885 2151.330 3419.485 2152.035 ;
      LAYER met4 ;
        RECT 3419.885 2151.730 3423.335 2299.000 ;
      LAYER met4 ;
        RECT 3423.735 2151.330 3424.335 2152.035 ;
      LAYER met4 ;
        RECT 3424.735 2151.730 3428.185 2299.000 ;
      LAYER met4 ;
        RECT 3428.585 2151.330 3429.185 2152.035 ;
      LAYER met4 ;
        RECT 3429.585 2151.730 3434.235 2299.000 ;
      LAYER met4 ;
        RECT 3434.635 2151.330 3435.335 2152.035 ;
      LAYER met4 ;
        RECT 3435.735 2151.730 3436.065 2299.000 ;
      LAYER met4 ;
        RECT 3390.035 2079.670 3435.965 2151.330 ;
        RECT 198.365 2066.330 199.465 2066.970 ;
        RECT 152.665 2034.690 199.465 2066.330 ;
        RECT 152.035 1991.010 199.465 2034.690 ;
        RECT 147.275 1824.545 151.535 1826.065 ;
        RECT 147.275 1810.360 148.255 1824.545 ;
        RECT 0.000 1808.840 148.255 1810.360 ;
        RECT 0.000 1775.010 143.495 1808.840 ;
        RECT 0.000 1773.670 142.865 1775.010 ;
      LAYER met4 ;
        RECT 0.000 1772.000 24.215 1773.270 ;
      LAYER met4 ;
        RECT 24.615 1772.965 104.600 1773.670 ;
        RECT 0.000 1636.000 104.600 1772.000 ;
      LAYER met4 ;
        RECT 0.000 1634.730 24.215 1636.000 ;
      LAYER met4 ;
        RECT 24.615 1634.330 104.600 1634.970 ;
      LAYER met4 ;
        RECT 105.000 1634.730 129.965 1773.270 ;
      LAYER met4 ;
        RECT 130.365 1772.965 131.065 1773.670 ;
        RECT 130.365 1636.000 131.065 1772.000 ;
        RECT 130.365 1634.330 131.065 1634.970 ;
      LAYER met4 ;
        RECT 131.465 1634.730 135.915 1773.270 ;
      LAYER met4 ;
        RECT 136.315 1772.965 136.915 1773.670 ;
        RECT 136.315 1636.000 136.915 1772.000 ;
        RECT 136.315 1634.330 136.915 1634.970 ;
      LAYER met4 ;
        RECT 137.315 1634.730 141.765 1773.270 ;
      LAYER met4 ;
        RECT 142.165 1772.965 142.865 1773.670 ;
        RECT 142.165 1636.000 142.865 1772.000 ;
        RECT 142.165 1634.330 142.865 1634.970 ;
        RECT 0.000 1602.690 142.865 1634.330 ;
      LAYER met4 ;
        RECT 143.265 1603.090 143.595 1774.610 ;
      LAYER met4 ;
        RECT 0.000 1594.360 143.495 1602.690 ;
      LAYER met4 ;
        RECT 143.895 1594.760 146.875 1808.440 ;
      LAYER met4 ;
        RECT 147.275 1773.670 148.255 1808.840 ;
      LAYER met4 ;
        RECT 147.175 1772.000 148.355 1773.270 ;
      LAYER met4 ;
        RECT 147.175 1636.000 148.355 1772.000 ;
      LAYER met4 ;
        RECT 147.175 1634.730 148.355 1636.000 ;
      LAYER met4 ;
        RECT 147.275 1610.065 148.255 1634.330 ;
      LAYER met4 ;
        RECT 148.655 1610.465 151.635 1824.145 ;
        RECT 151.935 1819.090 152.265 1990.610 ;
      LAYER met4 ;
        RECT 152.665 1989.670 199.465 1991.010 ;
        RECT 152.665 1988.965 153.365 1989.670 ;
        RECT 152.665 1850.330 153.365 1850.970 ;
      LAYER met4 ;
        RECT 153.765 1850.730 158.415 1989.270 ;
      LAYER met4 ;
        RECT 158.815 1988.965 159.415 1989.670 ;
        RECT 158.815 1850.330 159.415 1850.970 ;
      LAYER met4 ;
        RECT 159.815 1850.730 163.265 1989.270 ;
      LAYER met4 ;
        RECT 163.665 1988.965 164.265 1989.670 ;
        RECT 163.665 1850.330 164.265 1850.970 ;
      LAYER met4 ;
        RECT 164.665 1850.730 168.115 1989.270 ;
      LAYER met4 ;
        RECT 168.515 1988.965 169.115 1989.670 ;
        RECT 168.515 1850.330 169.115 1850.970 ;
      LAYER met4 ;
        RECT 169.515 1850.730 174.165 1989.270 ;
      LAYER met4 ;
        RECT 174.565 1988.965 175.165 1989.670 ;
        RECT 180.615 1989.365 186.065 1989.670 ;
        RECT 174.565 1850.330 175.165 1850.970 ;
      LAYER met4 ;
        RECT 175.565 1850.730 180.215 1989.270 ;
      LAYER met4 ;
        RECT 180.615 1988.965 181.215 1989.365 ;
        RECT 185.465 1988.965 186.065 1989.365 ;
      LAYER met4 ;
        RECT 181.615 1850.970 185.065 1988.965 ;
      LAYER met4 ;
        RECT 180.615 1850.570 181.215 1850.970 ;
        RECT 185.465 1850.570 186.065 1850.970 ;
      LAYER met4 ;
        RECT 186.465 1850.730 191.115 1989.270 ;
      LAYER met4 ;
        RECT 191.515 1988.965 192.115 1989.670 ;
        RECT 180.615 1850.330 186.065 1850.570 ;
        RECT 191.515 1850.330 192.115 1850.970 ;
      LAYER met4 ;
        RECT 192.515 1850.730 197.965 1989.270 ;
      LAYER met4 ;
        RECT 198.365 1988.965 199.465 1989.670 ;
        RECT 3388.535 1931.330 3389.635 1932.035 ;
      LAYER met4 ;
        RECT 3390.035 1931.730 3395.485 2079.270 ;
      LAYER met4 ;
        RECT 3395.885 2078.965 3396.485 2079.670 ;
        RECT 3401.935 2079.365 3407.385 2079.670 ;
        RECT 3395.885 1931.330 3396.485 1932.035 ;
      LAYER met4 ;
        RECT 3396.885 1931.730 3401.535 2079.270 ;
      LAYER met4 ;
        RECT 3401.935 2078.965 3402.535 2079.365 ;
        RECT 3406.785 2078.965 3407.385 2079.365 ;
      LAYER met4 ;
        RECT 3402.935 1932.035 3406.385 2078.965 ;
      LAYER met4 ;
        RECT 3401.935 1931.635 3402.535 1932.035 ;
        RECT 3406.785 1931.635 3407.385 1932.035 ;
      LAYER met4 ;
        RECT 3407.785 1931.730 3412.435 2079.270 ;
      LAYER met4 ;
        RECT 3412.835 2078.965 3413.435 2079.670 ;
        RECT 3401.935 1931.330 3407.385 1931.635 ;
        RECT 3412.835 1931.330 3413.435 1932.035 ;
      LAYER met4 ;
        RECT 3413.835 1931.730 3418.485 2079.270 ;
      LAYER met4 ;
        RECT 3418.885 2078.965 3419.485 2079.670 ;
        RECT 3418.885 1931.330 3419.485 1932.035 ;
      LAYER met4 ;
        RECT 3419.885 1931.730 3423.335 2079.270 ;
      LAYER met4 ;
        RECT 3423.735 2078.965 3424.335 2079.670 ;
        RECT 3423.735 1931.330 3424.335 1932.035 ;
      LAYER met4 ;
        RECT 3424.735 1931.730 3428.185 2079.270 ;
      LAYER met4 ;
        RECT 3428.585 2078.965 3429.185 2079.670 ;
        RECT 3428.585 1931.330 3429.185 1932.035 ;
      LAYER met4 ;
        RECT 3429.585 1931.730 3434.235 2079.270 ;
      LAYER met4 ;
        RECT 3434.635 2078.965 3435.335 2079.670 ;
        RECT 3434.635 1931.330 3435.335 1932.035 ;
        RECT 3388.535 1929.990 3435.335 1931.330 ;
      LAYER met4 ;
        RECT 3435.735 1930.390 3436.065 2079.270 ;
      LAYER met4 ;
        RECT 3388.535 1886.310 3435.965 1929.990 ;
        RECT 3388.535 1854.670 3435.335 1886.310 ;
        RECT 3388.535 1854.030 3389.635 1854.670 ;
        RECT 198.365 1850.330 199.465 1850.970 ;
        RECT 152.665 1818.690 199.465 1850.330 ;
        RECT 152.035 1775.010 199.465 1818.690 ;
        RECT 147.275 1608.545 151.535 1610.065 ;
        RECT 147.275 1594.360 148.255 1608.545 ;
        RECT 0.000 1592.840 148.255 1594.360 ;
        RECT 0.000 1559.010 143.495 1592.840 ;
        RECT 0.000 1557.670 142.865 1559.010 ;
      LAYER met4 ;
        RECT 0.000 1556.000 24.215 1557.270 ;
      LAYER met4 ;
        RECT 24.615 1556.965 104.600 1557.670 ;
        RECT 0.000 1420.000 104.600 1556.000 ;
      LAYER met4 ;
        RECT 0.000 1418.730 24.215 1420.000 ;
      LAYER met4 ;
        RECT 24.615 1418.330 104.600 1418.970 ;
      LAYER met4 ;
        RECT 105.000 1418.730 129.965 1557.270 ;
      LAYER met4 ;
        RECT 130.365 1556.965 131.065 1557.670 ;
        RECT 130.365 1420.000 131.065 1556.000 ;
        RECT 130.365 1418.330 131.065 1418.970 ;
      LAYER met4 ;
        RECT 131.465 1418.730 135.915 1557.270 ;
      LAYER met4 ;
        RECT 136.315 1556.965 136.915 1557.670 ;
        RECT 136.315 1420.000 136.915 1556.000 ;
        RECT 136.315 1418.330 136.915 1418.970 ;
      LAYER met4 ;
        RECT 137.315 1418.730 141.765 1557.270 ;
      LAYER met4 ;
        RECT 142.165 1556.965 142.865 1557.670 ;
        RECT 142.165 1420.000 142.865 1556.000 ;
        RECT 142.165 1418.330 142.865 1418.970 ;
        RECT 0.000 1386.690 142.865 1418.330 ;
      LAYER met4 ;
        RECT 143.265 1387.090 143.595 1558.610 ;
      LAYER met4 ;
        RECT 0.000 1378.360 143.495 1386.690 ;
      LAYER met4 ;
        RECT 143.895 1378.760 146.875 1592.440 ;
      LAYER met4 ;
        RECT 147.275 1557.670 148.255 1592.840 ;
      LAYER met4 ;
        RECT 147.175 1556.000 148.355 1557.270 ;
      LAYER met4 ;
        RECT 147.175 1420.000 148.355 1556.000 ;
      LAYER met4 ;
        RECT 147.175 1418.730 148.355 1420.000 ;
      LAYER met4 ;
        RECT 147.275 1394.065 148.255 1418.330 ;
      LAYER met4 ;
        RECT 148.655 1394.465 151.635 1608.145 ;
        RECT 151.935 1603.090 152.265 1774.610 ;
      LAYER met4 ;
        RECT 152.665 1773.670 199.465 1775.010 ;
        RECT 152.665 1772.965 153.365 1773.670 ;
        RECT 152.665 1634.330 153.365 1634.970 ;
      LAYER met4 ;
        RECT 153.765 1634.730 158.415 1773.270 ;
      LAYER met4 ;
        RECT 158.815 1772.965 159.415 1773.670 ;
        RECT 158.815 1634.330 159.415 1634.970 ;
      LAYER met4 ;
        RECT 159.815 1634.730 163.265 1773.270 ;
      LAYER met4 ;
        RECT 163.665 1772.965 164.265 1773.670 ;
        RECT 163.665 1634.330 164.265 1634.970 ;
      LAYER met4 ;
        RECT 164.665 1634.730 168.115 1773.270 ;
      LAYER met4 ;
        RECT 168.515 1772.965 169.115 1773.670 ;
        RECT 168.515 1634.330 169.115 1634.970 ;
      LAYER met4 ;
        RECT 169.515 1634.730 174.165 1773.270 ;
      LAYER met4 ;
        RECT 174.565 1772.965 175.165 1773.670 ;
        RECT 180.615 1773.365 186.065 1773.670 ;
        RECT 174.565 1634.330 175.165 1634.970 ;
      LAYER met4 ;
        RECT 175.565 1634.730 180.215 1773.270 ;
      LAYER met4 ;
        RECT 180.615 1772.965 181.215 1773.365 ;
        RECT 185.465 1772.965 186.065 1773.365 ;
      LAYER met4 ;
        RECT 181.615 1634.970 185.065 1772.965 ;
      LAYER met4 ;
        RECT 180.615 1634.570 181.215 1634.970 ;
        RECT 185.465 1634.570 186.065 1634.970 ;
      LAYER met4 ;
        RECT 186.465 1634.730 191.115 1773.270 ;
      LAYER met4 ;
        RECT 191.515 1772.965 192.115 1773.670 ;
        RECT 180.615 1634.330 186.065 1634.570 ;
        RECT 191.515 1634.330 192.115 1634.970 ;
      LAYER met4 ;
        RECT 192.515 1634.730 197.965 1773.270 ;
      LAYER met4 ;
        RECT 198.365 1772.965 199.465 1773.670 ;
        RECT 3388.535 1705.330 3389.635 1706.035 ;
      LAYER met4 ;
        RECT 3390.035 1705.730 3395.485 1854.270 ;
      LAYER met4 ;
        RECT 3395.885 1854.030 3396.485 1854.670 ;
        RECT 3401.935 1854.430 3407.385 1854.670 ;
        RECT 3395.885 1705.330 3396.485 1706.035 ;
      LAYER met4 ;
        RECT 3396.885 1705.730 3401.535 1854.270 ;
      LAYER met4 ;
        RECT 3401.935 1854.030 3402.535 1854.430 ;
        RECT 3406.785 1854.030 3407.385 1854.430 ;
      LAYER met4 ;
        RECT 3402.935 1706.035 3406.385 1854.030 ;
      LAYER met4 ;
        RECT 3401.935 1705.635 3402.535 1706.035 ;
        RECT 3406.785 1705.635 3407.385 1706.035 ;
      LAYER met4 ;
        RECT 3407.785 1705.730 3412.435 1854.270 ;
      LAYER met4 ;
        RECT 3412.835 1854.030 3413.435 1854.670 ;
        RECT 3401.935 1705.330 3407.385 1705.635 ;
        RECT 3412.835 1705.330 3413.435 1706.035 ;
      LAYER met4 ;
        RECT 3413.835 1705.730 3418.485 1854.270 ;
      LAYER met4 ;
        RECT 3418.885 1854.030 3419.485 1854.670 ;
        RECT 3418.885 1705.330 3419.485 1706.035 ;
      LAYER met4 ;
        RECT 3419.885 1705.730 3423.335 1854.270 ;
      LAYER met4 ;
        RECT 3423.735 1854.030 3424.335 1854.670 ;
        RECT 3423.735 1705.330 3424.335 1706.035 ;
      LAYER met4 ;
        RECT 3424.735 1705.730 3428.185 1854.270 ;
      LAYER met4 ;
        RECT 3428.585 1854.030 3429.185 1854.670 ;
        RECT 3428.585 1705.330 3429.185 1706.035 ;
      LAYER met4 ;
        RECT 3429.585 1705.730 3434.235 1854.270 ;
      LAYER met4 ;
        RECT 3434.635 1854.030 3435.335 1854.670 ;
        RECT 3434.635 1705.330 3435.335 1706.035 ;
        RECT 3388.535 1703.990 3435.335 1705.330 ;
      LAYER met4 ;
        RECT 3435.735 1704.390 3436.065 1885.910 ;
        RECT 3436.365 1880.855 3439.345 2299.000 ;
      LAYER met4 ;
        RECT 3439.645 2153.000 3440.825 2299.000 ;
      LAYER met4 ;
        RECT 3439.645 2151.730 3440.825 2153.000 ;
      LAYER met4 ;
        RECT 3439.745 2079.670 3440.725 2151.330 ;
      LAYER met4 ;
        RECT 3439.645 2078.000 3440.825 2079.270 ;
      LAYER met4 ;
        RECT 3439.645 1933.000 3440.825 2078.000 ;
      LAYER met4 ;
        RECT 3439.645 1931.730 3440.825 1933.000 ;
      LAYER met4 ;
        RECT 3439.745 1896.160 3440.725 1931.330 ;
      LAYER met4 ;
        RECT 3441.125 1896.560 3444.105 2299.000 ;
      LAYER met4 ;
        RECT 3445.135 2153.000 3445.835 2299.000 ;
        RECT 3445.135 2151.330 3445.835 2152.035 ;
      LAYER met4 ;
        RECT 3446.235 2151.730 3450.685 2299.000 ;
      LAYER met4 ;
        RECT 3451.085 2153.000 3451.685 2299.000 ;
        RECT 3451.085 2151.330 3451.685 2152.035 ;
      LAYER met4 ;
        RECT 3452.085 2151.730 3456.535 2299.000 ;
      LAYER met4 ;
        RECT 3456.935 2153.000 3457.635 2299.000 ;
        RECT 3456.935 2151.330 3457.635 2152.035 ;
      LAYER met4 ;
        RECT 3458.035 2151.730 3483.000 2299.000 ;
      LAYER met4 ;
        RECT 3483.400 2153.000 3588.000 2299.000 ;
        RECT 3483.400 2151.330 3563.385 2152.035 ;
      LAYER met4 ;
        RECT 3563.785 2151.730 3588.000 2153.000 ;
      LAYER met4 ;
        RECT 3444.505 2079.670 3588.000 2151.330 ;
      LAYER met4 ;
        RECT 3444.405 1930.390 3444.735 2079.270 ;
      LAYER met4 ;
        RECT 3445.135 2078.965 3445.835 2079.670 ;
        RECT 3445.135 1933.000 3445.835 2078.000 ;
        RECT 3445.135 1931.330 3445.835 1932.035 ;
      LAYER met4 ;
        RECT 3446.235 1931.730 3450.685 2079.270 ;
      LAYER met4 ;
        RECT 3451.085 2078.965 3451.685 2079.670 ;
        RECT 3451.085 1933.000 3451.685 2078.000 ;
        RECT 3451.085 1931.330 3451.685 1932.035 ;
      LAYER met4 ;
        RECT 3452.085 1931.730 3456.535 2079.270 ;
      LAYER met4 ;
        RECT 3456.935 2078.965 3457.635 2079.670 ;
        RECT 3456.935 1933.000 3457.635 2078.000 ;
        RECT 3456.935 1931.330 3457.635 1932.035 ;
      LAYER met4 ;
        RECT 3458.035 1931.730 3483.000 2079.270 ;
      LAYER met4 ;
        RECT 3483.400 2078.965 3563.385 2079.670 ;
      LAYER met4 ;
        RECT 3563.785 2078.000 3588.000 2079.270 ;
      LAYER met4 ;
        RECT 3483.400 1933.000 3588.000 2078.000 ;
        RECT 3483.400 1931.330 3563.385 1932.035 ;
      LAYER met4 ;
        RECT 3563.785 1931.730 3588.000 1933.000 ;
      LAYER met4 ;
        RECT 3445.135 1929.990 3588.000 1931.330 ;
        RECT 3444.505 1896.160 3588.000 1929.990 ;
        RECT 3439.745 1894.640 3588.000 1896.160 ;
        RECT 3439.745 1880.455 3440.725 1894.640 ;
        RECT 3436.465 1878.935 3440.725 1880.455 ;
        RECT 3388.535 1660.310 3435.965 1703.990 ;
        RECT 198.365 1634.330 199.465 1634.970 ;
        RECT 152.665 1602.690 199.465 1634.330 ;
        RECT 3388.535 1628.670 3435.335 1660.310 ;
        RECT 3388.535 1628.030 3389.635 1628.670 ;
        RECT 152.035 1559.010 199.465 1602.690 ;
        RECT 147.275 1392.545 151.535 1394.065 ;
        RECT 147.275 1378.360 148.255 1392.545 ;
        RECT 0.000 1376.840 148.255 1378.360 ;
        RECT 0.000 1343.010 143.495 1376.840 ;
        RECT 0.000 1341.670 142.865 1343.010 ;
      LAYER met4 ;
        RECT 0.000 1340.000 24.215 1341.270 ;
      LAYER met4 ;
        RECT 24.615 1340.965 104.600 1341.670 ;
        RECT 0.000 1204.000 104.600 1340.000 ;
      LAYER met4 ;
        RECT 0.000 1202.730 24.215 1204.000 ;
      LAYER met4 ;
        RECT 24.615 1202.330 104.600 1202.970 ;
      LAYER met4 ;
        RECT 105.000 1202.730 129.965 1341.270 ;
      LAYER met4 ;
        RECT 130.365 1340.965 131.065 1341.670 ;
        RECT 130.365 1204.000 131.065 1340.000 ;
        RECT 130.365 1202.330 131.065 1202.970 ;
      LAYER met4 ;
        RECT 131.465 1202.730 135.915 1341.270 ;
      LAYER met4 ;
        RECT 136.315 1340.965 136.915 1341.670 ;
        RECT 136.315 1204.000 136.915 1340.000 ;
        RECT 136.315 1202.330 136.915 1202.970 ;
      LAYER met4 ;
        RECT 137.315 1202.730 141.765 1341.270 ;
      LAYER met4 ;
        RECT 142.165 1340.965 142.865 1341.670 ;
        RECT 142.165 1204.000 142.865 1340.000 ;
        RECT 142.165 1202.330 142.865 1202.970 ;
        RECT 0.000 1170.690 142.865 1202.330 ;
      LAYER met4 ;
        RECT 143.265 1171.090 143.595 1342.610 ;
      LAYER met4 ;
        RECT 0.000 1162.360 143.495 1170.690 ;
      LAYER met4 ;
        RECT 143.895 1162.760 146.875 1376.440 ;
      LAYER met4 ;
        RECT 147.275 1341.670 148.255 1376.840 ;
      LAYER met4 ;
        RECT 147.175 1340.000 148.355 1341.270 ;
      LAYER met4 ;
        RECT 147.175 1204.000 148.355 1340.000 ;
      LAYER met4 ;
        RECT 147.175 1202.730 148.355 1204.000 ;
      LAYER met4 ;
        RECT 147.275 1178.065 148.255 1202.330 ;
      LAYER met4 ;
        RECT 148.655 1178.465 151.635 1392.145 ;
        RECT 151.935 1387.090 152.265 1558.610 ;
      LAYER met4 ;
        RECT 152.665 1557.670 199.465 1559.010 ;
        RECT 152.665 1556.965 153.365 1557.670 ;
        RECT 152.665 1418.330 153.365 1418.970 ;
      LAYER met4 ;
        RECT 153.765 1418.730 158.415 1557.270 ;
      LAYER met4 ;
        RECT 158.815 1556.965 159.415 1557.670 ;
        RECT 158.815 1418.330 159.415 1418.970 ;
      LAYER met4 ;
        RECT 159.815 1418.730 163.265 1557.270 ;
      LAYER met4 ;
        RECT 163.665 1556.965 164.265 1557.670 ;
        RECT 163.665 1418.330 164.265 1418.970 ;
      LAYER met4 ;
        RECT 164.665 1418.730 168.115 1557.270 ;
      LAYER met4 ;
        RECT 168.515 1556.965 169.115 1557.670 ;
        RECT 168.515 1418.330 169.115 1418.970 ;
      LAYER met4 ;
        RECT 169.515 1418.730 174.165 1557.270 ;
      LAYER met4 ;
        RECT 174.565 1556.965 175.165 1557.670 ;
        RECT 180.615 1557.365 186.065 1557.670 ;
        RECT 174.565 1418.330 175.165 1418.970 ;
      LAYER met4 ;
        RECT 175.565 1418.730 180.215 1557.270 ;
      LAYER met4 ;
        RECT 180.615 1556.965 181.215 1557.365 ;
        RECT 185.465 1556.965 186.065 1557.365 ;
      LAYER met4 ;
        RECT 181.615 1418.970 185.065 1556.965 ;
      LAYER met4 ;
        RECT 180.615 1418.570 181.215 1418.970 ;
        RECT 185.465 1418.570 186.065 1418.970 ;
      LAYER met4 ;
        RECT 186.465 1418.730 191.115 1557.270 ;
      LAYER met4 ;
        RECT 191.515 1556.965 192.115 1557.670 ;
        RECT 180.615 1418.330 186.065 1418.570 ;
        RECT 191.515 1418.330 192.115 1418.970 ;
      LAYER met4 ;
        RECT 192.515 1418.730 197.965 1557.270 ;
      LAYER met4 ;
        RECT 198.365 1556.965 199.465 1557.670 ;
        RECT 3388.535 1480.330 3389.635 1481.035 ;
      LAYER met4 ;
        RECT 3390.035 1480.730 3395.485 1628.270 ;
      LAYER met4 ;
        RECT 3395.885 1628.030 3396.485 1628.670 ;
        RECT 3401.935 1628.430 3407.385 1628.670 ;
        RECT 3395.885 1480.330 3396.485 1481.035 ;
      LAYER met4 ;
        RECT 3396.885 1480.730 3401.535 1628.270 ;
      LAYER met4 ;
        RECT 3401.935 1628.030 3402.535 1628.430 ;
        RECT 3406.785 1628.030 3407.385 1628.430 ;
      LAYER met4 ;
        RECT 3402.935 1481.035 3406.385 1628.030 ;
      LAYER met4 ;
        RECT 3401.935 1480.635 3402.535 1481.035 ;
        RECT 3406.785 1480.635 3407.385 1481.035 ;
      LAYER met4 ;
        RECT 3407.785 1480.730 3412.435 1628.270 ;
      LAYER met4 ;
        RECT 3412.835 1628.030 3413.435 1628.670 ;
        RECT 3401.935 1480.330 3407.385 1480.635 ;
        RECT 3412.835 1480.330 3413.435 1481.035 ;
      LAYER met4 ;
        RECT 3413.835 1480.730 3418.485 1628.270 ;
      LAYER met4 ;
        RECT 3418.885 1628.030 3419.485 1628.670 ;
        RECT 3418.885 1480.330 3419.485 1481.035 ;
      LAYER met4 ;
        RECT 3419.885 1480.730 3423.335 1628.270 ;
      LAYER met4 ;
        RECT 3423.735 1628.030 3424.335 1628.670 ;
        RECT 3423.735 1480.330 3424.335 1481.035 ;
      LAYER met4 ;
        RECT 3424.735 1480.730 3428.185 1628.270 ;
      LAYER met4 ;
        RECT 3428.585 1628.030 3429.185 1628.670 ;
        RECT 3428.585 1480.330 3429.185 1481.035 ;
      LAYER met4 ;
        RECT 3429.585 1480.730 3434.235 1628.270 ;
      LAYER met4 ;
        RECT 3434.635 1628.030 3435.335 1628.670 ;
        RECT 3434.635 1480.330 3435.335 1481.035 ;
        RECT 3388.535 1478.990 3435.335 1480.330 ;
      LAYER met4 ;
        RECT 3435.735 1479.390 3436.065 1659.910 ;
        RECT 3436.365 1654.855 3439.345 1878.535 ;
      LAYER met4 ;
        RECT 3439.745 1854.670 3440.725 1878.935 ;
      LAYER met4 ;
        RECT 3439.645 1853.000 3440.825 1854.270 ;
      LAYER met4 ;
        RECT 3439.645 1707.000 3440.825 1853.000 ;
      LAYER met4 ;
        RECT 3439.645 1705.730 3440.825 1707.000 ;
      LAYER met4 ;
        RECT 3439.745 1670.160 3440.725 1705.330 ;
      LAYER met4 ;
        RECT 3441.125 1670.560 3444.105 1894.240 ;
      LAYER met4 ;
        RECT 3444.505 1886.310 3588.000 1894.640 ;
      LAYER met4 ;
        RECT 3444.405 1704.390 3444.735 1885.910 ;
      LAYER met4 ;
        RECT 3445.135 1854.670 3588.000 1886.310 ;
        RECT 3445.135 1854.030 3445.835 1854.670 ;
        RECT 3445.135 1707.000 3445.835 1853.000 ;
        RECT 3445.135 1705.330 3445.835 1706.035 ;
      LAYER met4 ;
        RECT 3446.235 1705.730 3450.685 1854.270 ;
      LAYER met4 ;
        RECT 3451.085 1854.030 3451.685 1854.670 ;
        RECT 3451.085 1707.000 3451.685 1853.000 ;
        RECT 3451.085 1705.330 3451.685 1706.035 ;
      LAYER met4 ;
        RECT 3452.085 1705.730 3456.535 1854.270 ;
      LAYER met4 ;
        RECT 3456.935 1854.030 3457.635 1854.670 ;
        RECT 3456.935 1707.000 3457.635 1853.000 ;
        RECT 3456.935 1705.330 3457.635 1706.035 ;
      LAYER met4 ;
        RECT 3458.035 1705.730 3483.000 1854.270 ;
      LAYER met4 ;
        RECT 3483.400 1854.030 3563.385 1854.670 ;
      LAYER met4 ;
        RECT 3563.785 1853.000 3588.000 1854.270 ;
      LAYER met4 ;
        RECT 3483.400 1707.000 3588.000 1853.000 ;
        RECT 3483.400 1705.330 3563.385 1706.035 ;
      LAYER met4 ;
        RECT 3563.785 1705.730 3588.000 1707.000 ;
      LAYER met4 ;
        RECT 3445.135 1703.990 3588.000 1705.330 ;
        RECT 3444.505 1670.160 3588.000 1703.990 ;
        RECT 3439.745 1668.640 3588.000 1670.160 ;
        RECT 3439.745 1654.455 3440.725 1668.640 ;
        RECT 3436.465 1652.935 3440.725 1654.455 ;
        RECT 3388.535 1435.310 3435.965 1478.990 ;
        RECT 198.365 1418.330 199.465 1418.970 ;
        RECT 152.665 1386.690 199.465 1418.330 ;
        RECT 3388.535 1403.670 3435.335 1435.310 ;
        RECT 3388.535 1403.030 3389.635 1403.670 ;
        RECT 152.035 1343.010 199.465 1386.690 ;
        RECT 147.275 1176.545 151.535 1178.065 ;
        RECT 147.275 1162.360 148.255 1176.545 ;
        RECT 0.000 1160.840 148.255 1162.360 ;
        RECT 0.000 1127.010 143.495 1160.840 ;
        RECT 0.000 1125.670 142.865 1127.010 ;
      LAYER met4 ;
        RECT 0.000 1124.000 24.215 1125.270 ;
      LAYER met4 ;
        RECT 24.615 1124.965 104.600 1125.670 ;
        RECT 0.000 988.000 104.600 1124.000 ;
      LAYER met4 ;
        RECT 0.000 986.730 24.215 988.000 ;
      LAYER met4 ;
        RECT 24.615 986.330 104.600 986.970 ;
      LAYER met4 ;
        RECT 105.000 986.730 129.965 1125.270 ;
      LAYER met4 ;
        RECT 130.365 1124.965 131.065 1125.670 ;
        RECT 130.365 988.000 131.065 1124.000 ;
        RECT 130.365 986.330 131.065 986.970 ;
      LAYER met4 ;
        RECT 131.465 986.730 135.915 1125.270 ;
      LAYER met4 ;
        RECT 136.315 1124.965 136.915 1125.670 ;
        RECT 136.315 988.000 136.915 1124.000 ;
        RECT 136.315 986.330 136.915 986.970 ;
      LAYER met4 ;
        RECT 137.315 986.730 141.765 1125.270 ;
      LAYER met4 ;
        RECT 142.165 1124.965 142.865 1125.670 ;
        RECT 142.165 988.000 142.865 1124.000 ;
        RECT 142.165 986.330 142.865 986.970 ;
        RECT 0.000 954.690 142.865 986.330 ;
      LAYER met4 ;
        RECT 143.265 955.090 143.595 1126.610 ;
      LAYER met4 ;
        RECT 0.000 946.360 143.495 954.690 ;
      LAYER met4 ;
        RECT 143.895 946.760 146.875 1160.440 ;
      LAYER met4 ;
        RECT 147.275 1125.670 148.255 1160.840 ;
      LAYER met4 ;
        RECT 147.175 1124.000 148.355 1125.270 ;
      LAYER met4 ;
        RECT 147.175 988.000 148.355 1124.000 ;
      LAYER met4 ;
        RECT 147.175 986.730 148.355 988.000 ;
      LAYER met4 ;
        RECT 147.275 962.065 148.255 986.330 ;
      LAYER met4 ;
        RECT 148.655 962.465 151.635 1176.145 ;
        RECT 151.935 1171.090 152.265 1342.610 ;
      LAYER met4 ;
        RECT 152.665 1341.670 199.465 1343.010 ;
        RECT 152.665 1340.965 153.365 1341.670 ;
        RECT 152.665 1202.330 153.365 1202.970 ;
      LAYER met4 ;
        RECT 153.765 1202.730 158.415 1341.270 ;
      LAYER met4 ;
        RECT 158.815 1340.965 159.415 1341.670 ;
        RECT 158.815 1202.330 159.415 1202.970 ;
      LAYER met4 ;
        RECT 159.815 1202.730 163.265 1341.270 ;
      LAYER met4 ;
        RECT 163.665 1340.965 164.265 1341.670 ;
        RECT 163.665 1202.330 164.265 1202.970 ;
      LAYER met4 ;
        RECT 164.665 1202.730 168.115 1341.270 ;
      LAYER met4 ;
        RECT 168.515 1340.965 169.115 1341.670 ;
        RECT 168.515 1202.330 169.115 1202.970 ;
      LAYER met4 ;
        RECT 169.515 1202.730 174.165 1341.270 ;
      LAYER met4 ;
        RECT 174.565 1340.965 175.165 1341.670 ;
        RECT 180.615 1341.365 186.065 1341.670 ;
        RECT 174.565 1202.330 175.165 1202.970 ;
      LAYER met4 ;
        RECT 175.565 1202.730 180.215 1341.270 ;
      LAYER met4 ;
        RECT 180.615 1340.965 181.215 1341.365 ;
        RECT 185.465 1340.965 186.065 1341.365 ;
      LAYER met4 ;
        RECT 181.615 1202.970 185.065 1340.965 ;
      LAYER met4 ;
        RECT 180.615 1202.570 181.215 1202.970 ;
        RECT 185.465 1202.570 186.065 1202.970 ;
      LAYER met4 ;
        RECT 186.465 1202.730 191.115 1341.270 ;
      LAYER met4 ;
        RECT 191.515 1340.965 192.115 1341.670 ;
        RECT 180.615 1202.330 186.065 1202.570 ;
        RECT 191.515 1202.330 192.115 1202.970 ;
      LAYER met4 ;
        RECT 192.515 1202.730 197.965 1341.270 ;
      LAYER met4 ;
        RECT 198.365 1340.965 199.465 1341.670 ;
        RECT 3388.535 1255.330 3389.635 1256.035 ;
      LAYER met4 ;
        RECT 3390.035 1255.730 3395.485 1403.270 ;
      LAYER met4 ;
        RECT 3395.885 1403.030 3396.485 1403.670 ;
        RECT 3401.935 1403.430 3407.385 1403.670 ;
        RECT 3395.885 1255.330 3396.485 1256.035 ;
      LAYER met4 ;
        RECT 3396.885 1255.730 3401.535 1403.270 ;
      LAYER met4 ;
        RECT 3401.935 1403.030 3402.535 1403.430 ;
        RECT 3406.785 1403.030 3407.385 1403.430 ;
      LAYER met4 ;
        RECT 3402.935 1256.035 3406.385 1403.030 ;
      LAYER met4 ;
        RECT 3401.935 1255.635 3402.535 1256.035 ;
        RECT 3406.785 1255.635 3407.385 1256.035 ;
      LAYER met4 ;
        RECT 3407.785 1255.730 3412.435 1403.270 ;
      LAYER met4 ;
        RECT 3412.835 1403.030 3413.435 1403.670 ;
        RECT 3401.935 1255.330 3407.385 1255.635 ;
        RECT 3412.835 1255.330 3413.435 1256.035 ;
      LAYER met4 ;
        RECT 3413.835 1255.730 3418.485 1403.270 ;
      LAYER met4 ;
        RECT 3418.885 1403.030 3419.485 1403.670 ;
        RECT 3418.885 1255.330 3419.485 1256.035 ;
      LAYER met4 ;
        RECT 3419.885 1255.730 3423.335 1403.270 ;
      LAYER met4 ;
        RECT 3423.735 1403.030 3424.335 1403.670 ;
        RECT 3423.735 1255.330 3424.335 1256.035 ;
      LAYER met4 ;
        RECT 3424.735 1255.730 3428.185 1403.270 ;
      LAYER met4 ;
        RECT 3428.585 1403.030 3429.185 1403.670 ;
        RECT 3428.585 1255.330 3429.185 1256.035 ;
      LAYER met4 ;
        RECT 3429.585 1255.730 3434.235 1403.270 ;
      LAYER met4 ;
        RECT 3434.635 1403.030 3435.335 1403.670 ;
        RECT 3434.635 1255.330 3435.335 1256.035 ;
        RECT 3388.535 1253.990 3435.335 1255.330 ;
      LAYER met4 ;
        RECT 3435.735 1254.390 3436.065 1434.910 ;
        RECT 3436.365 1429.855 3439.345 1652.535 ;
      LAYER met4 ;
        RECT 3439.745 1628.670 3440.725 1652.935 ;
      LAYER met4 ;
        RECT 3439.645 1627.000 3440.825 1628.270 ;
      LAYER met4 ;
        RECT 3439.645 1482.000 3440.825 1627.000 ;
      LAYER met4 ;
        RECT 3439.645 1480.730 3440.825 1482.000 ;
      LAYER met4 ;
        RECT 3439.745 1445.160 3440.725 1480.330 ;
      LAYER met4 ;
        RECT 3441.125 1445.560 3444.105 1668.240 ;
      LAYER met4 ;
        RECT 3444.505 1660.310 3588.000 1668.640 ;
      LAYER met4 ;
        RECT 3444.405 1479.390 3444.735 1659.910 ;
      LAYER met4 ;
        RECT 3445.135 1628.670 3588.000 1660.310 ;
        RECT 3445.135 1628.030 3445.835 1628.670 ;
        RECT 3445.135 1482.000 3445.835 1627.000 ;
        RECT 3445.135 1480.330 3445.835 1481.035 ;
      LAYER met4 ;
        RECT 3446.235 1480.730 3450.685 1628.270 ;
      LAYER met4 ;
        RECT 3451.085 1628.030 3451.685 1628.670 ;
        RECT 3451.085 1482.000 3451.685 1627.000 ;
        RECT 3451.085 1480.330 3451.685 1481.035 ;
      LAYER met4 ;
        RECT 3452.085 1480.730 3456.535 1628.270 ;
      LAYER met4 ;
        RECT 3456.935 1628.030 3457.635 1628.670 ;
        RECT 3456.935 1482.000 3457.635 1627.000 ;
        RECT 3456.935 1480.330 3457.635 1481.035 ;
      LAYER met4 ;
        RECT 3458.035 1480.730 3483.000 1628.270 ;
      LAYER met4 ;
        RECT 3483.400 1628.030 3563.385 1628.670 ;
      LAYER met4 ;
        RECT 3563.785 1627.000 3588.000 1628.270 ;
      LAYER met4 ;
        RECT 3483.400 1482.000 3588.000 1627.000 ;
        RECT 3483.400 1480.330 3563.385 1481.035 ;
      LAYER met4 ;
        RECT 3563.785 1480.730 3588.000 1482.000 ;
      LAYER met4 ;
        RECT 3445.135 1478.990 3588.000 1480.330 ;
        RECT 3444.505 1445.160 3588.000 1478.990 ;
        RECT 3439.745 1443.640 3588.000 1445.160 ;
        RECT 3439.745 1429.455 3440.725 1443.640 ;
        RECT 3436.465 1427.935 3440.725 1429.455 ;
        RECT 3388.535 1210.310 3435.965 1253.990 ;
        RECT 198.365 1202.330 199.465 1202.970 ;
        RECT 152.665 1170.690 199.465 1202.330 ;
        RECT 3388.535 1178.670 3435.335 1210.310 ;
        RECT 3388.535 1178.030 3389.635 1178.670 ;
        RECT 152.035 1127.010 199.465 1170.690 ;
        RECT 147.275 960.545 151.535 962.065 ;
        RECT 147.275 946.360 148.255 960.545 ;
        RECT 0.000 944.840 148.255 946.360 ;
        RECT 0.000 911.010 143.495 944.840 ;
        RECT 0.000 909.670 142.865 911.010 ;
      LAYER met4 ;
        RECT 0.000 908.000 24.215 909.270 ;
      LAYER met4 ;
        RECT 24.615 908.965 104.600 909.670 ;
        RECT 0.000 631.000 104.600 908.000 ;
        RECT 0.000 626.000 24.215 631.000 ;
      LAYER met4 ;
        RECT 0.000 624.730 24.215 626.000 ;
      LAYER met4 ;
        RECT 24.615 624.330 104.600 625.035 ;
      LAYER met4 ;
        RECT 105.000 624.730 129.965 909.270 ;
      LAYER met4 ;
        RECT 130.365 908.965 131.065 909.670 ;
        RECT 130.365 631.000 131.065 908.000 ;
        RECT 130.365 624.330 131.065 625.035 ;
      LAYER met4 ;
        RECT 131.465 624.730 135.915 909.270 ;
      LAYER met4 ;
        RECT 136.315 908.965 136.915 909.670 ;
        RECT 136.315 631.000 136.915 908.000 ;
        RECT 136.315 624.330 136.915 625.035 ;
      LAYER met4 ;
        RECT 137.315 624.730 141.765 909.270 ;
      LAYER met4 ;
        RECT 142.165 908.965 142.865 909.670 ;
        RECT 142.165 631.000 142.865 908.000 ;
      LAYER met4 ;
        RECT 143.265 631.000 143.595 910.610 ;
      LAYER met4 ;
        RECT 142.165 624.330 142.865 625.035 ;
        RECT 0.000 552.670 142.865 624.330 ;
      LAYER met4 ;
        RECT 0.000 551.000 24.215 552.270 ;
      LAYER met4 ;
        RECT 24.615 551.965 104.600 552.670 ;
        RECT 0.000 415.000 104.600 551.000 ;
      LAYER met4 ;
        RECT 0.000 413.730 24.215 415.000 ;
      LAYER met4 ;
        RECT 24.615 413.330 104.600 415.000 ;
      LAYER met4 ;
        RECT 105.000 413.730 129.965 552.270 ;
      LAYER met4 ;
        RECT 130.365 551.965 131.065 552.670 ;
        RECT 130.365 413.330 131.065 551.000 ;
      LAYER met4 ;
        RECT 131.465 413.730 135.915 552.270 ;
      LAYER met4 ;
        RECT 136.315 551.965 136.915 552.670 ;
        RECT 136.315 413.330 136.915 551.000 ;
      LAYER met4 ;
        RECT 137.315 413.730 141.765 552.270 ;
      LAYER met4 ;
        RECT 142.165 551.965 142.865 552.670 ;
        RECT 142.165 413.330 142.865 551.000 ;
        RECT 0.000 341.670 142.865 413.330 ;
      LAYER met4 ;
        RECT 0.000 340.000 24.215 341.270 ;
      LAYER met4 ;
        RECT 24.615 340.965 104.600 341.670 ;
        RECT 0.000 204.000 104.600 340.000 ;
      LAYER met4 ;
        RECT 0.000 202.730 24.215 204.000 ;
      LAYER met4 ;
        RECT 24.615 202.330 104.600 202.745 ;
        RECT 0.000 201.745 104.600 202.330 ;
      LAYER met4 ;
        RECT 105.000 202.145 129.965 341.270 ;
      LAYER met4 ;
        RECT 130.365 340.965 131.065 341.670 ;
        RECT 130.365 204.000 131.065 340.000 ;
        RECT 130.365 202.330 131.065 202.745 ;
      LAYER met4 ;
        RECT 131.465 202.730 135.915 341.270 ;
      LAYER met4 ;
        RECT 136.315 340.965 136.915 341.670 ;
        RECT 136.315 204.000 136.915 340.000 ;
        RECT 136.315 202.330 136.915 202.745 ;
      LAYER met4 ;
        RECT 137.315 202.730 141.765 341.270 ;
      LAYER met4 ;
        RECT 142.165 340.965 142.865 341.670 ;
        RECT 142.165 204.000 142.865 340.000 ;
        RECT 142.165 202.330 142.865 202.745 ;
        RECT 130.365 201.745 142.865 202.330 ;
        RECT 0.000 176.425 142.865 201.745 ;
      LAYER met4 ;
        RECT 143.265 176.825 143.595 626.000 ;
        RECT 143.895 177.090 146.875 944.440 ;
      LAYER met4 ;
        RECT 147.275 909.670 148.255 944.840 ;
      LAYER met4 ;
        RECT 147.175 908.000 148.355 909.270 ;
      LAYER met4 ;
        RECT 147.175 631.000 148.355 908.000 ;
      LAYER met4 ;
        RECT 147.175 624.730 148.355 626.000 ;
      LAYER met4 ;
        RECT 147.275 552.670 148.255 624.330 ;
      LAYER met4 ;
        RECT 147.175 551.000 148.355 552.270 ;
      LAYER met4 ;
        RECT 147.175 415.000 148.355 551.000 ;
      LAYER met4 ;
        RECT 147.175 413.730 148.355 415.000 ;
      LAYER met4 ;
        RECT 147.275 341.670 148.255 413.330 ;
      LAYER met4 ;
        RECT 147.175 340.000 148.355 341.270 ;
      LAYER met4 ;
        RECT 147.175 204.000 148.355 340.000 ;
      LAYER met4 ;
        RECT 147.175 182.445 148.355 204.000 ;
        RECT 148.655 183.125 151.635 960.145 ;
        RECT 151.935 955.090 152.265 1126.610 ;
      LAYER met4 ;
        RECT 152.665 1125.670 199.465 1127.010 ;
        RECT 152.665 1124.965 153.365 1125.670 ;
        RECT 152.665 986.330 153.365 986.970 ;
      LAYER met4 ;
        RECT 153.765 986.730 158.415 1125.270 ;
      LAYER met4 ;
        RECT 158.815 1124.965 159.415 1125.670 ;
        RECT 158.815 986.330 159.415 986.970 ;
      LAYER met4 ;
        RECT 159.815 986.730 163.265 1125.270 ;
      LAYER met4 ;
        RECT 163.665 1124.965 164.265 1125.670 ;
        RECT 163.665 986.330 164.265 986.970 ;
      LAYER met4 ;
        RECT 164.665 986.730 168.115 1125.270 ;
      LAYER met4 ;
        RECT 168.515 1124.965 169.115 1125.670 ;
        RECT 168.515 986.330 169.115 986.970 ;
      LAYER met4 ;
        RECT 169.515 986.730 174.165 1125.270 ;
      LAYER met4 ;
        RECT 174.565 1124.965 175.165 1125.670 ;
        RECT 180.615 1125.365 186.065 1125.670 ;
        RECT 174.565 986.330 175.165 986.970 ;
      LAYER met4 ;
        RECT 175.565 986.730 180.215 1125.270 ;
      LAYER met4 ;
        RECT 180.615 1124.965 181.215 1125.365 ;
        RECT 185.465 1124.965 186.065 1125.365 ;
      LAYER met4 ;
        RECT 181.615 986.970 185.065 1124.965 ;
      LAYER met4 ;
        RECT 180.615 986.570 181.215 986.970 ;
        RECT 185.465 986.570 186.065 986.970 ;
      LAYER met4 ;
        RECT 186.465 986.730 191.115 1125.270 ;
      LAYER met4 ;
        RECT 191.515 1124.965 192.115 1125.670 ;
        RECT 180.615 986.330 186.065 986.570 ;
        RECT 191.515 986.330 192.115 986.970 ;
      LAYER met4 ;
        RECT 192.515 986.730 197.965 1125.270 ;
      LAYER met4 ;
        RECT 198.365 1124.965 199.465 1125.670 ;
        RECT 3388.535 1029.330 3389.635 1030.035 ;
      LAYER met4 ;
        RECT 3390.035 1029.730 3395.485 1178.270 ;
      LAYER met4 ;
        RECT 3395.885 1178.030 3396.485 1178.670 ;
        RECT 3401.935 1178.430 3407.385 1178.670 ;
        RECT 3395.885 1029.330 3396.485 1030.035 ;
      LAYER met4 ;
        RECT 3396.885 1029.730 3401.535 1178.270 ;
      LAYER met4 ;
        RECT 3401.935 1178.030 3402.535 1178.430 ;
        RECT 3406.785 1178.030 3407.385 1178.430 ;
      LAYER met4 ;
        RECT 3402.935 1030.035 3406.385 1178.030 ;
      LAYER met4 ;
        RECT 3401.935 1029.635 3402.535 1030.035 ;
        RECT 3406.785 1029.635 3407.385 1030.035 ;
      LAYER met4 ;
        RECT 3407.785 1029.730 3412.435 1178.270 ;
      LAYER met4 ;
        RECT 3412.835 1178.030 3413.435 1178.670 ;
        RECT 3401.935 1029.330 3407.385 1029.635 ;
        RECT 3412.835 1029.330 3413.435 1030.035 ;
      LAYER met4 ;
        RECT 3413.835 1029.730 3418.485 1178.270 ;
      LAYER met4 ;
        RECT 3418.885 1178.030 3419.485 1178.670 ;
        RECT 3418.885 1029.330 3419.485 1030.035 ;
      LAYER met4 ;
        RECT 3419.885 1029.730 3423.335 1178.270 ;
      LAYER met4 ;
        RECT 3423.735 1178.030 3424.335 1178.670 ;
        RECT 3423.735 1029.330 3424.335 1030.035 ;
      LAYER met4 ;
        RECT 3424.735 1029.730 3428.185 1178.270 ;
      LAYER met4 ;
        RECT 3428.585 1178.030 3429.185 1178.670 ;
        RECT 3428.585 1029.330 3429.185 1030.035 ;
      LAYER met4 ;
        RECT 3429.585 1029.730 3434.235 1178.270 ;
      LAYER met4 ;
        RECT 3434.635 1178.030 3435.335 1178.670 ;
        RECT 3434.635 1029.330 3435.335 1030.035 ;
        RECT 3388.535 1027.990 3435.335 1029.330 ;
      LAYER met4 ;
        RECT 3435.735 1028.390 3436.065 1209.910 ;
        RECT 3436.365 1204.855 3439.345 1427.535 ;
      LAYER met4 ;
        RECT 3439.745 1403.670 3440.725 1427.935 ;
      LAYER met4 ;
        RECT 3439.645 1402.000 3440.825 1403.270 ;
      LAYER met4 ;
        RECT 3439.645 1257.000 3440.825 1402.000 ;
      LAYER met4 ;
        RECT 3439.645 1255.730 3440.825 1257.000 ;
      LAYER met4 ;
        RECT 3439.745 1220.160 3440.725 1255.330 ;
      LAYER met4 ;
        RECT 3441.125 1220.560 3444.105 1443.240 ;
      LAYER met4 ;
        RECT 3444.505 1435.310 3588.000 1443.640 ;
      LAYER met4 ;
        RECT 3444.405 1254.390 3444.735 1434.910 ;
      LAYER met4 ;
        RECT 3445.135 1403.670 3588.000 1435.310 ;
        RECT 3445.135 1403.030 3445.835 1403.670 ;
        RECT 3445.135 1257.000 3445.835 1402.000 ;
        RECT 3445.135 1255.330 3445.835 1256.035 ;
      LAYER met4 ;
        RECT 3446.235 1255.730 3450.685 1403.270 ;
      LAYER met4 ;
        RECT 3451.085 1403.030 3451.685 1403.670 ;
        RECT 3451.085 1257.000 3451.685 1402.000 ;
        RECT 3451.085 1255.330 3451.685 1256.035 ;
      LAYER met4 ;
        RECT 3452.085 1255.730 3456.535 1403.270 ;
      LAYER met4 ;
        RECT 3456.935 1403.030 3457.635 1403.670 ;
        RECT 3456.935 1257.000 3457.635 1402.000 ;
        RECT 3456.935 1255.330 3457.635 1256.035 ;
      LAYER met4 ;
        RECT 3458.035 1255.730 3483.000 1403.270 ;
      LAYER met4 ;
        RECT 3483.400 1403.030 3563.385 1403.670 ;
      LAYER met4 ;
        RECT 3563.785 1402.000 3588.000 1403.270 ;
      LAYER met4 ;
        RECT 3483.400 1257.000 3588.000 1402.000 ;
        RECT 3483.400 1255.330 3563.385 1256.035 ;
      LAYER met4 ;
        RECT 3563.785 1255.730 3588.000 1257.000 ;
      LAYER met4 ;
        RECT 3445.135 1253.990 3588.000 1255.330 ;
        RECT 3444.505 1220.160 3588.000 1253.990 ;
        RECT 3439.745 1218.640 3588.000 1220.160 ;
        RECT 3439.745 1204.455 3440.725 1218.640 ;
        RECT 3436.465 1202.935 3440.725 1204.455 ;
        RECT 198.365 986.330 199.465 986.970 ;
        RECT 152.665 954.690 199.465 986.330 ;
        RECT 152.035 911.010 199.465 954.690 ;
        RECT 3388.535 984.310 3435.965 1027.990 ;
        RECT 3388.535 952.670 3435.335 984.310 ;
        RECT 3388.535 952.030 3389.635 952.670 ;
      LAYER met4 ;
        RECT 151.935 631.000 152.265 910.610 ;
      LAYER met4 ;
        RECT 152.665 909.670 199.465 911.010 ;
        RECT 152.665 908.965 153.365 909.670 ;
        RECT 148.755 182.045 151.535 182.725 ;
        RECT 147.275 180.025 151.535 182.045 ;
      LAYER met4 ;
        RECT 151.935 180.425 152.265 626.000 ;
      LAYER met4 ;
        RECT 152.665 624.330 153.365 625.035 ;
      LAYER met4 ;
        RECT 153.765 624.730 158.415 909.270 ;
      LAYER met4 ;
        RECT 158.815 908.965 159.415 909.670 ;
      LAYER met4 ;
        RECT 159.815 631.000 163.265 909.270 ;
      LAYER met4 ;
        RECT 163.665 908.965 164.265 909.670 ;
        RECT 158.815 624.330 159.415 625.035 ;
      LAYER met4 ;
        RECT 159.815 624.730 163.265 626.000 ;
      LAYER met4 ;
        RECT 163.665 624.330 164.265 625.035 ;
      LAYER met4 ;
        RECT 164.665 624.730 168.115 909.270 ;
      LAYER met4 ;
        RECT 168.515 908.965 169.115 909.670 ;
        RECT 168.515 624.330 169.115 625.035 ;
      LAYER met4 ;
        RECT 169.515 624.730 174.165 909.270 ;
      LAYER met4 ;
        RECT 174.565 908.965 175.165 909.670 ;
        RECT 180.615 909.365 186.065 909.670 ;
        RECT 174.565 624.330 175.165 625.035 ;
      LAYER met4 ;
        RECT 175.565 624.730 180.215 909.270 ;
      LAYER met4 ;
        RECT 180.615 908.965 181.215 909.365 ;
        RECT 185.465 908.965 186.065 909.365 ;
      LAYER met4 ;
        RECT 181.615 631.000 185.065 908.965 ;
        RECT 181.615 625.035 185.065 626.000 ;
      LAYER met4 ;
        RECT 180.615 624.635 181.215 625.035 ;
        RECT 185.465 624.635 186.065 625.035 ;
      LAYER met4 ;
        RECT 186.465 624.730 191.115 909.270 ;
      LAYER met4 ;
        RECT 191.515 908.965 192.115 909.670 ;
        RECT 180.615 624.330 186.065 624.635 ;
        RECT 191.515 624.330 192.115 625.035 ;
      LAYER met4 ;
        RECT 192.515 624.730 197.965 909.270 ;
      LAYER met4 ;
        RECT 198.365 908.965 199.465 909.670 ;
        RECT 3388.535 804.330 3389.635 805.035 ;
      LAYER met4 ;
        RECT 3390.035 804.730 3395.485 952.270 ;
      LAYER met4 ;
        RECT 3395.885 952.030 3396.485 952.670 ;
        RECT 3401.935 952.430 3407.385 952.670 ;
        RECT 3395.885 804.330 3396.485 805.035 ;
      LAYER met4 ;
        RECT 3396.885 804.730 3401.535 952.270 ;
      LAYER met4 ;
        RECT 3401.935 952.030 3402.535 952.430 ;
        RECT 3406.785 952.030 3407.385 952.430 ;
      LAYER met4 ;
        RECT 3402.935 805.035 3406.385 952.030 ;
      LAYER met4 ;
        RECT 3401.935 804.635 3402.535 805.035 ;
        RECT 3406.785 804.635 3407.385 805.035 ;
      LAYER met4 ;
        RECT 3407.785 804.730 3412.435 952.270 ;
      LAYER met4 ;
        RECT 3412.835 952.030 3413.435 952.670 ;
        RECT 3401.935 804.330 3407.385 804.635 ;
        RECT 3412.835 804.330 3413.435 805.035 ;
      LAYER met4 ;
        RECT 3413.835 804.730 3418.485 952.270 ;
      LAYER met4 ;
        RECT 3418.885 952.030 3419.485 952.670 ;
        RECT 3418.885 804.330 3419.485 805.035 ;
      LAYER met4 ;
        RECT 3419.885 804.730 3423.335 952.270 ;
      LAYER met4 ;
        RECT 3423.735 952.030 3424.335 952.670 ;
        RECT 3423.735 804.330 3424.335 805.035 ;
      LAYER met4 ;
        RECT 3424.735 804.730 3428.185 952.270 ;
      LAYER met4 ;
        RECT 3428.585 952.030 3429.185 952.670 ;
        RECT 3428.585 804.330 3429.185 805.035 ;
      LAYER met4 ;
        RECT 3429.585 804.730 3434.235 952.270 ;
      LAYER met4 ;
        RECT 3434.635 952.030 3435.335 952.670 ;
        RECT 3434.635 804.330 3435.335 805.035 ;
        RECT 3388.535 802.990 3435.335 804.330 ;
      LAYER met4 ;
        RECT 3435.735 803.390 3436.065 983.910 ;
        RECT 3436.365 978.855 3439.345 1202.535 ;
      LAYER met4 ;
        RECT 3439.745 1178.670 3440.725 1202.935 ;
      LAYER met4 ;
        RECT 3439.645 1177.000 3440.825 1178.270 ;
      LAYER met4 ;
        RECT 3439.645 1031.000 3440.825 1177.000 ;
      LAYER met4 ;
        RECT 3439.645 1029.730 3440.825 1031.000 ;
      LAYER met4 ;
        RECT 3439.745 994.160 3440.725 1029.330 ;
      LAYER met4 ;
        RECT 3441.125 994.560 3444.105 1218.240 ;
      LAYER met4 ;
        RECT 3444.505 1210.310 3588.000 1218.640 ;
      LAYER met4 ;
        RECT 3444.405 1028.390 3444.735 1209.910 ;
      LAYER met4 ;
        RECT 3445.135 1178.670 3588.000 1210.310 ;
        RECT 3445.135 1178.030 3445.835 1178.670 ;
        RECT 3445.135 1031.000 3445.835 1177.000 ;
        RECT 3445.135 1029.330 3445.835 1030.035 ;
      LAYER met4 ;
        RECT 3446.235 1029.730 3450.685 1178.270 ;
      LAYER met4 ;
        RECT 3451.085 1178.030 3451.685 1178.670 ;
        RECT 3451.085 1031.000 3451.685 1177.000 ;
        RECT 3451.085 1029.330 3451.685 1030.035 ;
      LAYER met4 ;
        RECT 3452.085 1029.730 3456.535 1178.270 ;
      LAYER met4 ;
        RECT 3456.935 1178.030 3457.635 1178.670 ;
        RECT 3456.935 1031.000 3457.635 1177.000 ;
        RECT 3456.935 1029.330 3457.635 1030.035 ;
      LAYER met4 ;
        RECT 3458.035 1029.730 3483.000 1178.270 ;
      LAYER met4 ;
        RECT 3483.400 1178.030 3563.385 1178.670 ;
      LAYER met4 ;
        RECT 3563.785 1177.000 3588.000 1178.270 ;
      LAYER met4 ;
        RECT 3483.400 1031.000 3588.000 1177.000 ;
        RECT 3483.400 1029.330 3563.385 1030.035 ;
      LAYER met4 ;
        RECT 3563.785 1029.730 3588.000 1031.000 ;
      LAYER met4 ;
        RECT 3445.135 1027.990 3588.000 1029.330 ;
        RECT 3444.505 994.160 3588.000 1027.990 ;
        RECT 3439.745 992.640 3588.000 994.160 ;
        RECT 3439.745 978.455 3440.725 992.640 ;
        RECT 3436.465 976.935 3440.725 978.455 ;
        RECT 3388.535 759.310 3435.965 802.990 ;
        RECT 3388.535 727.670 3435.335 759.310 ;
        RECT 3388.535 727.030 3389.635 727.670 ;
        RECT 152.665 552.670 197.965 624.330 ;
        RECT 3388.535 578.330 3389.635 579.035 ;
      LAYER met4 ;
        RECT 3390.035 578.730 3395.485 727.270 ;
      LAYER met4 ;
        RECT 3395.885 727.030 3396.485 727.670 ;
        RECT 3401.935 727.430 3407.385 727.670 ;
        RECT 3395.885 578.330 3396.485 579.035 ;
      LAYER met4 ;
        RECT 3396.885 578.730 3401.535 727.270 ;
      LAYER met4 ;
        RECT 3401.935 727.030 3402.535 727.430 ;
        RECT 3406.785 727.030 3407.385 727.430 ;
      LAYER met4 ;
        RECT 3402.935 579.035 3406.385 727.030 ;
      LAYER met4 ;
        RECT 3401.935 578.635 3402.535 579.035 ;
        RECT 3406.785 578.635 3407.385 579.035 ;
      LAYER met4 ;
        RECT 3407.785 578.730 3412.435 727.270 ;
      LAYER met4 ;
        RECT 3412.835 727.030 3413.435 727.670 ;
        RECT 3401.935 578.330 3407.385 578.635 ;
        RECT 3412.835 578.330 3413.435 579.035 ;
      LAYER met4 ;
        RECT 3413.835 578.730 3418.485 727.270 ;
      LAYER met4 ;
        RECT 3418.885 727.030 3419.485 727.670 ;
        RECT 3418.885 578.330 3419.485 579.035 ;
      LAYER met4 ;
        RECT 3419.885 578.730 3423.335 727.270 ;
      LAYER met4 ;
        RECT 3423.735 727.030 3424.335 727.670 ;
        RECT 3423.735 578.330 3424.335 579.035 ;
      LAYER met4 ;
        RECT 3424.735 578.730 3428.185 727.270 ;
      LAYER met4 ;
        RECT 3428.585 727.030 3429.185 727.670 ;
        RECT 3428.585 578.330 3429.185 579.035 ;
      LAYER met4 ;
        RECT 3429.585 578.730 3434.235 727.270 ;
      LAYER met4 ;
        RECT 3434.635 727.030 3435.335 727.670 ;
        RECT 3434.635 578.330 3435.335 579.035 ;
        RECT 3388.535 576.990 3435.335 578.330 ;
      LAYER met4 ;
        RECT 3435.735 577.390 3436.065 758.910 ;
        RECT 3436.365 753.855 3439.345 976.535 ;
      LAYER met4 ;
        RECT 3439.745 952.670 3440.725 976.935 ;
      LAYER met4 ;
        RECT 3439.645 951.000 3440.825 952.270 ;
      LAYER met4 ;
        RECT 3439.645 806.000 3440.825 951.000 ;
      LAYER met4 ;
        RECT 3439.645 804.730 3440.825 806.000 ;
      LAYER met4 ;
        RECT 3439.745 769.160 3440.725 804.330 ;
      LAYER met4 ;
        RECT 3441.125 769.560 3444.105 992.240 ;
      LAYER met4 ;
        RECT 3444.505 984.310 3588.000 992.640 ;
      LAYER met4 ;
        RECT 3444.405 803.390 3444.735 983.910 ;
      LAYER met4 ;
        RECT 3445.135 952.670 3588.000 984.310 ;
        RECT 3445.135 952.030 3445.835 952.670 ;
        RECT 3445.135 806.000 3445.835 951.000 ;
        RECT 3445.135 804.330 3445.835 805.035 ;
      LAYER met4 ;
        RECT 3446.235 804.730 3450.685 952.270 ;
      LAYER met4 ;
        RECT 3451.085 952.030 3451.685 952.670 ;
        RECT 3451.085 806.000 3451.685 951.000 ;
        RECT 3451.085 804.330 3451.685 805.035 ;
      LAYER met4 ;
        RECT 3452.085 804.730 3456.535 952.270 ;
      LAYER met4 ;
        RECT 3456.935 952.030 3457.635 952.670 ;
        RECT 3456.935 806.000 3457.635 951.000 ;
        RECT 3456.935 804.330 3457.635 805.035 ;
      LAYER met4 ;
        RECT 3458.035 804.730 3483.000 952.270 ;
      LAYER met4 ;
        RECT 3483.400 952.030 3563.385 952.670 ;
      LAYER met4 ;
        RECT 3563.785 951.000 3588.000 952.270 ;
      LAYER met4 ;
        RECT 3483.400 806.000 3588.000 951.000 ;
        RECT 3483.400 804.330 3563.385 805.035 ;
      LAYER met4 ;
        RECT 3563.785 804.730 3588.000 806.000 ;
      LAYER met4 ;
        RECT 3445.135 802.990 3588.000 804.330 ;
        RECT 3444.505 769.160 3588.000 802.990 ;
        RECT 3439.745 767.640 3588.000 769.160 ;
        RECT 3439.745 753.455 3440.725 767.640 ;
        RECT 3436.465 751.935 3440.725 753.455 ;
        RECT 152.665 551.965 153.365 552.670 ;
        RECT 152.665 413.330 153.365 415.000 ;
      LAYER met4 ;
        RECT 153.765 413.730 158.415 552.270 ;
      LAYER met4 ;
        RECT 158.815 551.965 159.415 552.670 ;
        RECT 158.815 413.330 159.415 415.000 ;
      LAYER met4 ;
        RECT 159.815 413.730 163.265 552.270 ;
      LAYER met4 ;
        RECT 163.665 551.965 164.265 552.670 ;
        RECT 163.665 413.330 164.265 415.000 ;
      LAYER met4 ;
        RECT 164.665 413.730 168.115 552.270 ;
      LAYER met4 ;
        RECT 168.515 551.965 169.115 552.670 ;
        RECT 168.515 413.330 169.115 415.000 ;
      LAYER met4 ;
        RECT 169.515 413.730 174.165 552.270 ;
      LAYER met4 ;
        RECT 174.565 551.965 175.165 552.670 ;
        RECT 180.615 552.365 186.065 552.670 ;
        RECT 174.565 413.330 175.165 415.000 ;
      LAYER met4 ;
        RECT 175.565 413.730 180.215 552.270 ;
      LAYER met4 ;
        RECT 180.615 551.965 181.215 552.365 ;
        RECT 185.465 551.965 186.065 552.365 ;
        RECT 180.615 413.635 181.215 415.000 ;
      LAYER met4 ;
        RECT 181.615 414.035 185.065 551.965 ;
      LAYER met4 ;
        RECT 185.465 413.635 186.065 415.000 ;
      LAYER met4 ;
        RECT 186.465 413.730 191.115 552.270 ;
      LAYER met4 ;
        RECT 191.515 551.965 192.115 552.670 ;
        RECT 180.615 413.330 186.065 413.635 ;
        RECT 191.515 413.330 192.115 415.000 ;
      LAYER met4 ;
        RECT 192.515 413.730 197.965 552.270 ;
      LAYER met4 ;
        RECT 3388.535 533.310 3435.965 576.990 ;
        RECT 3388.535 501.670 3435.335 533.310 ;
        RECT 3388.535 501.030 3389.635 501.670 ;
        RECT 152.665 341.670 197.965 413.330 ;
        RECT 152.665 340.965 153.365 341.670 ;
        RECT 152.665 202.330 153.365 202.745 ;
      LAYER met4 ;
        RECT 153.765 202.730 158.415 341.270 ;
      LAYER met4 ;
        RECT 158.815 340.965 159.415 341.670 ;
        RECT 158.815 202.330 159.415 202.745 ;
      LAYER met4 ;
        RECT 159.815 202.730 163.265 341.270 ;
      LAYER met4 ;
        RECT 163.665 340.965 164.265 341.670 ;
        RECT 163.665 202.330 164.265 202.745 ;
      LAYER met4 ;
        RECT 164.665 202.730 168.115 341.270 ;
      LAYER met4 ;
        RECT 168.515 340.965 169.115 341.670 ;
        RECT 168.515 202.330 169.115 202.745 ;
      LAYER met4 ;
        RECT 169.515 202.730 174.165 341.270 ;
      LAYER met4 ;
        RECT 174.565 340.965 175.165 341.670 ;
        RECT 180.615 341.365 186.065 341.670 ;
        RECT 174.565 202.330 175.165 202.745 ;
      LAYER met4 ;
        RECT 175.565 202.730 180.215 341.270 ;
      LAYER met4 ;
        RECT 180.615 340.965 181.215 341.365 ;
        RECT 185.465 340.965 186.065 341.365 ;
      LAYER met4 ;
        RECT 181.615 202.745 185.065 340.965 ;
      LAYER met4 ;
        RECT 180.615 202.345 181.215 202.745 ;
        RECT 185.465 202.345 186.065 202.745 ;
      LAYER met4 ;
        RECT 186.465 202.730 191.115 341.270 ;
      LAYER met4 ;
        RECT 191.515 340.965 192.115 341.670 ;
        RECT 180.615 202.330 186.065 202.345 ;
        RECT 191.515 202.330 192.115 202.745 ;
      LAYER met4 ;
        RECT 192.515 202.730 197.965 341.270 ;
      LAYER met4 ;
        RECT 198.365 202.330 200.000 202.745 ;
        RECT 152.665 198.365 200.000 202.330 ;
        RECT 3385.255 199.600 3389.635 200.000 ;
        POLYGON 3390.035 200.000 3390.035 199.600 3389.635 199.600 ;
        RECT 933.030 198.365 1011.035 199.465 ;
        RECT 1476.030 198.365 1554.035 199.465 ;
        RECT 1750.030 198.365 1828.035 199.465 ;
        RECT 2024.030 198.365 2102.035 199.465 ;
        RECT 2298.030 198.365 2376.035 199.465 ;
        RECT 2572.030 198.365 2650.035 199.465 ;
        RECT 3385.255 198.365 3390.035 199.600 ;
        RECT 152.665 192.115 197.250 198.365 ;
        RECT 197.965 197.965 199.600 198.365 ;
        POLYGON 199.600 198.365 200.000 197.965 199.600 197.965 ;
      LAYER met4 ;
        RECT 197.650 192.515 395.270 197.965 ;
      LAYER met4 ;
        RECT 395.670 192.115 467.330 197.965 ;
      LAYER met4 ;
        RECT 467.730 192.515 664.270 197.965 ;
      LAYER met4 ;
        RECT 664.670 192.115 736.330 197.965 ;
      LAYER met4 ;
        RECT 736.730 192.515 933.270 197.965 ;
      LAYER met4 ;
        RECT 933.670 192.115 1010.330 198.365 ;
      LAYER met4 ;
        RECT 1010.730 192.515 1207.270 197.965 ;
      LAYER met4 ;
        RECT 1207.670 192.115 1279.330 197.965 ;
      LAYER met4 ;
        RECT 1279.730 192.515 1476.270 197.965 ;
      LAYER met4 ;
        RECT 1476.670 192.115 1553.330 198.365 ;
      LAYER met4 ;
        RECT 1553.730 192.515 1750.270 197.965 ;
      LAYER met4 ;
        RECT 1750.670 192.115 1827.330 198.365 ;
      LAYER met4 ;
        RECT 1827.730 192.515 2024.270 197.965 ;
      LAYER met4 ;
        RECT 2024.670 192.115 2101.330 198.365 ;
      LAYER met4 ;
        RECT 2101.730 192.515 2298.270 197.965 ;
      LAYER met4 ;
        RECT 2298.670 192.115 2375.330 198.365 ;
      LAYER met4 ;
        RECT 2375.730 192.515 2572.270 197.965 ;
      LAYER met4 ;
        RECT 2572.670 192.115 2649.330 198.365 ;
        RECT 3385.670 197.965 3390.035 198.365 ;
      LAYER met4 ;
        RECT 2649.730 192.515 2846.270 197.965 ;
      LAYER met4 ;
        RECT 2846.670 192.115 2918.330 197.965 ;
      LAYER met4 ;
        RECT 2918.730 192.515 3115.270 197.965 ;
      LAYER met4 ;
        RECT 3115.670 192.115 3187.330 197.965 ;
      LAYER met4 ;
        RECT 3187.730 192.515 3385.270 197.965 ;
      LAYER met4 ;
        RECT 3385.670 197.250 3389.635 197.965 ;
      LAYER met4 ;
        RECT 3390.035 197.650 3395.485 501.270 ;
      LAYER met4 ;
        RECT 3395.885 501.030 3396.485 501.670 ;
        RECT 3401.935 501.430 3407.385 501.670 ;
        RECT 3395.885 197.250 3396.485 200.000 ;
        RECT 3385.670 195.815 3396.485 197.250 ;
      LAYER met4 ;
        RECT 3396.885 196.215 3401.535 501.270 ;
      LAYER met4 ;
        RECT 3401.935 501.030 3402.535 501.430 ;
        RECT 3406.785 501.030 3407.385 501.430 ;
      LAYER met4 ;
        RECT 3402.935 350.000 3406.385 501.030 ;
      LAYER met4 ;
        RECT 3401.935 198.130 3402.535 200.000 ;
      LAYER met4 ;
        RECT 3402.935 198.530 3406.385 345.000 ;
      LAYER met4 ;
        RECT 3406.785 198.130 3407.385 200.000 ;
      LAYER met4 ;
        RECT 3407.785 198.475 3412.435 501.270 ;
      LAYER met4 ;
        RECT 3412.835 501.030 3413.435 501.670 ;
        RECT 3401.935 198.075 3407.385 198.130 ;
        RECT 3412.835 198.075 3413.435 200.000 ;
      LAYER met4 ;
        RECT 3413.835 198.400 3418.485 501.270 ;
      LAYER met4 ;
        RECT 3418.885 501.030 3419.485 501.670 ;
        RECT 3401.935 198.000 3413.435 198.075 ;
        RECT 3418.885 198.215 3419.485 200.000 ;
      LAYER met4 ;
        RECT 3419.885 198.615 3423.335 501.270 ;
      LAYER met4 ;
        RECT 3423.735 501.030 3424.335 501.670 ;
      LAYER met4 ;
        RECT 3424.735 350.000 3428.185 501.270 ;
      LAYER met4 ;
        RECT 3428.585 501.030 3429.185 501.670 ;
        RECT 3423.735 198.265 3424.335 200.000 ;
      LAYER met4 ;
        RECT 3424.735 198.665 3428.185 345.000 ;
      LAYER met4 ;
        RECT 3428.585 198.265 3429.185 200.000 ;
      LAYER met4 ;
        RECT 3429.585 198.525 3434.235 501.270 ;
      LAYER met4 ;
        RECT 3434.635 501.030 3435.335 501.670 ;
      LAYER met4 ;
        RECT 3435.735 350.000 3436.065 532.910 ;
        RECT 3436.365 527.855 3439.345 751.535 ;
      LAYER met4 ;
        RECT 3439.745 727.670 3440.725 751.935 ;
      LAYER met4 ;
        RECT 3439.645 726.000 3440.825 727.270 ;
      LAYER met4 ;
        RECT 3439.645 580.000 3440.825 726.000 ;
      LAYER met4 ;
        RECT 3439.645 578.730 3440.825 580.000 ;
      LAYER met4 ;
        RECT 3439.745 543.160 3440.725 578.330 ;
      LAYER met4 ;
        RECT 3441.125 543.560 3444.105 767.240 ;
      LAYER met4 ;
        RECT 3444.505 759.310 3588.000 767.640 ;
      LAYER met4 ;
        RECT 3444.405 577.390 3444.735 758.910 ;
      LAYER met4 ;
        RECT 3445.135 727.670 3588.000 759.310 ;
        RECT 3445.135 727.030 3445.835 727.670 ;
        RECT 3445.135 580.000 3445.835 726.000 ;
        RECT 3445.135 578.330 3445.835 579.035 ;
      LAYER met4 ;
        RECT 3446.235 578.730 3450.685 727.270 ;
      LAYER met4 ;
        RECT 3451.085 727.030 3451.685 727.670 ;
        RECT 3451.085 580.000 3451.685 726.000 ;
        RECT 3451.085 578.330 3451.685 579.035 ;
      LAYER met4 ;
        RECT 3452.085 578.730 3456.535 727.270 ;
      LAYER met4 ;
        RECT 3456.935 727.030 3457.635 727.670 ;
        RECT 3456.935 580.000 3457.635 726.000 ;
        RECT 3456.935 578.330 3457.635 579.035 ;
      LAYER met4 ;
        RECT 3458.035 578.730 3483.000 727.270 ;
      LAYER met4 ;
        RECT 3483.400 727.030 3563.385 727.670 ;
      LAYER met4 ;
        RECT 3563.785 726.000 3588.000 727.270 ;
      LAYER met4 ;
        RECT 3483.400 580.000 3588.000 726.000 ;
        RECT 3483.400 578.330 3563.385 579.035 ;
      LAYER met4 ;
        RECT 3563.785 578.730 3588.000 580.000 ;
      LAYER met4 ;
        RECT 3445.135 576.990 3588.000 578.330 ;
        RECT 3444.505 543.160 3588.000 576.990 ;
        RECT 3439.745 541.640 3588.000 543.160 ;
        RECT 3439.745 527.455 3440.725 541.640 ;
        RECT 3436.465 525.935 3440.725 527.455 ;
        RECT 3423.735 198.215 3429.185 198.265 ;
        RECT 3418.885 198.125 3429.185 198.215 ;
        RECT 3434.635 198.125 3435.335 200.000 ;
        RECT 3418.885 198.000 3435.335 198.125 ;
        RECT 3401.935 195.815 3435.335 198.000 ;
        RECT 3385.670 192.115 3435.335 195.815 ;
        RECT 152.665 191.515 200.000 192.115 ;
        RECT 394.965 191.515 468.035 192.115 ;
        RECT 663.965 191.515 737.035 192.115 ;
        RECT 933.030 191.515 1011.035 192.115 ;
        RECT 1206.000 191.515 1280.035 192.115 ;
        RECT 1476.030 191.515 1554.035 192.115 ;
        RECT 1750.030 191.515 1828.035 192.115 ;
        RECT 2024.030 191.515 2102.035 192.115 ;
        RECT 2298.030 191.515 2376.035 192.115 ;
        RECT 2572.030 191.515 2650.035 192.115 ;
        RECT 2845.965 191.515 2919.035 192.115 ;
        RECT 3114.965 191.515 3188.035 192.115 ;
        RECT 3385.255 191.515 3435.335 192.115 ;
        RECT 152.665 186.065 195.815 191.515 ;
      LAYER met4 ;
        RECT 196.215 186.465 395.270 191.115 ;
      LAYER met4 ;
        RECT 395.670 186.065 467.330 191.515 ;
      LAYER met4 ;
        RECT 467.730 186.465 664.270 191.115 ;
      LAYER met4 ;
        RECT 664.670 186.065 736.330 191.515 ;
      LAYER met4 ;
        RECT 736.730 186.465 933.270 191.115 ;
      LAYER met4 ;
        RECT 933.670 186.065 1010.330 191.515 ;
      LAYER met4 ;
        RECT 1010.730 186.465 1207.270 191.115 ;
      LAYER met4 ;
        RECT 1207.670 186.065 1279.330 191.515 ;
      LAYER met4 ;
        RECT 1279.730 186.465 1476.270 191.115 ;
      LAYER met4 ;
        RECT 1476.670 186.065 1553.330 191.515 ;
      LAYER met4 ;
        RECT 1553.730 186.465 1750.270 191.115 ;
      LAYER met4 ;
        RECT 1750.670 186.065 1827.330 191.515 ;
      LAYER met4 ;
        RECT 1827.730 186.465 2024.270 191.115 ;
      LAYER met4 ;
        RECT 2024.670 186.065 2101.330 191.515 ;
      LAYER met4 ;
        RECT 2101.730 186.465 2298.270 191.115 ;
      LAYER met4 ;
        RECT 2298.670 186.065 2375.330 191.515 ;
      LAYER met4 ;
        RECT 2375.730 186.465 2572.270 191.115 ;
      LAYER met4 ;
        RECT 2572.670 186.065 2649.330 191.515 ;
      LAYER met4 ;
        RECT 2649.730 186.465 2846.270 191.115 ;
      LAYER met4 ;
        RECT 2846.670 186.065 2918.330 191.515 ;
      LAYER met4 ;
        RECT 2918.730 186.465 3115.270 191.115 ;
      LAYER met4 ;
        RECT 3115.670 186.065 3187.330 191.515 ;
      LAYER met4 ;
        RECT 3187.730 186.465 3385.270 191.115 ;
      LAYER met4 ;
        RECT 3385.670 186.065 3435.335 191.515 ;
        RECT 152.665 185.465 200.000 186.065 ;
        RECT 394.965 185.465 468.035 186.065 ;
        RECT 663.965 185.465 737.035 186.065 ;
        RECT 933.030 185.465 1011.035 186.065 ;
        RECT 1206.000 185.465 1280.035 186.065 ;
        RECT 1476.030 185.465 1554.035 186.065 ;
        RECT 1750.030 185.465 1828.035 186.065 ;
        RECT 2024.030 185.465 2102.035 186.065 ;
        RECT 2298.030 185.465 2376.035 186.065 ;
        RECT 2572.030 185.465 2650.035 186.065 ;
        RECT 2845.965 185.465 2919.035 186.065 ;
        RECT 3114.965 185.465 3188.035 186.065 ;
        RECT 3385.255 185.465 3435.335 186.065 ;
        RECT 152.665 181.215 198.130 185.465 ;
      LAYER met4 ;
        RECT 198.530 181.615 394.965 185.065 ;
      LAYER met4 ;
        RECT 395.365 181.215 467.635 185.465 ;
        RECT 664.365 181.215 736.635 185.465 ;
      LAYER met4 ;
        RECT 737.035 181.615 933.030 185.065 ;
      LAYER met4 ;
        RECT 933.430 181.215 1010.635 185.465 ;
      LAYER met4 ;
        RECT 1011.035 181.615 1206.965 185.065 ;
      LAYER met4 ;
        RECT 1207.365 181.215 1279.635 185.465 ;
      LAYER met4 ;
        RECT 1280.035 181.615 1476.030 185.065 ;
      LAYER met4 ;
        RECT 1476.430 181.215 1553.635 185.465 ;
      LAYER met4 ;
        RECT 1554.035 181.615 1750.030 185.065 ;
      LAYER met4 ;
        RECT 1750.430 181.215 1827.635 185.465 ;
      LAYER met4 ;
        RECT 1828.035 181.615 2024.030 185.065 ;
      LAYER met4 ;
        RECT 2024.430 181.215 2101.635 185.465 ;
      LAYER met4 ;
        RECT 2102.035 181.615 2298.030 185.065 ;
      LAYER met4 ;
        RECT 2298.430 181.215 2375.635 185.465 ;
      LAYER met4 ;
        RECT 2376.035 181.615 2572.030 185.065 ;
      LAYER met4 ;
        RECT 2572.430 181.215 2649.635 185.465 ;
      LAYER met4 ;
        RECT 2650.035 181.615 2845.965 185.065 ;
      LAYER met4 ;
        RECT 2846.365 181.215 2918.635 185.465 ;
      LAYER met4 ;
        RECT 2919.035 181.615 3114.965 185.065 ;
      LAYER met4 ;
        RECT 3115.365 181.215 3187.635 185.465 ;
      LAYER met4 ;
        RECT 3188.035 181.615 3385.255 185.065 ;
      LAYER met4 ;
        RECT 3385.655 181.215 3435.335 185.465 ;
        RECT 152.665 180.615 200.000 181.215 ;
        RECT 394.965 180.615 468.035 181.215 ;
        RECT 663.965 180.615 737.035 181.215 ;
        RECT 933.030 180.615 1011.035 181.215 ;
        RECT 1206.000 180.615 1280.035 181.215 ;
        RECT 1476.030 180.615 1554.035 181.215 ;
        RECT 1750.030 180.615 1828.035 181.215 ;
        RECT 2024.030 180.615 2102.035 181.215 ;
        RECT 2298.030 180.615 2376.035 181.215 ;
        RECT 2572.030 180.615 2650.035 181.215 ;
        RECT 2845.965 180.615 2919.035 181.215 ;
        RECT 3114.965 180.615 3188.035 181.215 ;
        RECT 3385.255 180.615 3435.335 181.215 ;
        RECT 152.665 180.025 198.075 180.615 ;
        RECT 147.275 176.690 198.075 180.025 ;
        RECT 143.995 176.425 198.075 176.690 ;
        RECT 0.000 175.165 198.075 176.425 ;
      LAYER met4 ;
        RECT 198.475 175.565 395.270 180.215 ;
      LAYER met4 ;
        RECT 395.670 175.165 467.330 180.615 ;
      LAYER met4 ;
        RECT 467.730 175.565 664.270 180.215 ;
      LAYER met4 ;
        RECT 664.670 175.165 736.330 180.615 ;
      LAYER met4 ;
        RECT 736.730 175.565 933.270 180.215 ;
      LAYER met4 ;
        RECT 933.670 175.165 1010.330 180.615 ;
      LAYER met4 ;
        RECT 1010.730 175.565 1207.270 180.215 ;
      LAYER met4 ;
        RECT 1207.670 175.165 1279.330 180.615 ;
      LAYER met4 ;
        RECT 1279.730 175.565 1476.270 180.215 ;
      LAYER met4 ;
        RECT 1476.670 175.165 1553.330 180.615 ;
      LAYER met4 ;
        RECT 1553.730 175.565 1750.270 180.215 ;
      LAYER met4 ;
        RECT 1750.670 175.165 1827.330 180.615 ;
      LAYER met4 ;
        RECT 1827.730 175.565 2024.270 180.215 ;
      LAYER met4 ;
        RECT 2024.670 175.165 2101.330 180.615 ;
      LAYER met4 ;
        RECT 2101.730 175.565 2298.270 180.215 ;
      LAYER met4 ;
        RECT 2298.670 175.165 2375.330 180.615 ;
      LAYER met4 ;
        RECT 2375.730 175.565 2572.270 180.215 ;
      LAYER met4 ;
        RECT 2572.670 175.165 2649.330 180.615 ;
      LAYER met4 ;
        RECT 2649.730 175.565 2846.270 180.215 ;
      LAYER met4 ;
        RECT 2846.670 175.165 2918.330 180.615 ;
      LAYER met4 ;
        RECT 2918.730 175.565 3115.270 180.215 ;
      LAYER met4 ;
        RECT 3115.670 175.165 3187.330 180.615 ;
      LAYER met4 ;
        RECT 3187.730 175.565 3385.270 180.215 ;
      LAYER met4 ;
        RECT 3385.670 180.025 3435.335 180.615 ;
      LAYER met4 ;
        RECT 3435.735 180.425 3436.065 345.000 ;
      LAYER met4 ;
        RECT 3385.670 178.665 3435.965 180.025 ;
      LAYER met4 ;
        RECT 3436.365 179.065 3439.345 525.535 ;
      LAYER met4 ;
        RECT 3439.745 501.670 3440.725 525.935 ;
      LAYER met4 ;
        RECT 3439.645 500.000 3440.825 501.270 ;
      LAYER met4 ;
        RECT 3439.645 350.000 3440.825 500.000 ;
        RECT 3439.645 200.000 3440.825 345.000 ;
        RECT 3385.670 178.050 3439.245 178.665 ;
      LAYER met4 ;
        RECT 3439.645 178.450 3440.825 200.000 ;
      LAYER met4 ;
        RECT 3385.670 176.690 3440.725 178.050 ;
      LAYER met4 ;
        RECT 3441.125 177.090 3444.105 541.240 ;
      LAYER met4 ;
        RECT 3444.505 533.310 3588.000 541.640 ;
      LAYER met4 ;
        RECT 3444.405 350.000 3444.735 532.910 ;
      LAYER met4 ;
        RECT 3445.135 501.670 3588.000 533.310 ;
        RECT 3445.135 501.030 3445.835 501.670 ;
        RECT 3445.135 350.000 3445.835 500.000 ;
      LAYER met4 ;
        RECT 3444.405 176.825 3444.735 345.000 ;
      LAYER met4 ;
        RECT 3445.135 197.975 3445.835 345.000 ;
      LAYER met4 ;
        RECT 3446.235 198.375 3450.685 501.270 ;
      LAYER met4 ;
        RECT 3451.085 501.030 3451.685 501.670 ;
        RECT 3451.085 350.000 3451.685 500.000 ;
        RECT 3451.085 198.120 3451.685 345.000 ;
      LAYER met4 ;
        RECT 3452.085 198.520 3456.535 501.270 ;
      LAYER met4 ;
        RECT 3456.935 501.030 3457.635 501.670 ;
        RECT 3456.935 350.000 3457.635 500.000 ;
        RECT 3456.935 198.120 3457.635 345.000 ;
        RECT 3451.085 197.975 3457.635 198.120 ;
        RECT 3445.135 196.955 3457.635 197.975 ;
      LAYER met4 ;
        RECT 3458.035 197.355 3483.000 501.270 ;
      LAYER met4 ;
        RECT 3483.400 501.030 3563.385 501.670 ;
      LAYER met4 ;
        RECT 3563.785 500.000 3588.000 501.270 ;
      LAYER met4 ;
        RECT 3483.400 350.000 3588.000 500.000 ;
        RECT 3563.785 345.000 3588.000 350.000 ;
        RECT 3483.400 200.000 3588.000 345.000 ;
        RECT 3483.400 198.165 3563.385 200.000 ;
      LAYER met4 ;
        RECT 3563.785 198.565 3588.000 200.000 ;
      LAYER met4 ;
        RECT 3483.400 196.955 3588.000 198.165 ;
        RECT 3385.670 176.425 3444.005 176.690 ;
        RECT 3445.135 176.425 3588.000 196.955 ;
        RECT 3385.670 175.165 3588.000 176.425 ;
        RECT 0.000 174.565 200.000 175.165 ;
        RECT 394.965 174.565 468.035 175.165 ;
        RECT 663.965 174.565 737.035 175.165 ;
        RECT 933.030 174.565 1011.035 175.165 ;
        RECT 1206.000 174.565 1280.035 175.165 ;
        RECT 1476.030 174.565 1554.035 175.165 ;
        RECT 1750.030 174.565 1828.035 175.165 ;
        RECT 2024.030 174.565 2102.035 175.165 ;
        RECT 2298.030 174.565 2376.035 175.165 ;
        RECT 2572.030 174.565 2650.035 175.165 ;
        RECT 2845.965 174.565 2919.035 175.165 ;
        RECT 3114.965 174.565 3188.035 175.165 ;
        RECT 3385.255 174.565 3588.000 175.165 ;
        RECT 0.000 169.115 198.000 174.565 ;
      LAYER met4 ;
        RECT 198.400 169.515 395.270 174.165 ;
      LAYER met4 ;
        RECT 395.670 169.115 467.330 174.565 ;
      LAYER met4 ;
        RECT 467.730 169.515 664.270 174.165 ;
      LAYER met4 ;
        RECT 664.670 169.115 736.330 174.565 ;
      LAYER met4 ;
        RECT 736.730 169.515 933.270 174.165 ;
      LAYER met4 ;
        RECT 933.670 169.115 1010.330 174.565 ;
      LAYER met4 ;
        RECT 1010.730 169.515 1207.270 174.165 ;
      LAYER met4 ;
        RECT 1207.670 169.115 1279.330 174.565 ;
      LAYER met4 ;
        RECT 1279.730 169.515 1476.270 174.165 ;
      LAYER met4 ;
        RECT 1476.670 169.115 1553.330 174.565 ;
      LAYER met4 ;
        RECT 1553.730 169.515 1750.270 174.165 ;
      LAYER met4 ;
        RECT 1750.670 169.115 1827.330 174.565 ;
      LAYER met4 ;
        RECT 1827.730 169.515 2024.270 174.165 ;
      LAYER met4 ;
        RECT 2024.670 169.115 2101.330 174.565 ;
      LAYER met4 ;
        RECT 2101.730 169.515 2298.270 174.165 ;
      LAYER met4 ;
        RECT 2298.670 169.115 2375.330 174.565 ;
      LAYER met4 ;
        RECT 2375.730 169.515 2572.270 174.165 ;
      LAYER met4 ;
        RECT 2572.670 169.115 2649.330 174.565 ;
      LAYER met4 ;
        RECT 2649.730 169.515 2846.270 174.165 ;
      LAYER met4 ;
        RECT 2846.670 169.115 2918.330 174.565 ;
      LAYER met4 ;
        RECT 2918.730 169.515 3115.270 174.165 ;
      LAYER met4 ;
        RECT 3115.670 169.115 3187.330 174.565 ;
      LAYER met4 ;
        RECT 3187.730 169.515 3385.270 174.165 ;
      LAYER met4 ;
        RECT 3385.670 169.115 3588.000 174.565 ;
        RECT 0.000 168.515 200.000 169.115 ;
        RECT 394.965 168.515 468.035 169.115 ;
        RECT 663.965 168.515 737.035 169.115 ;
        RECT 933.030 168.515 1011.035 169.115 ;
        RECT 1206.000 168.515 1280.035 169.115 ;
        RECT 1476.030 168.515 1554.035 169.115 ;
        RECT 1750.030 168.515 1828.035 169.115 ;
        RECT 2024.030 168.515 2102.035 169.115 ;
        RECT 2298.030 168.515 2376.035 169.115 ;
        RECT 2572.030 168.515 2650.035 169.115 ;
        RECT 2845.965 168.515 2919.035 169.115 ;
        RECT 3114.965 168.515 3188.035 169.115 ;
        RECT 3385.255 168.515 3588.000 169.115 ;
        RECT 0.000 164.265 198.215 168.515 ;
      LAYER met4 ;
        RECT 198.615 164.665 395.270 168.115 ;
      LAYER met4 ;
        RECT 395.670 164.265 467.330 168.515 ;
      LAYER met4 ;
        RECT 467.730 164.665 664.270 168.115 ;
      LAYER met4 ;
        RECT 664.670 164.265 736.330 168.515 ;
      LAYER met4 ;
        RECT 736.730 164.665 933.270 168.115 ;
      LAYER met4 ;
        RECT 933.670 164.265 1010.330 168.515 ;
      LAYER met4 ;
        RECT 1010.730 164.665 1207.270 168.115 ;
      LAYER met4 ;
        RECT 1207.670 164.265 1279.330 168.515 ;
      LAYER met4 ;
        RECT 1279.730 164.665 1476.270 168.115 ;
      LAYER met4 ;
        RECT 1476.670 164.265 1553.330 168.515 ;
      LAYER met4 ;
        RECT 1553.730 164.665 1750.270 168.115 ;
      LAYER met4 ;
        RECT 1750.670 164.265 1827.330 168.515 ;
      LAYER met4 ;
        RECT 1827.730 164.665 2024.270 168.115 ;
      LAYER met4 ;
        RECT 2024.670 164.265 2101.330 168.515 ;
      LAYER met4 ;
        RECT 2101.730 164.665 2298.270 168.115 ;
      LAYER met4 ;
        RECT 2298.670 164.265 2375.330 168.515 ;
      LAYER met4 ;
        RECT 2375.730 164.665 2572.270 168.115 ;
      LAYER met4 ;
        RECT 2572.670 164.265 2649.330 168.515 ;
      LAYER met4 ;
        RECT 2649.730 164.665 2846.270 168.115 ;
      LAYER met4 ;
        RECT 2846.670 164.265 2918.330 168.515 ;
      LAYER met4 ;
        RECT 2918.730 164.665 3115.270 168.115 ;
      LAYER met4 ;
        RECT 3115.670 164.265 3187.330 168.515 ;
      LAYER met4 ;
        RECT 3187.730 164.665 3385.270 168.115 ;
      LAYER met4 ;
        RECT 3385.670 164.265 3588.000 168.515 ;
        RECT 0.000 163.665 200.000 164.265 ;
        RECT 394.965 163.665 468.035 164.265 ;
        RECT 663.965 163.665 737.035 164.265 ;
        RECT 933.030 163.665 1011.035 164.265 ;
        RECT 1206.000 163.665 1280.035 164.265 ;
        RECT 1476.030 163.665 1554.035 164.265 ;
        RECT 1750.030 163.665 1828.035 164.265 ;
        RECT 2024.030 163.665 2102.035 164.265 ;
        RECT 2298.030 163.665 2376.035 164.265 ;
        RECT 2572.030 163.665 2650.035 164.265 ;
        RECT 2845.965 163.665 2919.035 164.265 ;
        RECT 3114.965 163.665 3188.035 164.265 ;
        RECT 3385.255 163.665 3588.000 164.265 ;
        RECT 0.000 159.415 198.265 163.665 ;
      LAYER met4 ;
        RECT 198.665 159.815 395.270 163.265 ;
      LAYER met4 ;
        RECT 395.670 159.415 467.330 163.665 ;
      LAYER met4 ;
        RECT 467.730 159.815 664.270 163.265 ;
      LAYER met4 ;
        RECT 664.670 159.415 736.330 163.665 ;
      LAYER met4 ;
        RECT 736.730 159.815 933.270 163.265 ;
      LAYER met4 ;
        RECT 933.670 159.415 1010.330 163.665 ;
      LAYER met4 ;
        RECT 1010.730 159.815 1207.270 163.265 ;
      LAYER met4 ;
        RECT 1207.670 159.415 1279.330 163.665 ;
      LAYER met4 ;
        RECT 1279.730 159.815 1476.270 163.265 ;
      LAYER met4 ;
        RECT 1476.670 159.415 1553.330 163.665 ;
      LAYER met4 ;
        RECT 1553.730 159.815 1750.270 163.265 ;
      LAYER met4 ;
        RECT 1750.670 159.415 1827.330 163.665 ;
      LAYER met4 ;
        RECT 1827.730 159.815 2024.270 163.265 ;
      LAYER met4 ;
        RECT 2024.670 159.415 2101.330 163.665 ;
      LAYER met4 ;
        RECT 2101.730 159.815 2298.270 163.265 ;
      LAYER met4 ;
        RECT 2298.670 159.415 2375.330 163.665 ;
      LAYER met4 ;
        RECT 2375.730 159.815 2572.270 163.265 ;
      LAYER met4 ;
        RECT 2572.670 159.415 2649.330 163.665 ;
      LAYER met4 ;
        RECT 2649.730 159.815 2846.270 163.265 ;
      LAYER met4 ;
        RECT 2846.670 159.415 2918.330 163.665 ;
      LAYER met4 ;
        RECT 2918.730 159.815 3115.270 163.265 ;
      LAYER met4 ;
        RECT 3115.670 159.415 3187.330 163.665 ;
      LAYER met4 ;
        RECT 3187.730 159.815 3385.270 163.265 ;
      LAYER met4 ;
        RECT 3385.670 159.415 3588.000 163.665 ;
        RECT 0.000 158.815 200.000 159.415 ;
        RECT 394.965 158.815 468.035 159.415 ;
        RECT 663.965 158.815 737.035 159.415 ;
        RECT 933.030 158.815 1011.035 159.415 ;
        RECT 1206.000 158.815 1280.035 159.415 ;
        RECT 1476.030 158.815 1554.035 159.415 ;
        RECT 1750.030 158.815 1828.035 159.415 ;
        RECT 2024.030 158.815 2102.035 159.415 ;
        RECT 2298.030 158.815 2376.035 159.415 ;
        RECT 2572.030 158.815 2650.035 159.415 ;
        RECT 2845.965 158.815 2919.035 159.415 ;
        RECT 3114.965 158.815 3188.035 159.415 ;
        RECT 3385.255 158.815 3588.000 159.415 ;
        RECT 0.000 153.365 198.125 158.815 ;
      LAYER met4 ;
        RECT 198.525 153.765 395.270 158.415 ;
      LAYER met4 ;
        RECT 395.670 153.365 467.330 158.815 ;
        RECT 664.670 158.770 736.330 158.815 ;
        RECT 664.745 153.410 736.330 158.770 ;
      LAYER met4 ;
        RECT 736.730 153.765 933.270 158.415 ;
      LAYER met4 ;
        RECT 664.670 153.365 736.330 153.410 ;
        RECT 933.670 153.365 1010.330 158.815 ;
      LAYER met4 ;
        RECT 1010.730 153.765 1207.270 158.415 ;
      LAYER met4 ;
        RECT 1207.670 153.365 1279.330 158.815 ;
      LAYER met4 ;
        RECT 1279.730 153.765 1476.270 158.415 ;
      LAYER met4 ;
        RECT 1476.670 153.365 1553.330 158.815 ;
      LAYER met4 ;
        RECT 1553.730 153.765 1750.270 158.415 ;
      LAYER met4 ;
        RECT 1750.670 153.365 1827.330 158.815 ;
      LAYER met4 ;
        RECT 1827.730 153.765 2024.270 158.415 ;
      LAYER met4 ;
        RECT 2024.670 153.365 2101.330 158.815 ;
      LAYER met4 ;
        RECT 2101.730 153.765 2298.270 158.415 ;
      LAYER met4 ;
        RECT 2298.670 153.365 2375.330 158.815 ;
      LAYER met4 ;
        RECT 2375.730 153.765 2572.270 158.415 ;
      LAYER met4 ;
        RECT 2572.670 153.365 2649.330 158.815 ;
      LAYER met4 ;
        RECT 2649.730 153.765 2846.270 158.415 ;
      LAYER met4 ;
        RECT 2846.670 153.365 2918.330 158.815 ;
      LAYER met4 ;
        RECT 2918.730 153.765 3115.270 158.415 ;
      LAYER met4 ;
        RECT 3115.670 153.365 3187.330 158.815 ;
      LAYER met4 ;
        RECT 3187.730 153.765 3385.270 158.415 ;
      LAYER met4 ;
        RECT 3385.670 153.365 3588.000 158.815 ;
        RECT 0.000 152.665 200.000 153.365 ;
        RECT 394.965 152.665 468.035 153.365 ;
        RECT 663.965 152.665 737.035 153.365 ;
        RECT 933.030 152.665 1011.035 153.365 ;
        RECT 1206.000 152.665 1280.035 153.365 ;
        RECT 1476.030 152.665 1554.035 153.365 ;
        RECT 1750.030 152.665 1828.035 153.365 ;
        RECT 2024.030 152.665 2102.035 153.365 ;
        RECT 2298.030 152.665 2376.035 153.365 ;
        RECT 2572.030 152.665 2650.035 153.365 ;
        RECT 2845.965 152.665 2919.035 153.365 ;
        RECT 3114.965 152.665 3188.035 153.365 ;
        RECT 3385.255 152.665 3588.000 153.365 ;
        RECT 0.000 152.035 180.025 152.665 ;
        RECT 0.000 148.755 178.665 152.035 ;
      LAYER met4 ;
        RECT 180.425 151.935 395.270 152.265 ;
      LAYER met4 ;
        RECT 395.670 152.035 467.330 152.665 ;
      LAYER met4 ;
        RECT 467.730 151.935 964.910 152.265 ;
      LAYER met4 ;
        RECT 965.310 152.035 1008.990 152.665 ;
      LAYER met4 ;
        RECT 1009.390 151.935 1507.910 152.265 ;
      LAYER met4 ;
        RECT 1508.310 152.035 1551.990 152.665 ;
      LAYER met4 ;
        RECT 1552.390 151.935 1781.910 152.265 ;
      LAYER met4 ;
        RECT 1782.310 152.035 1825.990 152.665 ;
      LAYER met4 ;
        RECT 1826.390 151.935 2055.910 152.265 ;
      LAYER met4 ;
        RECT 2056.310 152.035 2099.990 152.665 ;
      LAYER met4 ;
        RECT 2100.390 151.935 2329.910 152.265 ;
      LAYER met4 ;
        RECT 2330.310 152.035 2373.990 152.665 ;
      LAYER met4 ;
        RECT 2374.390 151.935 2603.910 152.265 ;
      LAYER met4 ;
        RECT 2604.310 152.035 2647.990 152.665 ;
      LAYER met4 ;
        RECT 2648.390 151.935 3407.575 152.265 ;
      LAYER met4 ;
        RECT 0.000 147.275 178.050 148.755 ;
      LAYER met4 ;
        RECT 179.065 148.655 957.535 151.635 ;
      LAYER met4 ;
        RECT 0.000 143.995 176.690 147.275 ;
      LAYER met4 ;
        RECT 178.450 147.175 200.000 148.355 ;
      LAYER met4 ;
        RECT 200.000 147.175 394.000 148.355 ;
      LAYER met4 ;
        RECT 394.000 147.175 395.270 148.355 ;
      LAYER met4 ;
        RECT 395.670 147.275 467.330 148.255 ;
      LAYER met4 ;
        RECT 467.730 147.175 469.000 148.355 ;
      LAYER met4 ;
        RECT 469.000 147.175 663.000 148.355 ;
      LAYER met4 ;
        RECT 663.000 147.175 664.270 148.355 ;
      LAYER met4 ;
        RECT 664.670 147.275 736.330 148.255 ;
      LAYER met4 ;
        RECT 736.730 147.175 738.000 148.355 ;
      LAYER met4 ;
        RECT 738.000 147.175 932.000 148.355 ;
      LAYER met4 ;
        RECT 932.000 147.175 933.270 148.355 ;
      LAYER met4 ;
        RECT 957.935 148.255 959.455 151.535 ;
      LAYER met4 ;
        RECT 959.855 148.655 1500.535 151.635 ;
      LAYER met4 ;
        RECT 933.670 147.275 1010.330 148.255 ;
        RECT 0.000 142.865 176.425 143.995 ;
      LAYER met4 ;
        RECT 177.090 143.895 973.240 146.875 ;
        RECT 176.825 143.265 395.270 143.595 ;
      LAYER met4 ;
        RECT 973.640 143.495 975.160 147.275 ;
      LAYER met4 ;
        RECT 1010.730 147.175 1012.000 148.355 ;
      LAYER met4 ;
        RECT 1012.000 147.175 1206.000 148.355 ;
      LAYER met4 ;
        RECT 1206.000 147.175 1207.270 148.355 ;
      LAYER met4 ;
        RECT 1207.670 147.275 1279.330 148.255 ;
      LAYER met4 ;
        RECT 1279.730 147.175 1281.000 148.355 ;
      LAYER met4 ;
        RECT 1281.000 147.175 1475.000 148.355 ;
      LAYER met4 ;
        RECT 1475.000 147.175 1476.270 148.355 ;
      LAYER met4 ;
        RECT 1500.935 148.255 1502.455 151.535 ;
      LAYER met4 ;
        RECT 1502.855 148.655 1774.535 151.635 ;
      LAYER met4 ;
        RECT 1476.670 147.275 1553.330 148.255 ;
      LAYER met4 ;
        RECT 975.560 143.895 1516.240 146.875 ;
      LAYER met4 ;
        RECT 395.670 142.865 467.330 143.495 ;
        RECT 965.310 142.865 1008.990 143.495 ;
      LAYER met4 ;
        RECT 1009.390 143.265 1507.910 143.595 ;
      LAYER met4 ;
        RECT 1516.640 143.495 1518.160 147.275 ;
      LAYER met4 ;
        RECT 1553.730 147.175 1555.000 148.355 ;
      LAYER met4 ;
        RECT 1555.000 147.175 1749.000 148.355 ;
      LAYER met4 ;
        RECT 1749.000 147.175 1750.270 148.355 ;
      LAYER met4 ;
        RECT 1774.935 148.255 1776.455 151.535 ;
      LAYER met4 ;
        RECT 1776.855 148.655 2048.535 151.635 ;
      LAYER met4 ;
        RECT 1750.670 147.275 1827.330 148.255 ;
      LAYER met4 ;
        RECT 1518.560 143.895 1790.240 146.875 ;
      LAYER met4 ;
        RECT 1508.310 142.865 1551.990 143.495 ;
      LAYER met4 ;
        RECT 1552.390 143.265 1781.910 143.595 ;
      LAYER met4 ;
        RECT 1790.640 143.495 1792.160 147.275 ;
      LAYER met4 ;
        RECT 1827.730 147.175 1829.000 148.355 ;
      LAYER met4 ;
        RECT 1829.000 147.175 2023.000 148.355 ;
      LAYER met4 ;
        RECT 2023.000 147.175 2024.270 148.355 ;
      LAYER met4 ;
        RECT 2048.935 148.255 2050.455 151.535 ;
      LAYER met4 ;
        RECT 2050.855 148.655 2322.535 151.635 ;
      LAYER met4 ;
        RECT 2024.670 147.275 2101.330 148.255 ;
      LAYER met4 ;
        RECT 1792.560 143.895 2064.240 146.875 ;
      LAYER met4 ;
        RECT 1782.310 142.865 1825.990 143.495 ;
      LAYER met4 ;
        RECT 1826.390 143.265 2055.910 143.595 ;
      LAYER met4 ;
        RECT 2064.640 143.495 2066.160 147.275 ;
      LAYER met4 ;
        RECT 2101.730 147.175 2103.000 148.355 ;
      LAYER met4 ;
        RECT 2103.000 147.175 2297.000 148.355 ;
      LAYER met4 ;
        RECT 2297.000 147.175 2298.270 148.355 ;
      LAYER met4 ;
        RECT 2322.935 148.255 2324.455 151.535 ;
      LAYER met4 ;
        RECT 2324.855 148.655 2596.535 151.635 ;
      LAYER met4 ;
        RECT 2298.670 147.275 2375.330 148.255 ;
      LAYER met4 ;
        RECT 2066.560 143.895 2338.240 146.875 ;
      LAYER met4 ;
        RECT 2056.310 142.865 2099.990 143.495 ;
      LAYER met4 ;
        RECT 2100.390 143.265 2329.910 143.595 ;
      LAYER met4 ;
        RECT 2338.640 143.495 2340.160 147.275 ;
      LAYER met4 ;
        RECT 2375.730 147.175 2377.000 148.355 ;
      LAYER met4 ;
        RECT 2377.000 147.175 2571.000 148.355 ;
      LAYER met4 ;
        RECT 2571.000 147.175 2572.270 148.355 ;
      LAYER met4 ;
        RECT 2596.935 148.255 2598.455 151.535 ;
      LAYER met4 ;
        RECT 2598.855 148.655 3404.875 151.635 ;
      LAYER met4 ;
        RECT 3407.975 151.535 3588.000 152.665 ;
        RECT 3405.275 148.755 3588.000 151.535 ;
        RECT 2572.670 147.275 2649.330 148.255 ;
      LAYER met4 ;
        RECT 2340.560 143.895 2612.240 146.875 ;
      LAYER met4 ;
        RECT 2330.310 142.865 2373.990 143.495 ;
      LAYER met4 ;
        RECT 2374.390 143.265 2603.910 143.595 ;
      LAYER met4 ;
        RECT 2612.640 143.495 2614.160 147.275 ;
      LAYER met4 ;
        RECT 2649.730 147.175 2651.000 148.355 ;
      LAYER met4 ;
        RECT 2651.000 147.175 2845.000 148.355 ;
      LAYER met4 ;
        RECT 2845.000 147.175 2846.270 148.355 ;
      LAYER met4 ;
        RECT 2846.670 147.275 2918.330 148.255 ;
      LAYER met4 ;
        RECT 2918.730 147.175 2920.000 148.355 ;
      LAYER met4 ;
        RECT 2920.000 147.175 3114.000 148.355 ;
      LAYER met4 ;
        RECT 3114.000 147.175 3115.270 148.355 ;
      LAYER met4 ;
        RECT 3115.670 147.275 3187.330 148.255 ;
      LAYER met4 ;
        RECT 3187.730 147.175 3189.000 148.355 ;
      LAYER met4 ;
        RECT 3189.000 147.175 3384.000 148.355 ;
      LAYER met4 ;
        RECT 3384.000 147.175 3405.555 148.355 ;
      LAYER met4 ;
        RECT 3405.955 147.275 3588.000 148.755 ;
      LAYER met4 ;
        RECT 2614.560 143.895 3410.910 146.875 ;
      LAYER met4 ;
        RECT 3411.310 143.995 3588.000 147.275 ;
        RECT 2604.310 142.865 2647.990 143.495 ;
      LAYER met4 ;
        RECT 2648.390 143.265 3411.175 143.595 ;
      LAYER met4 ;
        RECT 3411.575 142.865 3588.000 143.995 ;
        RECT 0.000 142.165 237.000 142.865 ;
        RECT 357.000 142.165 394.000 142.865 ;
        RECT 394.965 142.165 468.035 142.865 ;
        RECT 469.000 142.165 506.000 142.865 ;
        RECT 626.000 142.165 663.000 142.865 ;
        RECT 663.965 142.165 737.035 142.865 ;
        RECT 738.000 142.165 775.000 142.865 ;
        RECT 895.000 142.165 932.000 142.865 ;
        RECT 933.030 142.165 1011.035 142.865 ;
        RECT 1012.000 142.165 1049.000 142.865 ;
        RECT 1169.000 142.165 1280.035 142.865 ;
        RECT 1281.000 142.165 1318.000 142.865 ;
        RECT 1438.000 142.165 1475.000 142.865 ;
        RECT 1476.030 142.165 1554.035 142.865 ;
        RECT 1555.000 142.165 1592.000 142.865 ;
        RECT 1712.000 142.165 1749.000 142.865 ;
        RECT 1750.030 142.165 1828.035 142.865 ;
        RECT 1829.000 142.165 1866.000 142.865 ;
        RECT 1986.000 142.165 2023.000 142.865 ;
        RECT 2024.030 142.165 2102.035 142.865 ;
        RECT 2103.000 142.165 2140.000 142.865 ;
        RECT 2260.000 142.165 2297.000 142.865 ;
        RECT 2298.030 142.165 2376.035 142.865 ;
        RECT 2377.000 142.165 2414.000 142.865 ;
        RECT 2534.000 142.165 2571.000 142.865 ;
        RECT 2572.030 142.165 2650.035 142.865 ;
        RECT 2651.000 142.165 2688.000 142.865 ;
        RECT 2808.000 142.165 2845.000 142.865 ;
        RECT 2845.965 142.165 2919.035 142.865 ;
        RECT 2920.000 142.165 2957.000 142.865 ;
        RECT 3077.000 142.165 3114.000 142.865 ;
        RECT 3114.965 142.165 3188.035 142.865 ;
        RECT 3189.000 142.165 3226.000 142.865 ;
        RECT 3346.000 142.165 3384.000 142.865 ;
        RECT 3385.255 142.165 3588.000 142.865 ;
        RECT 0.000 136.915 197.975 142.165 ;
      LAYER met4 ;
        RECT 198.375 137.315 395.270 141.765 ;
      LAYER met4 ;
        RECT 395.670 136.915 467.330 142.165 ;
      LAYER met4 ;
        RECT 467.730 137.315 664.270 141.765 ;
      LAYER met4 ;
        RECT 664.670 136.915 736.330 142.165 ;
      LAYER met4 ;
        RECT 736.730 137.315 933.270 141.765 ;
      LAYER met4 ;
        RECT 933.670 136.915 1010.330 142.165 ;
      LAYER met4 ;
        RECT 1010.730 137.315 1207.270 141.765 ;
      LAYER met4 ;
        RECT 1207.670 136.915 1279.330 142.165 ;
      LAYER met4 ;
        RECT 1279.730 137.315 1476.270 141.765 ;
      LAYER met4 ;
        RECT 1476.670 136.915 1553.330 142.165 ;
      LAYER met4 ;
        RECT 1553.730 137.315 1750.270 141.765 ;
      LAYER met4 ;
        RECT 1750.670 136.915 1827.330 142.165 ;
      LAYER met4 ;
        RECT 1827.730 137.315 2024.270 141.765 ;
      LAYER met4 ;
        RECT 2024.670 136.915 2101.330 142.165 ;
      LAYER met4 ;
        RECT 2101.730 137.315 2298.270 141.765 ;
      LAYER met4 ;
        RECT 2298.670 136.915 2375.330 142.165 ;
      LAYER met4 ;
        RECT 2375.730 137.315 2572.270 141.765 ;
      LAYER met4 ;
        RECT 2572.670 136.915 2649.330 142.165 ;
      LAYER met4 ;
        RECT 2649.730 137.315 2846.270 141.765 ;
      LAYER met4 ;
        RECT 2846.670 136.915 2918.330 142.165 ;
      LAYER met4 ;
        RECT 2918.730 137.315 3115.270 141.765 ;
      LAYER met4 ;
        RECT 3115.670 136.915 3187.330 142.165 ;
      LAYER met4 ;
        RECT 3187.730 137.315 3385.270 141.765 ;
      LAYER met4 ;
        RECT 3385.670 136.915 3588.000 142.165 ;
        RECT 0.000 136.315 237.000 136.915 ;
        RECT 357.000 136.315 394.000 136.915 ;
        RECT 394.965 136.315 468.035 136.915 ;
        RECT 469.000 136.315 506.000 136.915 ;
        RECT 626.000 136.315 663.000 136.915 ;
        RECT 663.965 136.315 737.035 136.915 ;
        RECT 738.000 136.315 775.000 136.915 ;
        RECT 895.000 136.315 932.000 136.915 ;
        RECT 933.030 136.315 1011.035 136.915 ;
        RECT 1012.000 136.315 1049.000 136.915 ;
        RECT 1169.000 136.315 1280.035 136.915 ;
        RECT 1281.000 136.315 1318.000 136.915 ;
        RECT 1438.000 136.315 1475.000 136.915 ;
        RECT 1476.030 136.315 1554.035 136.915 ;
        RECT 1555.000 136.315 1592.000 136.915 ;
        RECT 1712.000 136.315 1749.000 136.915 ;
        RECT 1750.030 136.315 1828.035 136.915 ;
        RECT 1829.000 136.315 1866.000 136.915 ;
        RECT 1986.000 136.315 2023.000 136.915 ;
        RECT 2024.030 136.315 2102.035 136.915 ;
        RECT 2103.000 136.315 2140.000 136.915 ;
        RECT 2260.000 136.315 2297.000 136.915 ;
        RECT 2298.030 136.315 2376.035 136.915 ;
        RECT 2377.000 136.315 2414.000 136.915 ;
        RECT 2534.000 136.315 2571.000 136.915 ;
        RECT 2572.030 136.315 2650.035 136.915 ;
        RECT 2651.000 136.315 2688.000 136.915 ;
        RECT 2808.000 136.315 2845.000 136.915 ;
        RECT 2845.965 136.315 2919.035 136.915 ;
        RECT 2920.000 136.315 2957.000 136.915 ;
        RECT 3077.000 136.315 3114.000 136.915 ;
        RECT 3114.965 136.315 3188.035 136.915 ;
        RECT 3189.000 136.315 3226.000 136.915 ;
        RECT 3346.000 136.315 3384.000 136.915 ;
        RECT 3385.255 136.315 3588.000 136.915 ;
        RECT 0.000 131.065 198.120 136.315 ;
      LAYER met4 ;
        RECT 198.520 131.465 395.270 135.915 ;
      LAYER met4 ;
        RECT 395.670 131.065 467.330 136.315 ;
      LAYER met4 ;
        RECT 467.730 131.465 664.270 135.915 ;
      LAYER met4 ;
        RECT 664.670 131.065 736.330 136.315 ;
      LAYER met4 ;
        RECT 736.730 131.465 933.270 135.915 ;
      LAYER met4 ;
        RECT 933.670 131.065 1010.330 136.315 ;
      LAYER met4 ;
        RECT 1010.730 131.465 1207.270 135.915 ;
      LAYER met4 ;
        RECT 1207.670 131.065 1279.330 136.315 ;
      LAYER met4 ;
        RECT 1279.730 131.465 1476.270 135.915 ;
      LAYER met4 ;
        RECT 1476.670 131.065 1553.330 136.315 ;
      LAYER met4 ;
        RECT 1553.730 131.465 1750.270 135.915 ;
      LAYER met4 ;
        RECT 1750.670 131.065 1827.330 136.315 ;
      LAYER met4 ;
        RECT 1827.730 131.465 2024.270 135.915 ;
      LAYER met4 ;
        RECT 2024.670 131.065 2101.330 136.315 ;
      LAYER met4 ;
        RECT 2101.730 131.465 2298.270 135.915 ;
      LAYER met4 ;
        RECT 2298.670 131.065 2375.330 136.315 ;
      LAYER met4 ;
        RECT 2375.730 131.465 2572.270 135.915 ;
      LAYER met4 ;
        RECT 2572.670 131.065 2649.330 136.315 ;
      LAYER met4 ;
        RECT 2649.730 131.465 2846.270 135.915 ;
      LAYER met4 ;
        RECT 2846.670 131.065 2918.330 136.315 ;
      LAYER met4 ;
        RECT 2918.730 131.465 3115.270 135.915 ;
      LAYER met4 ;
        RECT 3115.670 131.065 3187.330 136.315 ;
      LAYER met4 ;
        RECT 3187.730 131.465 3385.270 135.915 ;
      LAYER met4 ;
        RECT 3385.670 131.065 3588.000 136.315 ;
        RECT 0.000 130.365 237.000 131.065 ;
        RECT 357.000 130.365 394.000 131.065 ;
        RECT 394.965 130.365 468.035 131.065 ;
        RECT 469.000 130.365 506.000 131.065 ;
        RECT 626.000 130.365 663.000 131.065 ;
        RECT 663.965 130.365 737.035 131.065 ;
        RECT 738.000 130.365 775.000 131.065 ;
        RECT 895.000 130.365 932.000 131.065 ;
        RECT 933.030 130.365 1011.035 131.065 ;
        RECT 1012.000 130.365 1049.000 131.065 ;
        RECT 1169.000 130.365 1280.035 131.065 ;
        RECT 1281.000 130.365 1318.000 131.065 ;
        RECT 1438.000 130.365 1475.000 131.065 ;
        RECT 1476.030 130.365 1554.035 131.065 ;
        RECT 1555.000 130.365 1592.000 131.065 ;
        RECT 1712.000 130.365 1749.000 131.065 ;
        RECT 1750.030 130.365 1828.035 131.065 ;
        RECT 1829.000 130.365 1866.000 131.065 ;
        RECT 1986.000 130.365 2023.000 131.065 ;
        RECT 2024.030 130.365 2102.035 131.065 ;
        RECT 2103.000 130.365 2140.000 131.065 ;
        RECT 2260.000 130.365 2297.000 131.065 ;
        RECT 2298.030 130.365 2376.035 131.065 ;
        RECT 2377.000 130.365 2414.000 131.065 ;
        RECT 2534.000 130.365 2571.000 131.065 ;
        RECT 2572.030 130.365 2650.035 131.065 ;
        RECT 2651.000 130.365 2688.000 131.065 ;
        RECT 2808.000 130.365 2845.000 131.065 ;
        RECT 2845.965 130.365 2919.035 131.065 ;
        RECT 2920.000 130.365 2957.000 131.065 ;
        RECT 3077.000 130.365 3114.000 131.065 ;
        RECT 3114.965 130.365 3188.035 131.065 ;
        RECT 3189.000 130.365 3226.000 131.065 ;
        RECT 3346.000 130.365 3384.000 131.065 ;
        RECT 3385.255 130.365 3588.000 131.065 ;
        RECT 0.000 104.600 196.955 130.365 ;
      LAYER met4 ;
        RECT 197.355 105.000 395.270 129.965 ;
      LAYER met4 ;
        RECT 395.670 104.600 467.330 130.365 ;
      LAYER met4 ;
        RECT 467.730 105.000 664.270 129.965 ;
      LAYER met4 ;
        RECT 664.670 104.600 736.330 130.365 ;
      LAYER met4 ;
        RECT 736.730 105.000 933.270 129.965 ;
      LAYER met4 ;
        RECT 933.670 104.600 1010.330 130.365 ;
      LAYER met4 ;
        RECT 1010.730 105.000 1207.270 129.965 ;
      LAYER met4 ;
        RECT 1207.670 104.600 1279.330 130.365 ;
      LAYER met4 ;
        RECT 1279.730 105.000 1476.270 129.965 ;
      LAYER met4 ;
        RECT 1476.670 104.600 1553.330 130.365 ;
      LAYER met4 ;
        RECT 1553.730 105.000 1750.270 129.965 ;
      LAYER met4 ;
        RECT 1750.670 104.600 1827.330 130.365 ;
      LAYER met4 ;
        RECT 1827.730 105.000 2024.270 129.965 ;
      LAYER met4 ;
        RECT 2024.670 104.600 2101.330 130.365 ;
      LAYER met4 ;
        RECT 2101.730 105.000 2298.270 129.965 ;
      LAYER met4 ;
        RECT 2298.670 104.600 2375.330 130.365 ;
      LAYER met4 ;
        RECT 2375.730 105.000 2572.270 129.965 ;
      LAYER met4 ;
        RECT 2572.670 104.600 2649.330 130.365 ;
      LAYER met4 ;
        RECT 2649.730 105.000 2846.270 129.965 ;
      LAYER met4 ;
        RECT 2846.670 104.600 2918.330 130.365 ;
      LAYER met4 ;
        RECT 2918.730 105.000 3115.270 129.965 ;
      LAYER met4 ;
        RECT 3115.670 104.600 3187.330 130.365 ;
      LAYER met4 ;
        RECT 3187.730 105.000 3385.855 129.965 ;
      LAYER met4 ;
        RECT 3386.255 104.600 3588.000 130.365 ;
        RECT 0.000 24.615 237.000 104.600 ;
        RECT 0.000 0.000 198.165 24.615 ;
        RECT 200.000 24.215 237.000 24.615 ;
        RECT 357.000 24.215 394.000 104.600 ;
        RECT 394.965 24.615 468.035 104.600 ;
      LAYER met4 ;
        RECT 198.565 0.000 200.000 24.215 ;
      LAYER met4 ;
        RECT 200.000 0.000 394.000 24.215 ;
      LAYER met4 ;
        RECT 394.000 0.000 395.270 24.215 ;
      LAYER met4 ;
        RECT 395.670 0.000 467.330 24.615 ;
        RECT 469.000 24.215 506.000 104.600 ;
        RECT 626.000 24.215 663.000 104.600 ;
        RECT 663.965 24.615 737.035 104.600 ;
      LAYER met4 ;
        RECT 467.730 0.000 469.000 24.215 ;
      LAYER met4 ;
        RECT 469.000 0.000 663.000 24.215 ;
      LAYER met4 ;
        RECT 663.000 0.000 664.270 24.215 ;
      LAYER met4 ;
        RECT 664.670 0.000 736.330 24.615 ;
        RECT 738.000 24.215 775.000 104.600 ;
        RECT 895.000 24.215 932.000 104.600 ;
        RECT 933.030 24.615 1011.035 104.600 ;
      LAYER met4 ;
        RECT 736.730 0.000 738.000 24.215 ;
      LAYER met4 ;
        RECT 738.000 0.000 932.000 24.215 ;
      LAYER met4 ;
        RECT 932.000 0.000 933.270 24.215 ;
      LAYER met4 ;
        RECT 933.670 0.000 1010.330 24.615 ;
        RECT 1012.000 24.215 1049.000 104.600 ;
        RECT 1169.000 24.615 1280.035 104.600 ;
        RECT 1169.000 24.215 1206.000 24.615 ;
      LAYER met4 ;
        RECT 1010.730 0.000 1012.000 24.215 ;
      LAYER met4 ;
        RECT 1012.000 0.000 1206.000 24.215 ;
      LAYER met4 ;
        RECT 1206.000 0.000 1207.270 24.215 ;
      LAYER met4 ;
        RECT 1207.670 0.000 1279.330 24.615 ;
        RECT 1281.000 24.215 1318.000 104.600 ;
        RECT 1438.000 24.215 1475.000 104.600 ;
        RECT 1476.030 24.615 1554.035 104.600 ;
      LAYER met4 ;
        RECT 1279.730 0.000 1281.000 24.215 ;
      LAYER met4 ;
        RECT 1281.000 0.000 1475.000 24.215 ;
      LAYER met4 ;
        RECT 1475.000 0.000 1476.270 24.215 ;
      LAYER met4 ;
        RECT 1476.670 0.000 1553.330 24.615 ;
        RECT 1555.000 24.215 1592.000 104.600 ;
        RECT 1712.000 24.215 1749.000 104.600 ;
        RECT 1750.030 24.615 1828.035 104.600 ;
      LAYER met4 ;
        RECT 1553.730 0.000 1555.000 24.215 ;
      LAYER met4 ;
        RECT 1555.000 0.000 1749.000 24.215 ;
      LAYER met4 ;
        RECT 1749.000 0.000 1750.270 24.215 ;
      LAYER met4 ;
        RECT 1750.670 0.000 1827.330 24.615 ;
        RECT 1829.000 24.215 1866.000 104.600 ;
        RECT 1986.000 24.215 2023.000 104.600 ;
        RECT 2024.030 24.615 2102.035 104.600 ;
      LAYER met4 ;
        RECT 1827.730 0.000 1829.000 24.215 ;
      LAYER met4 ;
        RECT 1829.000 0.000 2023.000 24.215 ;
      LAYER met4 ;
        RECT 2023.000 0.000 2024.270 24.215 ;
      LAYER met4 ;
        RECT 2024.670 0.000 2101.330 24.615 ;
        RECT 2103.000 24.215 2140.000 104.600 ;
        RECT 2260.000 24.215 2297.000 104.600 ;
        RECT 2298.030 24.615 2376.035 104.600 ;
      LAYER met4 ;
        RECT 2101.730 0.000 2103.000 24.215 ;
      LAYER met4 ;
        RECT 2103.000 0.000 2297.000 24.215 ;
      LAYER met4 ;
        RECT 2297.000 0.000 2298.270 24.215 ;
      LAYER met4 ;
        RECT 2298.670 0.000 2375.330 24.615 ;
        RECT 2377.000 24.215 2414.000 104.600 ;
        RECT 2534.000 24.215 2571.000 104.600 ;
        RECT 2572.030 24.615 2650.035 104.600 ;
      LAYER met4 ;
        RECT 2375.730 0.000 2377.000 24.215 ;
      LAYER met4 ;
        RECT 2377.000 0.000 2571.000 24.215 ;
      LAYER met4 ;
        RECT 2571.000 0.000 2572.270 24.215 ;
      LAYER met4 ;
        RECT 2572.670 0.000 2649.330 24.615 ;
        RECT 2651.000 24.215 2688.000 104.600 ;
        RECT 2808.000 24.215 2845.000 104.600 ;
        RECT 2845.965 24.615 2919.035 104.600 ;
      LAYER met4 ;
        RECT 2649.730 0.000 2651.000 24.215 ;
      LAYER met4 ;
        RECT 2651.000 0.000 2845.000 24.215 ;
      LAYER met4 ;
        RECT 2845.000 0.000 2846.270 24.215 ;
      LAYER met4 ;
        RECT 2846.670 0.000 2918.330 24.615 ;
        RECT 2920.000 24.215 2957.000 104.600 ;
        RECT 3077.000 24.215 3114.000 104.600 ;
        RECT 3114.965 24.615 3188.035 104.600 ;
      LAYER met4 ;
        RECT 2918.730 0.000 2920.000 24.215 ;
      LAYER met4 ;
        RECT 2920.000 0.000 3114.000 24.215 ;
      LAYER met4 ;
        RECT 3114.000 0.000 3115.270 24.215 ;
      LAYER met4 ;
        RECT 3115.670 0.000 3187.330 24.615 ;
        RECT 3189.000 24.215 3226.000 104.600 ;
        RECT 3346.000 24.215 3384.000 104.600 ;
        RECT 3385.255 24.615 3588.000 104.600 ;
      LAYER met4 ;
        RECT 3187.730 0.000 3189.000 24.215 ;
      LAYER met4 ;
        RECT 3189.000 0.000 3384.000 24.215 ;
      LAYER met4 ;
        RECT 3384.000 0.000 3385.270 24.215 ;
      LAYER met4 ;
        RECT 3385.670 0.000 3588.000 24.615 ;
      LAYER met5 ;
        RECT 0.000 5084.585 204.000 5188.000 ;
      LAYER met5 ;
        RECT 204.000 5163.785 387.270 5188.000 ;
      LAYER met5 ;
        RECT 388.870 5162.185 458.130 5188.000 ;
      LAYER met5 ;
        RECT 459.730 5163.785 644.270 5188.000 ;
      LAYER met5 ;
        RECT 645.870 5162.185 715.130 5188.000 ;
      LAYER met5 ;
        RECT 716.730 5163.785 901.270 5188.000 ;
      LAYER met5 ;
        RECT 902.870 5162.185 972.130 5188.000 ;
      LAYER met5 ;
        RECT 973.730 5163.785 1105.000 5188.000 ;
      LAYER met5 ;
        RECT 386.000 5155.545 461.000 5162.185 ;
        RECT 386.000 5091.520 391.450 5155.545 ;
        RECT 455.490 5091.520 461.000 5155.545 ;
        RECT 386.000 5084.585 461.000 5091.520 ;
        RECT 643.000 5155.545 718.000 5162.185 ;
        RECT 643.000 5091.520 648.450 5155.545 ;
        RECT 712.490 5091.520 718.000 5155.545 ;
        RECT 643.000 5084.585 718.000 5091.520 ;
        RECT 900.000 5155.545 975.000 5162.185 ;
        RECT 900.000 5091.520 905.450 5155.545 ;
        RECT 969.490 5091.520 975.000 5155.545 ;
        RECT 900.000 5084.585 975.000 5091.520 ;
        RECT 1105.000 5155.545 1274.000 5188.000 ;
      LAYER met5 ;
        RECT 1274.000 5163.785 1368.000 5188.000 ;
      LAYER met5 ;
        RECT 1105.000 5091.520 1157.450 5155.545 ;
        RECT 1221.490 5091.520 1274.000 5155.545 ;
        RECT 1105.000 5084.585 1274.000 5091.520 ;
        RECT 1368.000 5155.545 1537.000 5188.000 ;
      LAYER met5 ;
        RECT 1537.000 5163.785 1667.000 5188.000 ;
      LAYER met5 ;
        RECT 1368.000 5091.520 1420.450 5155.545 ;
        RECT 1484.490 5091.520 1537.000 5155.545 ;
        RECT 1368.000 5084.585 1537.000 5091.520 ;
        RECT 1667.000 5155.545 1742.000 5188.000 ;
      LAYER met5 ;
        RECT 1742.000 5163.785 1877.000 5188.000 ;
      LAYER met5 ;
        RECT 1667.000 5091.520 1672.450 5155.545 ;
        RECT 1736.490 5091.520 1742.000 5155.545 ;
        RECT 1667.000 5084.585 1742.000 5091.520 ;
        RECT 1877.000 5155.545 2046.000 5188.000 ;
      LAYER met5 ;
        RECT 2046.000 5163.785 2370.270 5188.000 ;
      LAYER met5 ;
        RECT 2371.870 5162.185 2441.130 5188.000 ;
      LAYER met5 ;
        RECT 2442.730 5163.785 2627.270 5188.000 ;
      LAYER met5 ;
        RECT 2628.870 5162.185 2698.130 5188.000 ;
      LAYER met5 ;
        RECT 2699.730 5163.785 2878.000 5188.000 ;
      LAYER met5 ;
        RECT 1877.000 5091.520 1929.450 5155.545 ;
        RECT 1993.490 5091.520 2046.000 5155.545 ;
        RECT 1877.000 5084.585 2046.000 5091.520 ;
        RECT 2369.000 5155.545 2444.000 5162.185 ;
        RECT 2369.000 5091.520 2374.450 5155.545 ;
        RECT 2438.490 5091.520 2444.000 5155.545 ;
        RECT 2369.000 5084.585 2444.000 5091.520 ;
        RECT 2626.000 5155.545 2701.000 5162.185 ;
        RECT 2626.000 5091.520 2631.450 5155.545 ;
        RECT 2695.490 5091.520 2701.000 5155.545 ;
        RECT 2626.000 5084.585 2701.000 5091.520 ;
        RECT 2878.000 5155.545 2953.000 5188.000 ;
      LAYER met5 ;
        RECT 2953.000 5163.785 3136.270 5188.000 ;
      LAYER met5 ;
        RECT 3137.870 5162.185 3207.130 5188.000 ;
      LAYER met5 ;
        RECT 3208.730 5163.785 3388.000 5188.000 ;
      LAYER met5 ;
        RECT 2878.000 5091.520 2883.450 5155.545 ;
        RECT 2947.490 5091.520 2953.000 5155.545 ;
        RECT 2878.000 5084.585 2953.000 5091.520 ;
        RECT 3135.000 5155.545 3210.000 5162.185 ;
        RECT 3135.000 5091.520 3140.450 5155.545 ;
        RECT 3204.490 5091.520 3210.000 5155.545 ;
        RECT 3135.000 5084.585 3210.000 5091.520 ;
        RECT 3388.000 5084.585 3588.000 5188.000 ;
        RECT 0.000 5056.435 200.545 5084.585 ;
      LAYER met5 ;
        RECT 202.145 5058.035 387.270 5082.985 ;
      LAYER met5 ;
        RECT 0.000 5046.335 201.130 5056.435 ;
      LAYER met5 ;
        RECT 202.730 5052.185 387.270 5056.435 ;
        RECT 202.730 5046.335 387.270 5050.585 ;
      LAYER met5 ;
        RECT 0.000 5034.135 175.245 5046.335 ;
      LAYER met5 ;
        RECT 176.845 5035.735 387.270 5044.735 ;
      LAYER met5 ;
        RECT 0.000 5012.755 201.130 5034.135 ;
      LAYER met5 ;
        RECT 202.730 5029.685 387.270 5034.135 ;
        RECT 202.730 5024.840 387.270 5028.085 ;
      LAYER met5 ;
        RECT 388.870 5024.840 458.130 5084.585 ;
      LAYER met5 ;
        RECT 459.730 5058.035 644.270 5082.985 ;
        RECT 459.730 5052.185 644.270 5056.435 ;
        RECT 459.730 5046.335 644.270 5050.585 ;
        RECT 459.730 5035.735 644.270 5044.735 ;
        RECT 459.730 5029.685 644.270 5034.135 ;
        RECT 459.730 5024.840 644.270 5028.085 ;
      LAYER met5 ;
        RECT 645.870 5024.840 715.130 5084.585 ;
      LAYER met5 ;
        RECT 716.730 5058.035 901.270 5082.985 ;
        RECT 716.730 5052.185 901.270 5056.435 ;
        RECT 716.730 5046.335 901.270 5050.585 ;
        RECT 716.730 5035.735 901.270 5044.735 ;
        RECT 716.730 5029.685 901.270 5034.135 ;
        RECT 716.730 5024.840 901.270 5028.085 ;
      LAYER met5 ;
        RECT 902.870 5024.840 972.130 5084.585 ;
      LAYER met5 ;
        RECT 973.730 5058.035 1152.715 5082.985 ;
        RECT 973.730 5052.185 1152.715 5056.435 ;
        RECT 973.730 5046.335 1152.715 5050.585 ;
      LAYER met5 ;
        RECT 1154.315 5044.735 1229.285 5084.585 ;
      LAYER met5 ;
        RECT 1230.885 5058.035 1415.715 5082.985 ;
        RECT 1230.885 5052.185 1415.715 5056.435 ;
        RECT 1230.885 5046.335 1415.715 5050.585 ;
      LAYER met5 ;
        RECT 1417.315 5044.735 1492.285 5084.585 ;
      LAYER met5 ;
        RECT 1493.885 5058.035 1668.270 5082.985 ;
        RECT 1493.885 5052.185 1668.270 5056.435 ;
        RECT 1493.885 5046.335 1668.270 5050.585 ;
        RECT 973.730 5035.735 1152.240 5044.735 ;
      LAYER met5 ;
        RECT 1153.840 5035.735 1229.285 5044.735 ;
      LAYER met5 ;
        RECT 1230.885 5035.735 1415.240 5044.735 ;
      LAYER met5 ;
        RECT 1416.840 5035.735 1492.285 5044.735 ;
      LAYER met5 ;
        RECT 1493.885 5035.735 1668.270 5044.735 ;
        RECT 973.730 5029.685 1152.715 5034.135 ;
        RECT 973.730 5024.840 1152.715 5028.085 ;
        RECT 204.000 5024.835 386.000 5024.840 ;
      LAYER met5 ;
        RECT 386.000 5024.835 461.000 5024.840 ;
      LAYER met5 ;
        RECT 461.000 5024.835 643.000 5024.840 ;
      LAYER met5 ;
        RECT 643.000 5024.835 718.000 5024.840 ;
      LAYER met5 ;
        RECT 718.000 5024.835 900.000 5024.840 ;
      LAYER met5 ;
        RECT 900.000 5024.835 975.000 5024.840 ;
      LAYER met5 ;
        RECT 975.000 5024.835 1152.715 5024.840 ;
        RECT 202.730 5019.985 387.270 5023.235 ;
        RECT 202.730 5013.935 387.270 5018.385 ;
      LAYER met5 ;
        RECT 0.000 4992.245 141.665 5012.755 ;
        RECT 0.000 4988.000 103.415 4992.245 ;
        RECT 131.565 4991.225 141.665 4992.245 ;
        RECT 131.565 4991.080 135.815 4991.225 ;
      LAYER met5 ;
        RECT 0.000 4849.730 24.215 4988.000 ;
      LAYER met5 ;
        RECT 25.815 4848.130 103.415 4851.000 ;
      LAYER met5 ;
        RECT 105.015 4849.730 129.965 4990.645 ;
        RECT 131.565 4849.730 135.815 4989.480 ;
        RECT 137.415 4849.730 141.665 4989.625 ;
        RECT 143.265 4849.730 152.265 5011.155 ;
      LAYER met5 ;
        RECT 153.865 5006.285 201.130 5012.755 ;
      LAYER met5 ;
        RECT 202.730 5007.885 387.270 5012.335 ;
      LAYER met5 ;
        RECT 388.870 5006.285 458.130 5024.835 ;
      LAYER met5 ;
        RECT 459.730 5019.985 644.270 5023.235 ;
        RECT 459.730 5013.935 644.270 5018.385 ;
        RECT 459.730 5007.885 644.270 5012.335 ;
      LAYER met5 ;
        RECT 645.870 5006.285 715.130 5024.835 ;
      LAYER met5 ;
        RECT 716.730 5019.985 901.270 5023.235 ;
        RECT 716.730 5013.935 901.270 5018.385 ;
        RECT 716.730 5007.885 901.270 5012.335 ;
      LAYER met5 ;
        RECT 902.870 5006.285 972.130 5024.835 ;
      LAYER met5 ;
        RECT 973.730 5019.985 1152.715 5023.235 ;
        RECT 973.730 5013.935 1152.715 5018.385 ;
        RECT 973.730 5007.885 1152.715 5012.335 ;
      LAYER met5 ;
        RECT 1154.315 5007.885 1229.285 5035.735 ;
      LAYER met5 ;
        RECT 1230.885 5029.685 1415.715 5034.135 ;
        RECT 1230.885 5024.835 1415.715 5028.085 ;
        RECT 1230.885 5019.985 1415.715 5023.235 ;
        RECT 1230.885 5013.935 1415.715 5018.385 ;
        RECT 1230.885 5007.885 1415.715 5012.335 ;
      LAYER met5 ;
        RECT 1417.315 5007.885 1492.285 5035.735 ;
      LAYER met5 ;
        RECT 1493.885 5029.685 1668.270 5034.135 ;
        RECT 1493.885 5024.840 1668.270 5028.085 ;
      LAYER met5 ;
        RECT 1669.870 5024.840 1739.130 5084.585 ;
      LAYER met5 ;
        RECT 1740.730 5058.035 1924.715 5082.985 ;
        RECT 1740.730 5052.185 1924.715 5056.435 ;
        RECT 1740.730 5046.335 1924.715 5050.585 ;
      LAYER met5 ;
        RECT 1926.315 5044.735 2001.285 5084.585 ;
      LAYER met5 ;
        RECT 2002.885 5058.035 2370.270 5082.985 ;
        RECT 2002.885 5052.185 2370.270 5056.435 ;
        RECT 2002.885 5046.335 2370.270 5050.585 ;
        RECT 1740.730 5035.735 1862.000 5044.735 ;
        RECT 1867.000 5035.735 1924.240 5044.735 ;
      LAYER met5 ;
        RECT 1925.840 5035.735 2001.285 5044.735 ;
      LAYER met5 ;
        RECT 2002.885 5035.735 2370.270 5044.735 ;
        RECT 1740.730 5029.685 1924.715 5034.135 ;
        RECT 1740.730 5024.840 1862.000 5028.085 ;
        RECT 1493.885 5024.835 1667.000 5024.840 ;
      LAYER met5 ;
        RECT 1667.000 5024.835 1742.000 5024.840 ;
      LAYER met5 ;
        RECT 1742.000 5024.835 1862.000 5024.840 ;
        RECT 1867.000 5024.835 1924.715 5028.085 ;
        RECT 1493.885 5019.985 1668.270 5023.235 ;
        RECT 1493.885 5013.935 1668.270 5018.385 ;
        RECT 1493.885 5007.885 1668.270 5012.335 ;
      LAYER met5 ;
        RECT 153.865 5003.035 201.145 5006.285 ;
      LAYER met5 ;
        RECT 202.745 5003.035 386.965 5006.285 ;
      LAYER met5 ;
        RECT 388.565 5003.035 458.435 5006.285 ;
      LAYER met5 ;
        RECT 460.035 5003.035 643.965 5006.285 ;
      LAYER met5 ;
        RECT 645.565 5003.035 715.435 5006.285 ;
      LAYER met5 ;
        RECT 717.035 5003.035 900.965 5006.285 ;
      LAYER met5 ;
        RECT 902.565 5003.035 972.435 5006.285 ;
      LAYER met5 ;
        RECT 974.035 5003.035 1152.715 5006.285 ;
      LAYER met5 ;
        RECT 153.865 4993.385 201.130 5003.035 ;
      LAYER met5 ;
        RECT 202.730 4996.985 387.270 5001.435 ;
      LAYER met5 ;
        RECT 153.865 4991.200 184.965 4993.385 ;
        RECT 192.615 4991.950 201.130 4993.385 ;
        RECT 153.865 4991.075 168.015 4991.200 ;
        RECT 175.665 4991.125 184.965 4991.200 ;
        RECT 159.915 4990.985 168.015 4991.075 ;
        RECT 181.715 4991.070 184.965 4991.125 ;
        RECT 159.915 4990.935 163.165 4990.985 ;
      LAYER met5 ;
        RECT 153.865 4849.730 158.315 4989.475 ;
        RECT 159.915 4851.000 163.165 4989.335 ;
        RECT 159.915 4849.730 163.160 4851.000 ;
      LAYER met5 ;
        RECT 163.160 4848.130 163.165 4851.000 ;
      LAYER met5 ;
        RECT 164.765 4849.730 168.015 4989.385 ;
        RECT 169.615 4849.730 174.065 4989.600 ;
        RECT 175.665 4849.730 180.115 4989.525 ;
        RECT 181.715 4850.035 184.965 4989.470 ;
        RECT 186.565 4849.730 191.015 4991.785 ;
        RECT 192.615 4849.730 197.865 4990.350 ;
      LAYER met5 ;
        RECT 199.465 4990.135 201.130 4991.950 ;
      LAYER met5 ;
        RECT 202.730 4990.135 387.270 4995.385 ;
      LAYER met5 ;
        RECT 388.870 4990.135 458.130 5003.035 ;
      LAYER met5 ;
        RECT 459.730 4996.985 644.270 5001.435 ;
        RECT 459.730 4990.135 644.270 4995.385 ;
      LAYER met5 ;
        RECT 645.870 4990.135 715.130 5003.035 ;
      LAYER met5 ;
        RECT 716.730 4996.985 901.270 5001.435 ;
        RECT 716.730 4990.135 901.270 4995.385 ;
      LAYER met5 ;
        RECT 902.870 4990.135 972.130 5003.035 ;
        RECT 1154.315 5001.435 1224.605 5007.885 ;
      LAYER met5 ;
        RECT 1226.205 5003.035 1415.715 5006.285 ;
      LAYER met5 ;
        RECT 1417.315 5001.435 1487.605 5007.885 ;
        RECT 1669.870 5006.285 1739.130 5024.835 ;
      LAYER met5 ;
        RECT 1740.730 5019.985 1924.715 5023.235 ;
        RECT 1740.730 5013.935 1924.715 5018.385 ;
        RECT 1740.730 5007.885 1924.715 5012.335 ;
      LAYER met5 ;
        RECT 1926.315 5007.885 2001.285 5035.735 ;
      LAYER met5 ;
        RECT 2002.885 5029.685 2370.270 5034.135 ;
        RECT 2002.885 5024.840 2370.270 5028.085 ;
      LAYER met5 ;
        RECT 2371.870 5024.840 2441.130 5084.585 ;
      LAYER met5 ;
        RECT 2442.730 5058.035 2627.270 5082.985 ;
        RECT 2442.730 5052.185 2627.270 5056.435 ;
        RECT 2442.730 5046.335 2627.270 5050.585 ;
        RECT 2442.730 5035.735 2627.270 5044.735 ;
        RECT 2442.730 5029.685 2627.270 5034.135 ;
        RECT 2442.730 5024.840 2627.270 5028.085 ;
      LAYER met5 ;
        RECT 2628.870 5024.840 2698.130 5084.585 ;
      LAYER met5 ;
        RECT 2699.730 5058.035 2879.270 5082.985 ;
        RECT 2699.730 5052.185 2879.270 5056.435 ;
        RECT 2699.730 5046.335 2879.270 5050.585 ;
        RECT 2699.730 5035.735 2879.270 5044.735 ;
        RECT 2699.730 5029.685 2879.270 5034.135 ;
        RECT 2699.730 5024.840 2879.270 5028.085 ;
      LAYER met5 ;
        RECT 2880.870 5024.840 2950.130 5084.585 ;
      LAYER met5 ;
        RECT 2951.730 5058.035 3136.270 5082.985 ;
        RECT 2951.730 5052.185 3136.270 5056.435 ;
        RECT 2951.730 5046.335 3136.270 5050.585 ;
        RECT 2951.730 5035.735 3136.270 5044.735 ;
        RECT 2951.730 5029.685 3136.270 5034.135 ;
        RECT 2951.730 5024.840 3136.270 5028.085 ;
      LAYER met5 ;
        RECT 3137.870 5024.840 3207.130 5084.585 ;
      LAYER met5 ;
        RECT 3208.730 5058.035 3390.645 5082.985 ;
      LAYER met5 ;
        RECT 3392.245 5056.435 3588.000 5084.585 ;
      LAYER met5 ;
        RECT 3208.730 5052.185 3389.480 5056.435 ;
      LAYER met5 ;
        RECT 3391.080 5052.185 3588.000 5056.435 ;
      LAYER met5 ;
        RECT 3208.730 5046.335 3389.625 5050.585 ;
      LAYER met5 ;
        RECT 3391.225 5046.335 3588.000 5052.185 ;
      LAYER met5 ;
        RECT 3208.730 5035.735 3411.155 5044.735 ;
      LAYER met5 ;
        RECT 3412.755 5034.135 3588.000 5046.335 ;
      LAYER met5 ;
        RECT 3208.730 5029.685 3389.475 5034.135 ;
      LAYER met5 ;
        RECT 3391.075 5028.085 3588.000 5034.135 ;
      LAYER met5 ;
        RECT 3208.730 5024.840 3389.335 5028.085 ;
        RECT 2002.885 5024.835 2369.000 5024.840 ;
      LAYER met5 ;
        RECT 2369.000 5024.835 2444.000 5024.840 ;
      LAYER met5 ;
        RECT 2444.000 5024.835 2626.000 5024.840 ;
      LAYER met5 ;
        RECT 2626.000 5024.835 2701.000 5024.840 ;
      LAYER met5 ;
        RECT 2701.000 5024.835 2878.000 5024.840 ;
      LAYER met5 ;
        RECT 2878.000 5024.835 2953.000 5024.840 ;
      LAYER met5 ;
        RECT 2953.000 5024.835 3135.000 5024.840 ;
      LAYER met5 ;
        RECT 3135.000 5024.835 3210.000 5024.840 ;
      LAYER met5 ;
        RECT 3210.000 5024.835 3389.335 5024.840 ;
      LAYER met5 ;
        RECT 3390.935 5024.835 3588.000 5028.085 ;
      LAYER met5 ;
        RECT 2002.885 5019.985 2370.270 5023.235 ;
        RECT 2002.885 5013.935 2370.270 5018.385 ;
        RECT 2002.885 5007.885 2370.270 5012.335 ;
        RECT 1489.205 5003.035 1667.965 5006.285 ;
      LAYER met5 ;
        RECT 1669.565 5003.035 1739.435 5006.285 ;
      LAYER met5 ;
        RECT 1741.035 5003.035 1862.000 5006.285 ;
        RECT 1867.000 5003.035 1924.715 5006.285 ;
        RECT 973.730 4996.985 1152.715 5001.435 ;
        RECT 973.730 4990.135 1152.715 4995.385 ;
      LAYER met5 ;
        RECT 1154.315 4990.135 1229.285 5001.435 ;
      LAYER met5 ;
        RECT 1230.885 4996.985 1415.715 5001.435 ;
        RECT 1230.885 4990.135 1415.715 4995.385 ;
      LAYER met5 ;
        RECT 1417.315 4990.135 1492.285 5001.435 ;
      LAYER met5 ;
        RECT 1493.885 4996.985 1668.270 5001.435 ;
        RECT 1493.885 4990.135 1668.270 4995.385 ;
      LAYER met5 ;
        RECT 1669.870 4990.135 1739.130 5003.035 ;
        RECT 1926.315 5001.435 1996.605 5007.885 ;
        RECT 2371.870 5006.285 2441.130 5024.835 ;
      LAYER met5 ;
        RECT 2442.730 5019.985 2627.270 5023.235 ;
        RECT 2442.730 5013.935 2627.270 5018.385 ;
        RECT 2442.730 5007.885 2627.270 5012.335 ;
      LAYER met5 ;
        RECT 2628.870 5006.285 2698.130 5024.835 ;
      LAYER met5 ;
        RECT 2699.730 5019.985 2879.270 5023.235 ;
        RECT 2699.730 5013.935 2879.270 5018.385 ;
        RECT 2699.730 5007.885 2879.270 5012.335 ;
      LAYER met5 ;
        RECT 2880.870 5006.285 2950.130 5024.835 ;
      LAYER met5 ;
        RECT 2951.730 5019.985 3136.270 5023.235 ;
        RECT 2951.730 5013.935 3136.270 5018.385 ;
        RECT 2951.730 5007.885 3136.270 5012.335 ;
      LAYER met5 ;
        RECT 3137.870 5006.285 3207.130 5024.835 ;
      LAYER met5 ;
        RECT 3208.730 5019.985 3389.385 5023.235 ;
      LAYER met5 ;
        RECT 3390.985 5019.985 3588.000 5024.835 ;
      LAYER met5 ;
        RECT 3208.730 5013.935 3389.600 5018.385 ;
      LAYER met5 ;
        RECT 3391.200 5012.755 3588.000 5019.985 ;
        RECT 3391.200 5012.335 3434.135 5012.755 ;
      LAYER met5 ;
        RECT 3208.730 5007.885 3389.525 5012.335 ;
      LAYER met5 ;
        RECT 3391.125 5006.285 3434.135 5012.335 ;
      LAYER met5 ;
        RECT 1998.205 5003.035 2369.965 5006.285 ;
      LAYER met5 ;
        RECT 2371.565 5003.035 2441.435 5006.285 ;
      LAYER met5 ;
        RECT 2443.035 5003.035 2626.965 5006.285 ;
      LAYER met5 ;
        RECT 2628.565 5003.035 2698.435 5006.285 ;
      LAYER met5 ;
        RECT 2700.035 5003.035 2878.965 5006.285 ;
      LAYER met5 ;
        RECT 2880.565 5003.035 2950.435 5006.285 ;
      LAYER met5 ;
        RECT 2952.035 5003.035 3135.965 5006.285 ;
      LAYER met5 ;
        RECT 3137.565 5003.035 3207.435 5006.285 ;
      LAYER met5 ;
        RECT 3209.035 5003.035 3389.470 5006.285 ;
      LAYER met5 ;
        RECT 3391.070 5003.035 3434.135 5006.285 ;
      LAYER met5 ;
        RECT 1740.730 4996.985 1924.715 5001.435 ;
        RECT 1740.730 4990.135 1924.715 4995.385 ;
      LAYER met5 ;
        RECT 1926.315 4990.135 2001.285 5001.435 ;
      LAYER met5 ;
        RECT 2002.885 4996.985 2370.270 5001.435 ;
        RECT 2002.885 4990.135 2370.270 4995.385 ;
      LAYER met5 ;
        RECT 2371.870 4990.135 2441.130 5003.035 ;
      LAYER met5 ;
        RECT 2442.730 4996.985 2627.270 5001.435 ;
        RECT 2442.730 4990.135 2627.270 4995.385 ;
      LAYER met5 ;
        RECT 2628.870 4990.135 2698.130 5003.035 ;
      LAYER met5 ;
        RECT 2699.730 4996.985 2879.270 5001.435 ;
        RECT 2699.730 4990.135 2879.270 4995.385 ;
      LAYER met5 ;
        RECT 2880.870 4990.135 2950.130 5003.035 ;
      LAYER met5 ;
        RECT 2951.730 4996.985 3136.270 5001.435 ;
        RECT 2951.730 4990.135 3136.270 4995.385 ;
      LAYER met5 ;
        RECT 3137.870 4990.135 3207.130 5003.035 ;
      LAYER met5 ;
        RECT 3208.730 4996.985 3391.785 5001.435 ;
      LAYER met5 ;
        RECT 3393.385 4995.385 3434.135 5003.035 ;
      LAYER met5 ;
        RECT 3208.730 4990.135 3390.350 4995.385 ;
      LAYER met5 ;
        RECT 197.865 4989.600 201.130 4990.135 ;
        POLYGON 197.865 4989.600 199.465 4989.600 197.865 4988.000 ;
        RECT 199.465 4988.535 201.130 4989.600 ;
        POLYGON 3388.000 4990.135 3389.600 4990.135 3389.600 4988.535 ;
        RECT 3389.600 4988.535 3390.135 4990.135 ;
        RECT 3391.950 4988.535 3434.135 4995.385 ;
        RECT 199.465 4988.000 204.000 4988.535 ;
        RECT 3388.000 4986.870 3434.135 4988.535 ;
        RECT 3388.000 4984.000 3388.535 4986.870 ;
        RECT 3403.035 4986.855 3406.285 4986.870 ;
        RECT 181.715 4848.130 184.965 4848.435 ;
        RECT 0.000 4845.490 197.865 4848.130 ;
        RECT 0.000 4781.450 32.455 4845.490 ;
        RECT 96.480 4781.450 197.865 4845.490 ;
      LAYER met5 ;
        RECT 3390.135 4831.730 3395.385 4985.270 ;
        RECT 3396.985 4831.730 3401.435 4985.270 ;
        RECT 3403.035 4832.035 3406.285 4985.255 ;
        RECT 3407.885 4831.730 3412.335 4985.270 ;
        RECT 3413.935 4831.730 3418.385 4985.270 ;
        RECT 3419.985 4831.730 3423.235 4985.270 ;
        RECT 3424.840 4984.000 3428.085 4985.270 ;
        RECT 3424.835 4833.000 3428.085 4984.000 ;
      LAYER met5 ;
        RECT 3403.035 4830.130 3406.285 4830.435 ;
        RECT 3424.835 4830.130 3424.840 4833.000 ;
      LAYER met5 ;
        RECT 3424.840 4831.730 3428.085 4833.000 ;
        RECT 3429.685 4831.730 3434.135 4985.270 ;
        RECT 3435.735 4831.730 3444.735 5011.155 ;
      LAYER met5 ;
        RECT 3446.335 4987.455 3588.000 5012.755 ;
        RECT 3446.335 4986.870 3456.435 4987.455 ;
      LAYER met5 ;
        RECT 3446.335 4831.730 3450.585 4985.270 ;
        RECT 3452.185 4831.730 3456.435 4985.270 ;
        RECT 3458.035 4831.730 3482.985 4985.855 ;
      LAYER met5 ;
        RECT 3484.585 4984.000 3588.000 4987.455 ;
        RECT 3484.585 4830.130 3562.185 4833.000 ;
      LAYER met5 ;
        RECT 3563.785 4831.730 3588.000 4984.000 ;
      LAYER met5 ;
        RECT 0.000 4778.870 197.865 4781.450 ;
        RECT 3390.135 4827.550 3588.000 4830.130 ;
      LAYER met5 ;
        RECT 0.000 4635.000 24.215 4777.270 ;
      LAYER met5 ;
        RECT 25.815 4776.000 103.415 4778.870 ;
      LAYER met5 ;
        RECT 105.015 4635.000 129.965 4777.270 ;
        RECT 131.565 4635.000 135.815 4777.270 ;
        RECT 137.415 4635.000 141.665 4777.270 ;
        RECT 143.265 4635.000 152.265 4777.270 ;
        RECT 153.865 4635.000 158.315 4777.270 ;
        RECT 159.915 4776.000 163.160 4777.270 ;
      LAYER met5 ;
        RECT 163.160 4776.000 163.165 4778.870 ;
        RECT 181.715 4778.565 184.965 4778.870 ;
      LAYER met5 ;
        RECT 159.915 4635.000 163.165 4776.000 ;
        RECT 164.765 4635.000 168.015 4777.270 ;
        RECT 169.615 4635.000 174.065 4777.270 ;
        RECT 175.665 4635.000 180.115 4777.270 ;
        RECT 181.715 4635.000 184.965 4776.965 ;
        RECT 186.565 4635.000 191.015 4777.270 ;
        RECT 192.615 4635.000 197.865 4777.270 ;
      LAYER met5 ;
        RECT 3390.135 4763.510 3491.520 4827.550 ;
        RECT 3555.545 4763.510 3588.000 4827.550 ;
        RECT 3390.135 4760.870 3588.000 4763.510 ;
        RECT 3403.035 4760.565 3406.285 4760.870 ;
      LAYER met5 ;
        RECT 3390.135 4613.000 3395.385 4759.270 ;
        RECT 3396.985 4613.000 3401.435 4759.270 ;
        RECT 3403.035 4613.000 3406.285 4758.965 ;
        RECT 3407.885 4613.000 3412.335 4759.270 ;
        RECT 3413.935 4613.000 3418.385 4759.270 ;
        RECT 3419.985 4613.000 3423.235 4759.270 ;
      LAYER met5 ;
        RECT 3424.835 4758.000 3424.840 4760.870 ;
      LAYER met5 ;
        RECT 3424.840 4758.000 3428.085 4759.270 ;
        RECT 3424.835 4613.000 3428.085 4758.000 ;
        RECT 3429.685 4613.000 3434.135 4759.270 ;
        RECT 3435.735 4613.000 3444.735 4759.270 ;
        RECT 3446.335 4613.000 3450.585 4759.270 ;
        RECT 3452.185 4613.000 3456.435 4759.270 ;
        RECT 3458.035 4613.000 3482.985 4759.270 ;
      LAYER met5 ;
        RECT 3484.585 4758.000 3562.185 4760.870 ;
      LAYER met5 ;
        RECT 3563.785 4613.000 3588.000 4759.270 ;
        RECT 0.000 4424.000 24.215 4560.000 ;
      LAYER met5 ;
        RECT 0.000 4421.130 103.415 4424.000 ;
      LAYER met5 ;
        RECT 105.015 4422.730 129.965 4560.000 ;
        RECT 131.565 4422.730 135.815 4560.000 ;
        RECT 137.415 4422.730 141.665 4560.000 ;
        RECT 143.265 4422.730 152.265 4560.000 ;
        RECT 153.865 4422.730 158.315 4560.000 ;
        RECT 159.915 4424.000 163.165 4560.000 ;
        RECT 159.915 4422.730 163.160 4424.000 ;
      LAYER met5 ;
        RECT 163.160 4421.130 163.165 4424.000 ;
      LAYER met5 ;
        RECT 164.765 4422.730 168.015 4560.000 ;
        RECT 169.615 4422.730 174.065 4560.000 ;
        RECT 175.665 4422.730 180.115 4560.000 ;
        RECT 181.715 4423.035 184.965 4560.000 ;
        RECT 186.565 4422.730 191.015 4560.000 ;
        RECT 192.615 4422.730 197.865 4560.000 ;
      LAYER met5 ;
        RECT 181.715 4421.130 184.965 4421.435 ;
        RECT 0.000 4418.490 197.865 4421.130 ;
        RECT 0.000 4354.450 32.455 4418.490 ;
        RECT 96.480 4354.450 197.865 4418.490 ;
      LAYER met5 ;
        RECT 3390.135 4390.730 3395.385 4538.000 ;
        RECT 3396.985 4390.730 3401.435 4538.000 ;
        RECT 3403.035 4391.035 3406.285 4538.000 ;
        RECT 3407.885 4390.730 3412.335 4538.000 ;
        RECT 3413.935 4390.730 3418.385 4538.000 ;
        RECT 3419.985 4390.730 3423.235 4538.000 ;
        RECT 3424.835 4392.000 3428.085 4538.000 ;
        RECT 3424.840 4390.730 3428.085 4392.000 ;
        RECT 3429.685 4390.730 3434.135 4538.000 ;
        RECT 3435.735 4390.730 3444.735 4538.000 ;
        RECT 3446.335 4390.730 3450.585 4538.000 ;
        RECT 3452.185 4390.730 3456.435 4538.000 ;
        RECT 3458.035 4390.730 3482.985 4538.000 ;
        RECT 3563.785 4392.000 3588.000 4538.000 ;
      LAYER met5 ;
        RECT 3403.035 4389.130 3406.285 4389.435 ;
        RECT 3484.585 4389.130 3588.000 4392.000 ;
        RECT 0.000 4351.870 197.865 4354.450 ;
        RECT 3390.135 4382.400 3588.000 4389.130 ;
        RECT 0.000 4349.000 103.415 4351.870 ;
      LAYER met5 ;
        RECT 0.000 4213.000 24.215 4349.000 ;
      LAYER met5 ;
        RECT 0.000 4210.130 103.415 4213.000 ;
      LAYER met5 ;
        RECT 105.015 4211.730 129.965 4350.270 ;
        RECT 131.565 4211.730 135.815 4350.270 ;
        RECT 137.415 4211.730 141.665 4350.270 ;
        RECT 143.265 4211.730 152.265 4350.270 ;
        RECT 153.865 4211.730 158.315 4350.270 ;
        RECT 159.915 4349.000 163.160 4350.270 ;
      LAYER met5 ;
        RECT 163.160 4349.000 163.165 4351.870 ;
        RECT 181.715 4351.565 184.965 4351.870 ;
      LAYER met5 ;
        RECT 159.915 4213.000 163.165 4349.000 ;
        RECT 159.915 4211.730 163.160 4213.000 ;
      LAYER met5 ;
        RECT 163.160 4210.130 163.165 4213.000 ;
      LAYER met5 ;
        RECT 164.765 4211.730 168.015 4350.270 ;
        RECT 169.615 4211.730 174.065 4350.270 ;
        RECT 175.665 4211.730 180.115 4350.270 ;
        RECT 181.715 4212.035 184.965 4349.965 ;
        RECT 186.565 4211.730 191.015 4350.270 ;
        RECT 192.615 4211.730 197.865 4350.270 ;
      LAYER met5 ;
        RECT 3390.135 4316.600 3490.960 4382.400 ;
        RECT 3556.610 4316.600 3588.000 4382.400 ;
        RECT 3390.135 4314.870 3588.000 4316.600 ;
        RECT 3403.035 4314.630 3406.285 4314.870 ;
        RECT 181.715 4210.130 184.965 4210.435 ;
        RECT 0.000 4207.490 197.865 4210.130 ;
        RECT 0.000 4143.450 32.455 4207.490 ;
        RECT 96.480 4143.450 197.865 4207.490 ;
      LAYER met5 ;
        RECT 3390.135 4165.730 3395.385 4313.270 ;
        RECT 3396.985 4165.730 3401.435 4313.270 ;
        RECT 3403.035 4166.035 3406.285 4313.030 ;
        RECT 3407.885 4165.730 3412.335 4313.270 ;
        RECT 3413.935 4165.730 3418.385 4313.270 ;
        RECT 3419.985 4165.730 3423.235 4313.270 ;
        RECT 3424.840 4312.000 3428.085 4313.270 ;
        RECT 3424.835 4167.000 3428.085 4312.000 ;
      LAYER met5 ;
        RECT 3403.035 4164.130 3406.285 4164.435 ;
        RECT 3424.835 4164.130 3424.840 4167.000 ;
      LAYER met5 ;
        RECT 3424.840 4165.730 3428.085 4167.000 ;
        RECT 3429.685 4165.730 3434.135 4313.270 ;
        RECT 3435.735 4165.730 3444.735 4313.270 ;
        RECT 3446.335 4165.730 3450.585 4313.270 ;
        RECT 3452.185 4165.730 3456.435 4313.270 ;
        RECT 3458.035 4165.730 3482.985 4313.270 ;
      LAYER met5 ;
        RECT 3484.585 4312.000 3588.000 4314.870 ;
      LAYER met5 ;
        RECT 3563.785 4167.000 3588.000 4312.000 ;
      LAYER met5 ;
        RECT 3484.585 4164.130 3588.000 4167.000 ;
        RECT 0.000 4140.870 197.865 4143.450 ;
        RECT 3390.135 4161.550 3588.000 4164.130 ;
        RECT 0.000 4138.000 103.415 4140.870 ;
      LAYER met5 ;
        RECT 0.000 4002.000 24.215 4138.000 ;
      LAYER met5 ;
        RECT 0.000 3999.130 103.415 4002.000 ;
      LAYER met5 ;
        RECT 105.015 4000.730 129.965 4139.270 ;
        RECT 131.565 4000.730 135.815 4139.270 ;
        RECT 137.415 4000.730 141.665 4139.270 ;
        RECT 143.265 4000.730 152.265 4139.270 ;
        RECT 153.865 4000.730 158.315 4139.270 ;
        RECT 159.915 4138.000 163.160 4139.270 ;
      LAYER met5 ;
        RECT 163.160 4138.000 163.165 4140.870 ;
        RECT 181.715 4140.565 184.965 4140.870 ;
      LAYER met5 ;
        RECT 159.915 4002.000 163.165 4138.000 ;
        RECT 159.915 4000.730 163.160 4002.000 ;
        RECT 164.765 4000.730 168.015 4139.270 ;
        RECT 169.615 4000.730 174.065 4139.270 ;
        RECT 175.665 4000.730 180.115 4139.270 ;
        RECT 181.715 4000.970 184.965 4138.965 ;
        RECT 186.565 4000.730 191.015 4139.270 ;
        RECT 192.615 4000.730 197.865 4139.270 ;
      LAYER met5 ;
        RECT 3390.135 4097.510 3491.520 4161.550 ;
        RECT 3555.545 4097.510 3588.000 4161.550 ;
        RECT 3390.135 4094.870 3588.000 4097.510 ;
        RECT 3403.035 4094.565 3406.285 4094.870 ;
        RECT 181.715 3999.130 184.965 3999.370 ;
        RECT 0.000 3997.400 197.865 3999.130 ;
        RECT 0.000 3931.600 31.390 3997.400 ;
        RECT 97.040 3931.600 197.865 3997.400 ;
      LAYER met5 ;
        RECT 3390.135 3944.730 3395.385 4093.270 ;
        RECT 3396.985 3944.730 3401.435 4093.270 ;
        RECT 3403.035 3945.035 3406.285 4092.965 ;
        RECT 3407.885 3944.730 3412.335 4093.270 ;
        RECT 3413.935 3944.730 3418.385 4093.270 ;
        RECT 3419.985 3944.730 3423.235 4093.270 ;
      LAYER met5 ;
        RECT 3424.835 4092.000 3424.840 4094.870 ;
      LAYER met5 ;
        RECT 3424.840 4092.000 3428.085 4093.270 ;
        RECT 3424.835 3946.000 3428.085 4092.000 ;
        RECT 3424.840 3944.730 3428.085 3946.000 ;
        RECT 3429.685 3944.730 3434.135 4093.270 ;
        RECT 3435.735 3944.730 3444.735 4093.270 ;
        RECT 3446.335 3944.730 3450.585 4093.270 ;
        RECT 3452.185 3944.730 3456.435 4093.270 ;
        RECT 3458.035 3944.730 3482.985 4093.270 ;
      LAYER met5 ;
        RECT 3484.585 4092.000 3588.000 4094.870 ;
      LAYER met5 ;
        RECT 3563.785 3946.000 3588.000 4092.000 ;
      LAYER met5 ;
        RECT 3403.035 3943.130 3406.285 3943.435 ;
        RECT 3484.585 3943.130 3588.000 3946.000 ;
        RECT 0.000 3924.870 197.865 3931.600 ;
        RECT 3390.135 3936.400 3588.000 3943.130 ;
        RECT 0.000 3922.000 103.415 3924.870 ;
        RECT 181.715 3924.565 184.965 3924.870 ;
      LAYER met5 ;
        RECT 0.000 3786.000 24.215 3922.000 ;
      LAYER met5 ;
        RECT 0.000 3783.130 103.415 3786.000 ;
      LAYER met5 ;
        RECT 105.015 3784.730 129.965 3923.270 ;
        RECT 131.565 3784.730 135.815 3923.270 ;
        RECT 137.415 3784.730 141.665 3923.270 ;
        RECT 143.265 3784.730 152.265 3923.270 ;
        RECT 153.865 3784.730 158.315 3923.270 ;
        RECT 159.915 3922.000 163.160 3923.270 ;
        RECT 159.915 3786.000 163.165 3922.000 ;
        RECT 159.915 3784.730 163.160 3786.000 ;
        RECT 164.765 3784.730 168.015 3923.270 ;
        RECT 169.615 3784.730 174.065 3923.270 ;
        RECT 175.665 3784.730 180.115 3923.270 ;
        RECT 181.715 3784.970 184.965 3922.965 ;
        RECT 186.565 3784.730 191.015 3923.270 ;
        RECT 192.615 3784.730 197.865 3923.270 ;
      LAYER met5 ;
        RECT 3390.135 3870.600 3490.960 3936.400 ;
        RECT 3556.610 3870.600 3588.000 3936.400 ;
        RECT 3390.135 3868.870 3588.000 3870.600 ;
        RECT 3403.035 3868.630 3406.285 3868.870 ;
        RECT 181.715 3783.130 184.965 3783.370 ;
        RECT 0.000 3781.400 197.865 3783.130 ;
        RECT 0.000 3715.600 31.390 3781.400 ;
        RECT 97.040 3715.600 197.865 3781.400 ;
      LAYER met5 ;
        RECT 3390.135 3719.730 3395.385 3867.270 ;
        RECT 3396.985 3719.730 3401.435 3867.270 ;
        RECT 3403.035 3720.035 3406.285 3867.030 ;
        RECT 3407.885 3719.730 3412.335 3867.270 ;
        RECT 3413.935 3719.730 3418.385 3867.270 ;
        RECT 3419.985 3719.730 3423.235 3867.270 ;
        RECT 3424.840 3866.000 3428.085 3867.270 ;
        RECT 3424.835 3721.000 3428.085 3866.000 ;
        RECT 3424.840 3719.730 3428.085 3721.000 ;
        RECT 3429.685 3719.730 3434.135 3867.270 ;
        RECT 3435.735 3719.730 3444.735 3867.270 ;
        RECT 3446.335 3719.730 3450.585 3867.270 ;
        RECT 3452.185 3719.730 3456.435 3867.270 ;
        RECT 3458.035 3719.730 3482.985 3867.270 ;
      LAYER met5 ;
        RECT 3484.585 3866.000 3588.000 3868.870 ;
      LAYER met5 ;
        RECT 3563.785 3721.000 3588.000 3866.000 ;
      LAYER met5 ;
        RECT 3403.035 3718.130 3406.285 3718.435 ;
        RECT 3484.585 3718.130 3588.000 3721.000 ;
        RECT 0.000 3708.870 197.865 3715.600 ;
        RECT 3390.135 3711.400 3588.000 3718.130 ;
        RECT 0.000 3706.000 103.415 3708.870 ;
        RECT 181.715 3708.565 184.965 3708.870 ;
      LAYER met5 ;
        RECT 0.000 3570.000 24.215 3706.000 ;
      LAYER met5 ;
        RECT 0.000 3567.130 103.415 3570.000 ;
      LAYER met5 ;
        RECT 105.015 3568.730 129.965 3707.270 ;
        RECT 131.565 3568.730 135.815 3707.270 ;
        RECT 137.415 3568.730 141.665 3707.270 ;
        RECT 143.265 3568.730 152.265 3707.270 ;
        RECT 153.865 3568.730 158.315 3707.270 ;
        RECT 159.915 3706.000 163.160 3707.270 ;
        RECT 159.915 3570.000 163.165 3706.000 ;
        RECT 159.915 3568.730 163.160 3570.000 ;
        RECT 164.765 3568.730 168.015 3707.270 ;
        RECT 169.615 3568.730 174.065 3707.270 ;
        RECT 175.665 3568.730 180.115 3707.270 ;
        RECT 181.715 3568.970 184.965 3706.965 ;
        RECT 186.565 3568.730 191.015 3707.270 ;
        RECT 192.615 3568.730 197.865 3707.270 ;
      LAYER met5 ;
        RECT 3390.135 3645.600 3490.960 3711.400 ;
        RECT 3556.610 3645.600 3588.000 3711.400 ;
        RECT 3390.135 3643.870 3588.000 3645.600 ;
        RECT 3403.035 3643.630 3406.285 3643.870 ;
        RECT 181.715 3567.130 184.965 3567.370 ;
        RECT 0.000 3565.400 197.865 3567.130 ;
        RECT 0.000 3499.600 31.390 3565.400 ;
        RECT 97.040 3499.600 197.865 3565.400 ;
        RECT 0.000 3492.870 197.865 3499.600 ;
      LAYER met5 ;
        RECT 3390.135 3494.730 3395.385 3642.270 ;
        RECT 3396.985 3494.730 3401.435 3642.270 ;
        RECT 3403.035 3495.035 3406.285 3642.030 ;
        RECT 3407.885 3494.730 3412.335 3642.270 ;
        RECT 3413.935 3494.730 3418.385 3642.270 ;
        RECT 3419.985 3494.730 3423.235 3642.270 ;
        RECT 3424.840 3641.000 3428.085 3642.270 ;
        RECT 3424.835 3496.000 3428.085 3641.000 ;
        RECT 3424.840 3494.730 3428.085 3496.000 ;
        RECT 3429.685 3494.730 3434.135 3642.270 ;
        RECT 3435.735 3494.730 3444.735 3642.270 ;
        RECT 3446.335 3494.730 3450.585 3642.270 ;
        RECT 3452.185 3494.730 3456.435 3642.270 ;
        RECT 3458.035 3494.730 3482.985 3642.270 ;
      LAYER met5 ;
        RECT 3484.585 3641.000 3588.000 3643.870 ;
      LAYER met5 ;
        RECT 3563.785 3496.000 3588.000 3641.000 ;
      LAYER met5 ;
        RECT 3403.035 3493.130 3406.285 3493.435 ;
        RECT 3484.585 3493.130 3588.000 3496.000 ;
        RECT 0.000 3490.000 103.415 3492.870 ;
        RECT 181.715 3492.565 184.965 3492.870 ;
      LAYER met5 ;
        RECT 0.000 3354.000 24.215 3490.000 ;
      LAYER met5 ;
        RECT 0.000 3351.130 103.415 3354.000 ;
      LAYER met5 ;
        RECT 105.015 3352.730 129.965 3491.270 ;
        RECT 131.565 3352.730 135.815 3491.270 ;
        RECT 137.415 3352.730 141.665 3491.270 ;
        RECT 143.265 3352.730 152.265 3491.270 ;
        RECT 153.865 3352.730 158.315 3491.270 ;
        RECT 159.915 3490.000 163.160 3491.270 ;
        RECT 159.915 3354.000 163.165 3490.000 ;
        RECT 159.915 3352.730 163.160 3354.000 ;
        RECT 164.765 3352.730 168.015 3491.270 ;
        RECT 169.615 3352.730 174.065 3491.270 ;
        RECT 175.665 3352.730 180.115 3491.270 ;
        RECT 181.715 3352.970 184.965 3490.965 ;
        RECT 186.565 3352.730 191.015 3491.270 ;
        RECT 192.615 3352.730 197.865 3491.270 ;
      LAYER met5 ;
        RECT 3390.135 3486.400 3588.000 3493.130 ;
        RECT 3390.135 3420.600 3490.960 3486.400 ;
        RECT 3556.610 3420.600 3588.000 3486.400 ;
        RECT 3390.135 3418.870 3588.000 3420.600 ;
        RECT 3403.035 3418.630 3406.285 3418.870 ;
        RECT 181.715 3351.130 184.965 3351.370 ;
        RECT 0.000 3349.400 197.865 3351.130 ;
        RECT 0.000 3283.600 31.390 3349.400 ;
        RECT 97.040 3283.600 197.865 3349.400 ;
        RECT 0.000 3276.870 197.865 3283.600 ;
        RECT 0.000 3274.000 103.415 3276.870 ;
        RECT 181.715 3276.565 184.965 3276.870 ;
      LAYER met5 ;
        RECT 0.000 3138.000 24.215 3274.000 ;
      LAYER met5 ;
        RECT 0.000 3135.130 103.415 3138.000 ;
      LAYER met5 ;
        RECT 105.015 3136.730 129.965 3275.270 ;
        RECT 131.565 3136.730 135.815 3275.270 ;
        RECT 137.415 3136.730 141.665 3275.270 ;
        RECT 143.265 3136.730 152.265 3275.270 ;
        RECT 153.865 3136.730 158.315 3275.270 ;
        RECT 159.915 3274.000 163.160 3275.270 ;
        RECT 159.915 3138.000 163.165 3274.000 ;
        RECT 159.915 3136.730 163.160 3138.000 ;
        RECT 164.765 3136.730 168.015 3275.270 ;
        RECT 169.615 3136.730 174.065 3275.270 ;
        RECT 175.665 3136.730 180.115 3275.270 ;
        RECT 181.715 3136.970 184.965 3274.965 ;
        RECT 186.565 3136.730 191.015 3275.270 ;
        RECT 192.615 3136.730 197.865 3275.270 ;
        RECT 3390.135 3268.730 3395.385 3417.270 ;
        RECT 3396.985 3268.730 3401.435 3417.270 ;
        RECT 3403.035 3269.035 3406.285 3417.030 ;
        RECT 3407.885 3268.730 3412.335 3417.270 ;
        RECT 3413.935 3268.730 3418.385 3417.270 ;
        RECT 3419.985 3268.730 3423.235 3417.270 ;
        RECT 3424.840 3416.000 3428.085 3417.270 ;
        RECT 3424.835 3270.000 3428.085 3416.000 ;
        RECT 3424.840 3268.730 3428.085 3270.000 ;
        RECT 3429.685 3268.730 3434.135 3417.270 ;
        RECT 3435.735 3268.730 3444.735 3417.270 ;
        RECT 3446.335 3268.730 3450.585 3417.270 ;
        RECT 3452.185 3268.730 3456.435 3417.270 ;
        RECT 3458.035 3268.730 3482.985 3417.270 ;
      LAYER met5 ;
        RECT 3484.585 3416.000 3588.000 3418.870 ;
      LAYER met5 ;
        RECT 3563.785 3270.000 3588.000 3416.000 ;
      LAYER met5 ;
        RECT 3403.035 3267.130 3406.285 3267.435 ;
        RECT 3484.585 3267.130 3588.000 3270.000 ;
        RECT 3390.135 3260.400 3588.000 3267.130 ;
        RECT 3390.135 3194.600 3490.960 3260.400 ;
        RECT 3556.610 3194.600 3588.000 3260.400 ;
        RECT 3390.135 3192.870 3588.000 3194.600 ;
        RECT 3403.035 3192.630 3406.285 3192.870 ;
        RECT 181.715 3135.130 184.965 3135.370 ;
        RECT 0.000 3133.400 197.865 3135.130 ;
        RECT 0.000 3067.600 31.390 3133.400 ;
        RECT 97.040 3067.600 197.865 3133.400 ;
        RECT 0.000 3060.870 197.865 3067.600 ;
        RECT 0.000 3058.000 103.415 3060.870 ;
        RECT 181.715 3060.565 184.965 3060.870 ;
      LAYER met5 ;
        RECT 0.000 2922.000 24.215 3058.000 ;
      LAYER met5 ;
        RECT 0.000 2919.130 103.415 2922.000 ;
      LAYER met5 ;
        RECT 105.015 2920.730 129.965 3059.270 ;
        RECT 131.565 2920.730 135.815 3059.270 ;
        RECT 137.415 2920.730 141.665 3059.270 ;
        RECT 143.265 2920.730 152.265 3059.270 ;
        RECT 153.865 2920.730 158.315 3059.270 ;
        RECT 159.915 3058.000 163.160 3059.270 ;
        RECT 159.915 2922.000 163.165 3058.000 ;
        RECT 159.915 2920.730 163.160 2922.000 ;
        RECT 164.765 2920.730 168.015 3059.270 ;
        RECT 169.615 2920.730 174.065 3059.270 ;
        RECT 175.665 2920.730 180.115 3059.270 ;
        RECT 181.715 2920.970 184.965 3058.965 ;
        RECT 186.565 2920.730 191.015 3059.270 ;
        RECT 192.615 2920.730 197.865 3059.270 ;
        RECT 3390.135 3043.730 3395.385 3191.270 ;
        RECT 3396.985 3043.730 3401.435 3191.270 ;
        RECT 3403.035 3044.035 3406.285 3191.030 ;
        RECT 3407.885 3043.730 3412.335 3191.270 ;
        RECT 3413.935 3043.730 3418.385 3191.270 ;
        RECT 3419.985 3043.730 3423.235 3191.270 ;
        RECT 3424.840 3190.000 3428.085 3191.270 ;
        RECT 3424.835 3045.000 3428.085 3190.000 ;
        RECT 3424.840 3043.730 3428.085 3045.000 ;
        RECT 3429.685 3043.730 3434.135 3191.270 ;
        RECT 3435.735 3043.730 3444.735 3191.270 ;
        RECT 3446.335 3043.730 3450.585 3191.270 ;
        RECT 3452.185 3043.730 3456.435 3191.270 ;
        RECT 3458.035 3043.730 3482.985 3191.270 ;
      LAYER met5 ;
        RECT 3484.585 3190.000 3588.000 3192.870 ;
      LAYER met5 ;
        RECT 3563.785 3045.000 3588.000 3190.000 ;
      LAYER met5 ;
        RECT 3403.035 3042.130 3406.285 3042.435 ;
        RECT 3484.585 3042.130 3588.000 3045.000 ;
        RECT 3390.135 3035.400 3588.000 3042.130 ;
        RECT 3390.135 2969.600 3490.960 3035.400 ;
        RECT 3556.610 2969.600 3588.000 3035.400 ;
        RECT 3390.135 2967.870 3588.000 2969.600 ;
        RECT 3403.035 2967.630 3406.285 2967.870 ;
        RECT 181.715 2919.130 184.965 2919.370 ;
        RECT 0.000 2917.400 197.865 2919.130 ;
        RECT 0.000 2851.600 31.390 2917.400 ;
        RECT 97.040 2851.600 197.865 2917.400 ;
        RECT 0.000 2844.870 197.865 2851.600 ;
        RECT 0.000 2842.000 103.415 2844.870 ;
        RECT 181.715 2844.565 184.965 2844.870 ;
      LAYER met5 ;
        RECT 0.000 2706.000 24.215 2842.000 ;
      LAYER met5 ;
        RECT 0.000 2703.130 103.415 2706.000 ;
      LAYER met5 ;
        RECT 105.015 2704.730 129.965 2843.270 ;
        RECT 131.565 2704.730 135.815 2843.270 ;
        RECT 137.415 2704.730 141.665 2843.270 ;
        RECT 143.265 2704.730 152.265 2843.270 ;
        RECT 153.865 2704.730 158.315 2843.270 ;
        RECT 159.915 2842.000 163.160 2843.270 ;
        RECT 159.915 2706.000 163.165 2842.000 ;
        RECT 159.915 2704.730 163.160 2706.000 ;
        RECT 164.765 2704.730 168.015 2843.270 ;
        RECT 169.615 2704.730 174.065 2843.270 ;
        RECT 175.665 2704.730 180.115 2843.270 ;
        RECT 181.715 2704.970 184.965 2842.965 ;
        RECT 186.565 2704.730 191.015 2843.270 ;
        RECT 192.615 2704.730 197.865 2843.270 ;
        RECT 3390.135 2817.730 3395.385 2966.270 ;
        RECT 3396.985 2817.730 3401.435 2966.270 ;
        RECT 3403.035 2818.035 3406.285 2966.030 ;
        RECT 3407.885 2817.730 3412.335 2966.270 ;
        RECT 3413.935 2817.730 3418.385 2966.270 ;
        RECT 3419.985 2817.730 3423.235 2966.270 ;
        RECT 3424.840 2965.000 3428.085 2966.270 ;
        RECT 3424.835 2819.000 3428.085 2965.000 ;
        RECT 3424.840 2817.730 3428.085 2819.000 ;
        RECT 3429.685 2817.730 3434.135 2966.270 ;
        RECT 3435.735 2817.730 3444.735 2966.270 ;
        RECT 3446.335 2817.730 3450.585 2966.270 ;
        RECT 3452.185 2817.730 3456.435 2966.270 ;
        RECT 3458.035 2817.730 3482.985 2966.270 ;
      LAYER met5 ;
        RECT 3484.585 2965.000 3588.000 2967.870 ;
      LAYER met5 ;
        RECT 3563.785 2819.000 3588.000 2965.000 ;
      LAYER met5 ;
        RECT 3403.035 2816.130 3406.285 2816.435 ;
        RECT 3484.585 2816.130 3588.000 2819.000 ;
        RECT 3390.135 2809.400 3588.000 2816.130 ;
        RECT 3390.135 2743.600 3490.960 2809.400 ;
        RECT 3556.610 2743.600 3588.000 2809.400 ;
        RECT 3390.135 2741.870 3588.000 2743.600 ;
        RECT 3403.035 2741.630 3406.285 2741.870 ;
        RECT 181.715 2703.130 184.965 2703.370 ;
        RECT 0.000 2701.400 197.865 2703.130 ;
        RECT 0.000 2635.600 31.390 2701.400 ;
        RECT 97.040 2635.600 197.865 2701.400 ;
        RECT 0.000 2628.870 197.865 2635.600 ;
        RECT 0.000 2626.000 103.415 2628.870 ;
        RECT 181.715 2628.565 184.965 2628.870 ;
      LAYER met5 ;
        RECT 0.000 2490.000 24.215 2626.000 ;
      LAYER met5 ;
        RECT 0.000 2487.130 103.415 2490.000 ;
      LAYER met5 ;
        RECT 105.015 2488.730 129.965 2627.270 ;
        RECT 131.565 2488.730 135.815 2627.270 ;
        RECT 137.415 2488.730 141.665 2627.270 ;
        RECT 143.265 2488.730 152.265 2627.270 ;
        RECT 153.865 2488.730 158.315 2627.270 ;
        RECT 159.915 2626.000 163.160 2627.270 ;
        RECT 159.915 2490.000 163.165 2626.000 ;
        RECT 159.915 2488.730 163.160 2490.000 ;
      LAYER met5 ;
        RECT 163.160 2487.130 163.165 2490.000 ;
      LAYER met5 ;
        RECT 164.765 2488.730 168.015 2627.270 ;
        RECT 169.615 2488.730 174.065 2627.270 ;
        RECT 175.665 2488.730 180.115 2627.270 ;
        RECT 181.715 2489.035 184.965 2626.965 ;
        RECT 186.565 2488.730 191.015 2627.270 ;
        RECT 192.615 2488.730 197.865 2627.270 ;
        RECT 3390.135 2592.730 3395.385 2740.270 ;
        RECT 3396.985 2592.730 3401.435 2740.270 ;
        RECT 3403.035 2593.035 3406.285 2740.030 ;
        RECT 3407.885 2592.730 3412.335 2740.270 ;
        RECT 3413.935 2592.730 3418.385 2740.270 ;
        RECT 3419.985 2592.730 3423.235 2740.270 ;
        RECT 3424.840 2739.000 3428.085 2740.270 ;
        RECT 3424.835 2594.000 3428.085 2739.000 ;
      LAYER met5 ;
        RECT 3403.035 2591.130 3406.285 2591.435 ;
        RECT 3424.835 2591.130 3424.840 2594.000 ;
      LAYER met5 ;
        RECT 3424.840 2592.730 3428.085 2594.000 ;
        RECT 3429.685 2592.730 3434.135 2740.270 ;
        RECT 3435.735 2592.730 3444.735 2740.270 ;
        RECT 3446.335 2592.730 3450.585 2740.270 ;
        RECT 3452.185 2592.730 3456.435 2740.270 ;
        RECT 3458.035 2592.730 3482.985 2740.270 ;
      LAYER met5 ;
        RECT 3484.585 2739.000 3588.000 2741.870 ;
      LAYER met5 ;
        RECT 3563.785 2594.000 3588.000 2739.000 ;
      LAYER met5 ;
        RECT 3484.585 2591.130 3588.000 2594.000 ;
        RECT 3390.135 2588.550 3588.000 2591.130 ;
        RECT 3390.135 2524.510 3491.520 2588.550 ;
        RECT 3555.545 2524.510 3588.000 2588.550 ;
        RECT 3390.135 2521.870 3588.000 2524.510 ;
        RECT 3403.035 2521.565 3406.285 2521.870 ;
        RECT 181.715 2487.130 184.965 2487.435 ;
        RECT 0.000 2484.490 197.865 2487.130 ;
        RECT 0.000 2420.450 32.455 2484.490 ;
        RECT 96.480 2420.450 197.865 2484.490 ;
        RECT 0.000 2417.870 197.865 2420.450 ;
        RECT 0.000 2415.000 103.415 2417.870 ;
      LAYER met5 ;
        RECT 0.000 2279.000 24.215 2415.000 ;
        RECT 105.015 2279.000 129.965 2416.270 ;
        RECT 131.565 2279.000 135.815 2416.270 ;
        RECT 137.415 2279.000 141.665 2416.270 ;
        RECT 143.265 2279.000 152.265 2416.270 ;
        RECT 153.865 2279.000 158.315 2416.270 ;
        RECT 159.915 2415.000 163.160 2416.270 ;
      LAYER met5 ;
        RECT 163.160 2415.000 163.165 2417.870 ;
        RECT 181.715 2417.565 184.965 2417.870 ;
      LAYER met5 ;
        RECT 159.915 2279.000 163.165 2415.000 ;
        RECT 164.765 2279.000 168.015 2416.270 ;
        RECT 169.615 2279.000 174.065 2416.270 ;
        RECT 175.665 2279.000 180.115 2416.270 ;
        RECT 181.715 2279.000 184.965 2415.965 ;
        RECT 186.565 2279.000 191.015 2416.270 ;
        RECT 192.615 2279.000 197.865 2416.270 ;
        RECT 3390.135 2374.000 3395.385 2520.270 ;
        RECT 3396.985 2374.000 3401.435 2520.270 ;
        RECT 3403.035 2374.000 3406.285 2519.965 ;
        RECT 3407.885 2374.000 3412.335 2520.270 ;
        RECT 3413.935 2374.000 3418.385 2520.270 ;
        RECT 3419.985 2374.000 3423.235 2520.270 ;
      LAYER met5 ;
        RECT 3424.835 2519.000 3424.840 2521.870 ;
      LAYER met5 ;
        RECT 3424.840 2519.000 3428.085 2520.270 ;
        RECT 3424.835 2374.000 3428.085 2519.000 ;
        RECT 3429.685 2374.000 3434.135 2520.270 ;
        RECT 3435.735 2374.000 3444.735 2520.270 ;
        RECT 3446.335 2374.000 3450.585 2520.270 ;
        RECT 3452.185 2374.000 3456.435 2520.270 ;
        RECT 3458.035 2374.000 3482.985 2520.270 ;
      LAYER met5 ;
        RECT 3484.585 2519.000 3588.000 2521.870 ;
      LAYER met5 ;
        RECT 3563.785 2374.000 3588.000 2519.000 ;
        RECT 0.000 2068.000 24.215 2204.000 ;
      LAYER met5 ;
        RECT 0.000 2065.130 103.415 2068.000 ;
      LAYER met5 ;
        RECT 105.015 2066.730 129.965 2204.000 ;
        RECT 131.565 2066.730 135.815 2204.000 ;
        RECT 137.415 2066.730 141.665 2204.000 ;
        RECT 143.265 2066.730 152.265 2204.000 ;
        RECT 153.865 2066.730 158.315 2204.000 ;
        RECT 159.915 2068.000 163.165 2204.000 ;
        RECT 159.915 2066.730 163.160 2068.000 ;
        RECT 164.765 2066.730 168.015 2204.000 ;
        RECT 169.615 2066.730 174.065 2204.000 ;
        RECT 175.665 2066.730 180.115 2204.000 ;
        RECT 181.715 2066.970 184.965 2204.000 ;
        RECT 186.565 2066.730 191.015 2204.000 ;
        RECT 192.615 2066.730 197.865 2204.000 ;
        RECT 3390.135 2151.730 3395.385 2299.000 ;
        RECT 3396.985 2151.730 3401.435 2299.000 ;
        RECT 3403.035 2152.035 3406.285 2299.000 ;
        RECT 3407.885 2151.730 3412.335 2299.000 ;
        RECT 3413.935 2151.730 3418.385 2299.000 ;
        RECT 3419.985 2151.730 3423.235 2299.000 ;
        RECT 3424.835 2153.000 3428.085 2299.000 ;
      LAYER met5 ;
        RECT 3403.035 2150.130 3406.285 2150.435 ;
        RECT 3424.835 2150.130 3424.840 2153.000 ;
      LAYER met5 ;
        RECT 3424.840 2151.730 3428.085 2153.000 ;
        RECT 3429.685 2151.730 3434.135 2299.000 ;
        RECT 3435.735 2151.730 3444.735 2299.000 ;
        RECT 3446.335 2151.730 3450.585 2299.000 ;
        RECT 3452.185 2151.730 3456.435 2299.000 ;
        RECT 3458.035 2151.730 3482.985 2299.000 ;
        RECT 3563.785 2153.000 3588.000 2299.000 ;
      LAYER met5 ;
        RECT 3484.585 2150.130 3588.000 2153.000 ;
        RECT 3390.135 2147.550 3588.000 2150.130 ;
        RECT 3390.135 2083.510 3491.520 2147.550 ;
        RECT 3555.545 2083.510 3588.000 2147.550 ;
        RECT 3390.135 2080.870 3588.000 2083.510 ;
        RECT 3403.035 2080.565 3406.285 2080.870 ;
        RECT 181.715 2065.130 184.965 2065.370 ;
        RECT 0.000 2063.400 197.865 2065.130 ;
        RECT 0.000 1997.600 31.390 2063.400 ;
        RECT 97.040 1997.600 197.865 2063.400 ;
        RECT 0.000 1990.870 197.865 1997.600 ;
        RECT 0.000 1988.000 103.415 1990.870 ;
        RECT 181.715 1990.565 184.965 1990.870 ;
      LAYER met5 ;
        RECT 0.000 1852.000 24.215 1988.000 ;
      LAYER met5 ;
        RECT 0.000 1849.130 103.415 1852.000 ;
      LAYER met5 ;
        RECT 105.015 1850.730 129.965 1989.270 ;
        RECT 131.565 1850.730 135.815 1989.270 ;
        RECT 137.415 1850.730 141.665 1989.270 ;
        RECT 143.265 1850.730 152.265 1989.270 ;
        RECT 153.865 1850.730 158.315 1989.270 ;
        RECT 159.915 1988.000 163.160 1989.270 ;
        RECT 159.915 1852.000 163.165 1988.000 ;
        RECT 159.915 1850.730 163.160 1852.000 ;
        RECT 164.765 1850.730 168.015 1989.270 ;
        RECT 169.615 1850.730 174.065 1989.270 ;
        RECT 175.665 1850.730 180.115 1989.270 ;
        RECT 181.715 1850.970 184.965 1988.965 ;
        RECT 186.565 1850.730 191.015 1989.270 ;
        RECT 192.615 1850.730 197.865 1989.270 ;
        RECT 3390.135 1931.730 3395.385 2079.270 ;
        RECT 3396.985 1931.730 3401.435 2079.270 ;
        RECT 3403.035 1932.035 3406.285 2078.965 ;
        RECT 3407.885 1931.730 3412.335 2079.270 ;
        RECT 3413.935 1931.730 3418.385 2079.270 ;
        RECT 3419.985 1931.730 3423.235 2079.270 ;
      LAYER met5 ;
        RECT 3424.835 2078.000 3424.840 2080.870 ;
      LAYER met5 ;
        RECT 3424.840 2078.000 3428.085 2079.270 ;
        RECT 3424.835 1933.000 3428.085 2078.000 ;
        RECT 3424.840 1931.730 3428.085 1933.000 ;
        RECT 3429.685 1931.730 3434.135 2079.270 ;
        RECT 3435.735 1931.730 3444.735 2079.270 ;
        RECT 3446.335 1931.730 3450.585 2079.270 ;
        RECT 3452.185 1931.730 3456.435 2079.270 ;
        RECT 3458.035 1931.730 3482.985 2079.270 ;
      LAYER met5 ;
        RECT 3484.585 2078.000 3588.000 2080.870 ;
      LAYER met5 ;
        RECT 3563.785 1933.000 3588.000 2078.000 ;
      LAYER met5 ;
        RECT 3403.035 1930.130 3406.285 1930.435 ;
        RECT 3484.585 1930.130 3588.000 1933.000 ;
        RECT 3390.135 1923.400 3588.000 1930.130 ;
        RECT 3390.135 1857.600 3490.960 1923.400 ;
        RECT 3556.610 1857.600 3588.000 1923.400 ;
        RECT 3390.135 1855.870 3588.000 1857.600 ;
        RECT 3403.035 1855.630 3406.285 1855.870 ;
        RECT 181.715 1849.130 184.965 1849.370 ;
        RECT 0.000 1847.400 197.865 1849.130 ;
        RECT 0.000 1781.600 31.390 1847.400 ;
        RECT 97.040 1781.600 197.865 1847.400 ;
        RECT 0.000 1774.870 197.865 1781.600 ;
        RECT 0.000 1772.000 103.415 1774.870 ;
        RECT 181.715 1774.565 184.965 1774.870 ;
      LAYER met5 ;
        RECT 0.000 1636.000 24.215 1772.000 ;
      LAYER met5 ;
        RECT 0.000 1633.130 103.415 1636.000 ;
      LAYER met5 ;
        RECT 105.015 1634.730 129.965 1773.270 ;
        RECT 131.565 1634.730 135.815 1773.270 ;
        RECT 137.415 1634.730 141.665 1773.270 ;
        RECT 143.265 1634.730 152.265 1773.270 ;
        RECT 153.865 1634.730 158.315 1773.270 ;
        RECT 159.915 1772.000 163.160 1773.270 ;
        RECT 159.915 1636.000 163.165 1772.000 ;
        RECT 159.915 1634.730 163.160 1636.000 ;
        RECT 164.765 1634.730 168.015 1773.270 ;
        RECT 169.615 1634.730 174.065 1773.270 ;
        RECT 175.665 1634.730 180.115 1773.270 ;
        RECT 181.715 1634.970 184.965 1772.965 ;
        RECT 186.565 1634.730 191.015 1773.270 ;
        RECT 192.615 1634.730 197.865 1773.270 ;
        RECT 3390.135 1705.730 3395.385 1854.270 ;
        RECT 3396.985 1705.730 3401.435 1854.270 ;
        RECT 3403.035 1706.035 3406.285 1854.030 ;
        RECT 3407.885 1705.730 3412.335 1854.270 ;
        RECT 3413.935 1705.730 3418.385 1854.270 ;
        RECT 3419.985 1705.730 3423.235 1854.270 ;
        RECT 3424.840 1853.000 3428.085 1854.270 ;
        RECT 3424.835 1707.000 3428.085 1853.000 ;
        RECT 3424.840 1705.730 3428.085 1707.000 ;
        RECT 3429.685 1705.730 3434.135 1854.270 ;
        RECT 3435.735 1705.730 3444.735 1854.270 ;
        RECT 3446.335 1705.730 3450.585 1854.270 ;
        RECT 3452.185 1705.730 3456.435 1854.270 ;
        RECT 3458.035 1705.730 3482.985 1854.270 ;
      LAYER met5 ;
        RECT 3484.585 1853.000 3588.000 1855.870 ;
      LAYER met5 ;
        RECT 3563.785 1707.000 3588.000 1853.000 ;
      LAYER met5 ;
        RECT 3403.035 1704.130 3406.285 1704.435 ;
        RECT 3484.585 1704.130 3588.000 1707.000 ;
        RECT 3390.135 1697.400 3588.000 1704.130 ;
        RECT 181.715 1633.130 184.965 1633.370 ;
        RECT 0.000 1631.400 197.865 1633.130 ;
        RECT 0.000 1565.600 31.390 1631.400 ;
        RECT 97.040 1565.600 197.865 1631.400 ;
        RECT 3390.135 1631.600 3490.960 1697.400 ;
        RECT 3556.610 1631.600 3588.000 1697.400 ;
        RECT 3390.135 1629.870 3588.000 1631.600 ;
        RECT 3403.035 1629.630 3406.285 1629.870 ;
        RECT 0.000 1558.870 197.865 1565.600 ;
        RECT 0.000 1556.000 103.415 1558.870 ;
        RECT 181.715 1558.565 184.965 1558.870 ;
      LAYER met5 ;
        RECT 0.000 1420.000 24.215 1556.000 ;
      LAYER met5 ;
        RECT 0.000 1417.130 103.415 1420.000 ;
      LAYER met5 ;
        RECT 105.015 1418.730 129.965 1557.270 ;
        RECT 131.565 1418.730 135.815 1557.270 ;
        RECT 137.415 1418.730 141.665 1557.270 ;
        RECT 143.265 1418.730 152.265 1557.270 ;
        RECT 153.865 1418.730 158.315 1557.270 ;
        RECT 159.915 1556.000 163.160 1557.270 ;
        RECT 159.915 1420.000 163.165 1556.000 ;
        RECT 159.915 1418.730 163.160 1420.000 ;
        RECT 164.765 1418.730 168.015 1557.270 ;
        RECT 169.615 1418.730 174.065 1557.270 ;
        RECT 175.665 1418.730 180.115 1557.270 ;
        RECT 181.715 1418.970 184.965 1556.965 ;
        RECT 186.565 1418.730 191.015 1557.270 ;
        RECT 192.615 1418.730 197.865 1557.270 ;
        RECT 3390.135 1480.730 3395.385 1628.270 ;
        RECT 3396.985 1480.730 3401.435 1628.270 ;
        RECT 3403.035 1481.035 3406.285 1628.030 ;
        RECT 3407.885 1480.730 3412.335 1628.270 ;
        RECT 3413.935 1480.730 3418.385 1628.270 ;
        RECT 3419.985 1480.730 3423.235 1628.270 ;
        RECT 3424.840 1627.000 3428.085 1628.270 ;
        RECT 3424.835 1482.000 3428.085 1627.000 ;
        RECT 3424.840 1480.730 3428.085 1482.000 ;
        RECT 3429.685 1480.730 3434.135 1628.270 ;
        RECT 3435.735 1480.730 3444.735 1628.270 ;
        RECT 3446.335 1480.730 3450.585 1628.270 ;
        RECT 3452.185 1480.730 3456.435 1628.270 ;
        RECT 3458.035 1480.730 3482.985 1628.270 ;
      LAYER met5 ;
        RECT 3484.585 1627.000 3588.000 1629.870 ;
      LAYER met5 ;
        RECT 3563.785 1482.000 3588.000 1627.000 ;
      LAYER met5 ;
        RECT 3403.035 1479.130 3406.285 1479.435 ;
        RECT 3484.585 1479.130 3588.000 1482.000 ;
        RECT 3390.135 1472.400 3588.000 1479.130 ;
        RECT 181.715 1417.130 184.965 1417.370 ;
        RECT 0.000 1415.400 197.865 1417.130 ;
        RECT 0.000 1349.600 31.390 1415.400 ;
        RECT 97.040 1349.600 197.865 1415.400 ;
        RECT 3390.135 1406.600 3490.960 1472.400 ;
        RECT 3556.610 1406.600 3588.000 1472.400 ;
        RECT 3390.135 1404.870 3588.000 1406.600 ;
        RECT 3403.035 1404.630 3406.285 1404.870 ;
        RECT 0.000 1342.870 197.865 1349.600 ;
        RECT 0.000 1340.000 103.415 1342.870 ;
        RECT 181.715 1342.565 184.965 1342.870 ;
      LAYER met5 ;
        RECT 0.000 1204.000 24.215 1340.000 ;
      LAYER met5 ;
        RECT 0.000 1201.130 103.415 1204.000 ;
      LAYER met5 ;
        RECT 105.015 1202.730 129.965 1341.270 ;
        RECT 131.565 1202.730 135.815 1341.270 ;
        RECT 137.415 1202.730 141.665 1341.270 ;
        RECT 143.265 1202.730 152.265 1341.270 ;
        RECT 153.865 1202.730 158.315 1341.270 ;
        RECT 159.915 1340.000 163.160 1341.270 ;
        RECT 159.915 1204.000 163.165 1340.000 ;
        RECT 159.915 1202.730 163.160 1204.000 ;
        RECT 164.765 1202.730 168.015 1341.270 ;
        RECT 169.615 1202.730 174.065 1341.270 ;
        RECT 175.665 1202.730 180.115 1341.270 ;
        RECT 181.715 1202.970 184.965 1340.965 ;
        RECT 186.565 1202.730 191.015 1341.270 ;
        RECT 192.615 1202.730 197.865 1341.270 ;
        RECT 3390.135 1255.730 3395.385 1403.270 ;
        RECT 3396.985 1255.730 3401.435 1403.270 ;
        RECT 3403.035 1256.035 3406.285 1403.030 ;
        RECT 3407.885 1255.730 3412.335 1403.270 ;
        RECT 3413.935 1255.730 3418.385 1403.270 ;
        RECT 3419.985 1255.730 3423.235 1403.270 ;
        RECT 3424.840 1402.000 3428.085 1403.270 ;
        RECT 3424.835 1257.000 3428.085 1402.000 ;
        RECT 3424.840 1255.730 3428.085 1257.000 ;
        RECT 3429.685 1255.730 3434.135 1403.270 ;
        RECT 3435.735 1255.730 3444.735 1403.270 ;
        RECT 3446.335 1255.730 3450.585 1403.270 ;
        RECT 3452.185 1255.730 3456.435 1403.270 ;
        RECT 3458.035 1255.730 3482.985 1403.270 ;
      LAYER met5 ;
        RECT 3484.585 1402.000 3588.000 1404.870 ;
      LAYER met5 ;
        RECT 3563.785 1257.000 3588.000 1402.000 ;
      LAYER met5 ;
        RECT 3403.035 1254.130 3406.285 1254.435 ;
        RECT 3484.585 1254.130 3588.000 1257.000 ;
        RECT 3390.135 1247.400 3588.000 1254.130 ;
        RECT 181.715 1201.130 184.965 1201.370 ;
        RECT 0.000 1199.400 197.865 1201.130 ;
        RECT 0.000 1133.600 31.390 1199.400 ;
        RECT 97.040 1133.600 197.865 1199.400 ;
        RECT 3390.135 1181.600 3490.960 1247.400 ;
        RECT 3556.610 1181.600 3588.000 1247.400 ;
        RECT 3390.135 1179.870 3588.000 1181.600 ;
        RECT 3403.035 1179.630 3406.285 1179.870 ;
        RECT 0.000 1126.870 197.865 1133.600 ;
        RECT 0.000 1124.000 103.415 1126.870 ;
        RECT 181.715 1126.565 184.965 1126.870 ;
      LAYER met5 ;
        RECT 0.000 988.000 24.215 1124.000 ;
      LAYER met5 ;
        RECT 0.000 985.130 103.415 988.000 ;
      LAYER met5 ;
        RECT 105.015 986.730 129.965 1125.270 ;
        RECT 131.565 986.730 135.815 1125.270 ;
        RECT 137.415 986.730 141.665 1125.270 ;
        RECT 143.265 986.730 152.265 1125.270 ;
        RECT 153.865 986.730 158.315 1125.270 ;
        RECT 159.915 1124.000 163.160 1125.270 ;
        RECT 159.915 988.000 163.165 1124.000 ;
        RECT 159.915 986.730 163.160 988.000 ;
        RECT 164.765 986.730 168.015 1125.270 ;
        RECT 169.615 986.730 174.065 1125.270 ;
        RECT 175.665 986.730 180.115 1125.270 ;
        RECT 181.715 986.970 184.965 1124.965 ;
        RECT 186.565 986.730 191.015 1125.270 ;
        RECT 192.615 986.730 197.865 1125.270 ;
        RECT 3390.135 1029.730 3395.385 1178.270 ;
        RECT 3396.985 1029.730 3401.435 1178.270 ;
        RECT 3403.035 1030.035 3406.285 1178.030 ;
        RECT 3407.885 1029.730 3412.335 1178.270 ;
        RECT 3413.935 1029.730 3418.385 1178.270 ;
        RECT 3419.985 1029.730 3423.235 1178.270 ;
        RECT 3424.840 1177.000 3428.085 1178.270 ;
        RECT 3424.835 1031.000 3428.085 1177.000 ;
        RECT 3424.840 1029.730 3428.085 1031.000 ;
        RECT 3429.685 1029.730 3434.135 1178.270 ;
        RECT 3435.735 1029.730 3444.735 1178.270 ;
        RECT 3446.335 1029.730 3450.585 1178.270 ;
        RECT 3452.185 1029.730 3456.435 1178.270 ;
        RECT 3458.035 1029.730 3482.985 1178.270 ;
      LAYER met5 ;
        RECT 3484.585 1177.000 3588.000 1179.870 ;
      LAYER met5 ;
        RECT 3563.785 1031.000 3588.000 1177.000 ;
      LAYER met5 ;
        RECT 3403.035 1028.130 3406.285 1028.435 ;
        RECT 3484.585 1028.130 3588.000 1031.000 ;
        RECT 3390.135 1021.400 3588.000 1028.130 ;
        RECT 181.715 985.130 184.965 985.370 ;
        RECT 0.000 983.400 197.865 985.130 ;
        RECT 0.000 917.600 31.390 983.400 ;
        RECT 97.040 917.600 197.865 983.400 ;
        RECT 3390.135 955.600 3490.960 1021.400 ;
        RECT 3556.610 955.600 3588.000 1021.400 ;
        RECT 3390.135 953.870 3588.000 955.600 ;
        RECT 3403.035 953.630 3406.285 953.870 ;
        RECT 0.000 910.870 197.865 917.600 ;
        RECT 0.000 908.000 103.415 910.870 ;
        RECT 181.715 910.565 184.965 910.870 ;
      LAYER met5 ;
        RECT 0.000 626.000 24.215 908.000 ;
      LAYER met5 ;
        RECT 0.000 623.130 103.415 626.000 ;
      LAYER met5 ;
        RECT 105.015 624.730 129.965 909.270 ;
        RECT 131.565 624.730 135.815 909.270 ;
        RECT 137.415 624.730 141.665 909.270 ;
        RECT 143.265 631.000 152.265 909.270 ;
        RECT 143.265 624.730 152.265 626.330 ;
        RECT 153.865 624.730 158.315 909.270 ;
        RECT 159.915 908.000 163.160 909.270 ;
        RECT 159.915 631.000 163.165 908.000 ;
        RECT 159.915 624.730 163.160 626.330 ;
      LAYER met5 ;
        RECT 163.160 623.130 163.165 626.000 ;
      LAYER met5 ;
        RECT 164.765 624.730 168.015 909.270 ;
        RECT 169.615 624.730 174.065 909.270 ;
        RECT 175.665 624.730 180.115 909.270 ;
        RECT 181.715 631.000 184.965 908.965 ;
        RECT 181.715 625.035 184.965 626.635 ;
        RECT 186.565 624.730 191.015 909.270 ;
        RECT 192.615 624.730 197.865 909.270 ;
        RECT 3390.135 804.730 3395.385 952.270 ;
        RECT 3396.985 804.730 3401.435 952.270 ;
        RECT 3403.035 805.035 3406.285 952.030 ;
        RECT 3407.885 804.730 3412.335 952.270 ;
        RECT 3413.935 804.730 3418.385 952.270 ;
        RECT 3419.985 804.730 3423.235 952.270 ;
        RECT 3424.840 951.000 3428.085 952.270 ;
        RECT 3424.835 806.000 3428.085 951.000 ;
        RECT 3424.840 804.730 3428.085 806.000 ;
        RECT 3429.685 804.730 3434.135 952.270 ;
        RECT 3435.735 804.730 3444.735 952.270 ;
        RECT 3446.335 804.730 3450.585 952.270 ;
        RECT 3452.185 804.730 3456.435 952.270 ;
        RECT 3458.035 804.730 3482.985 952.270 ;
      LAYER met5 ;
        RECT 3484.585 951.000 3588.000 953.870 ;
      LAYER met5 ;
        RECT 3563.785 806.000 3588.000 951.000 ;
      LAYER met5 ;
        RECT 3403.035 803.130 3406.285 803.435 ;
        RECT 3484.585 803.130 3588.000 806.000 ;
        RECT 3390.135 796.400 3588.000 803.130 ;
        RECT 3390.135 730.600 3490.960 796.400 ;
        RECT 3556.610 730.600 3588.000 796.400 ;
        RECT 3390.135 728.870 3588.000 730.600 ;
        RECT 3403.035 728.630 3406.285 728.870 ;
        RECT 181.715 623.130 184.965 623.435 ;
        RECT 0.000 620.490 197.865 623.130 ;
        RECT 0.000 556.450 32.455 620.490 ;
        RECT 96.480 556.450 197.865 620.490 ;
      LAYER met5 ;
        RECT 3390.135 578.730 3395.385 727.270 ;
        RECT 3396.985 578.730 3401.435 727.270 ;
        RECT 3403.035 579.035 3406.285 727.030 ;
        RECT 3407.885 578.730 3412.335 727.270 ;
        RECT 3413.935 578.730 3418.385 727.270 ;
        RECT 3419.985 578.730 3423.235 727.270 ;
        RECT 3424.840 726.000 3428.085 727.270 ;
        RECT 3424.835 580.000 3428.085 726.000 ;
        RECT 3424.840 578.730 3428.085 580.000 ;
        RECT 3429.685 578.730 3434.135 727.270 ;
        RECT 3435.735 578.730 3444.735 727.270 ;
        RECT 3446.335 578.730 3450.585 727.270 ;
        RECT 3452.185 578.730 3456.435 727.270 ;
        RECT 3458.035 578.730 3482.985 727.270 ;
      LAYER met5 ;
        RECT 3484.585 726.000 3588.000 728.870 ;
      LAYER met5 ;
        RECT 3563.785 580.000 3588.000 726.000 ;
      LAYER met5 ;
        RECT 3403.035 577.130 3406.285 577.435 ;
        RECT 3484.585 577.130 3588.000 580.000 ;
        RECT 0.000 553.870 197.865 556.450 ;
        RECT 3390.135 570.400 3588.000 577.130 ;
        RECT 0.000 551.000 103.415 553.870 ;
      LAYER met5 ;
        RECT 0.000 415.000 24.215 551.000 ;
      LAYER met5 ;
        RECT 0.000 412.130 103.415 415.000 ;
      LAYER met5 ;
        RECT 105.015 413.730 129.965 552.270 ;
        RECT 131.565 413.730 135.815 552.270 ;
        RECT 137.415 413.730 141.665 552.270 ;
        RECT 143.265 413.730 152.265 552.270 ;
        RECT 153.865 413.730 158.315 552.270 ;
        RECT 159.915 551.000 163.160 552.270 ;
      LAYER met5 ;
        RECT 163.160 551.000 163.165 553.870 ;
        RECT 181.715 553.565 184.965 553.870 ;
      LAYER met5 ;
        RECT 159.915 415.000 163.165 551.000 ;
        RECT 159.915 413.730 163.160 415.000 ;
      LAYER met5 ;
        RECT 163.160 412.130 163.165 415.000 ;
      LAYER met5 ;
        RECT 164.765 413.730 168.015 552.270 ;
        RECT 169.615 413.730 174.065 552.270 ;
        RECT 175.665 413.730 180.115 552.270 ;
        RECT 181.715 414.035 184.965 551.965 ;
        RECT 186.565 413.730 191.015 552.270 ;
        RECT 192.615 413.730 197.865 552.270 ;
      LAYER met5 ;
        RECT 3390.135 504.600 3490.960 570.400 ;
        RECT 3556.610 504.600 3588.000 570.400 ;
        RECT 3390.135 502.870 3588.000 504.600 ;
        RECT 3403.035 502.630 3406.285 502.870 ;
        RECT 181.715 412.130 184.965 412.435 ;
        RECT 0.000 406.270 197.865 412.130 ;
        RECT 0.000 348.670 29.235 406.270 ;
        RECT 99.700 348.670 197.865 406.270 ;
        RECT 0.000 342.870 197.865 348.670 ;
        RECT 0.000 340.000 103.415 342.870 ;
      LAYER met5 ;
        RECT 0.000 204.000 24.215 340.000 ;
      LAYER met5 ;
        RECT 0.000 200.545 103.415 204.000 ;
      LAYER met5 ;
        RECT 105.015 202.145 129.965 341.270 ;
        RECT 131.565 202.730 135.815 341.270 ;
        RECT 137.415 202.730 141.665 341.270 ;
      LAYER met5 ;
        RECT 131.565 200.545 141.665 201.130 ;
        RECT 0.000 175.245 141.665 200.545 ;
      LAYER met5 ;
        RECT 143.265 176.845 152.265 341.270 ;
        RECT 153.865 202.730 158.315 341.270 ;
        RECT 159.915 340.000 163.160 341.270 ;
      LAYER met5 ;
        RECT 163.160 340.000 163.165 342.870 ;
        RECT 181.715 342.565 184.965 342.870 ;
      LAYER met5 ;
        RECT 159.915 204.000 163.165 340.000 ;
        RECT 159.915 202.730 163.160 204.000 ;
        RECT 164.765 202.730 168.015 341.270 ;
        RECT 169.615 202.730 174.065 341.270 ;
        RECT 175.665 202.730 180.115 341.270 ;
        RECT 181.715 202.745 184.965 340.965 ;
        RECT 186.565 202.730 191.015 341.270 ;
        RECT 192.615 202.730 197.865 341.270 ;
      LAYER met5 ;
        RECT 181.715 201.130 184.965 201.145 ;
        RECT 199.465 201.130 200.000 204.000 ;
        RECT 153.865 199.465 200.000 201.130 ;
        RECT 3384.000 199.465 3388.535 200.000 ;
        RECT 153.865 192.615 196.050 199.465 ;
        RECT 197.865 197.865 198.400 199.465 ;
        POLYGON 198.400 199.465 200.000 197.865 198.400 197.865 ;
        RECT 3386.870 198.400 3388.535 199.465 ;
        POLYGON 3390.135 200.000 3390.135 198.400 3388.535 198.400 ;
        RECT 3386.870 197.865 3390.135 198.400 ;
      LAYER met5 ;
        RECT 197.650 192.615 395.270 197.865 ;
      LAYER met5 ;
        RECT 153.865 184.965 194.615 192.615 ;
      LAYER met5 ;
        RECT 237.000 191.015 357.000 192.615 ;
        RECT 196.215 186.565 395.270 191.015 ;
      LAYER met5 ;
        RECT 396.870 184.965 466.130 197.865 ;
      LAYER met5 ;
        RECT 467.730 192.615 664.270 197.865 ;
        RECT 506.000 191.015 626.000 192.615 ;
        RECT 467.730 186.565 664.270 191.015 ;
      LAYER met5 ;
        RECT 665.870 184.965 735.130 197.865 ;
      LAYER met5 ;
        RECT 736.730 192.615 933.270 197.865 ;
        RECT 775.000 191.015 895.000 192.615 ;
        RECT 736.730 186.565 933.270 191.015 ;
      LAYER met5 ;
        RECT 934.870 184.965 1009.130 197.865 ;
      LAYER met5 ;
        RECT 1010.730 192.615 1207.270 197.865 ;
        RECT 1049.000 191.015 1169.000 192.615 ;
        RECT 1010.730 186.565 1207.270 191.015 ;
      LAYER met5 ;
        RECT 1208.870 184.965 1278.130 197.865 ;
      LAYER met5 ;
        RECT 1279.730 192.615 1476.270 197.865 ;
        RECT 1318.000 191.015 1438.000 192.615 ;
        RECT 1279.730 186.565 1476.270 191.015 ;
      LAYER met5 ;
        RECT 1477.870 184.965 1552.130 197.865 ;
      LAYER met5 ;
        RECT 1553.730 192.615 1750.270 197.865 ;
        RECT 1592.000 191.015 1712.000 192.615 ;
        RECT 1553.730 186.565 1750.270 191.015 ;
      LAYER met5 ;
        RECT 1751.870 184.965 1826.130 197.865 ;
      LAYER met5 ;
        RECT 1827.730 192.615 2024.270 197.865 ;
        RECT 1866.000 191.015 1986.000 192.615 ;
        RECT 1827.730 186.565 2024.270 191.015 ;
      LAYER met5 ;
        RECT 2025.870 184.965 2100.130 197.865 ;
      LAYER met5 ;
        RECT 2101.730 192.615 2298.270 197.865 ;
        RECT 2140.000 191.015 2260.000 192.615 ;
        RECT 2101.730 186.565 2298.270 191.015 ;
      LAYER met5 ;
        RECT 2299.870 184.965 2374.130 197.865 ;
      LAYER met5 ;
        RECT 2375.730 192.615 2572.270 197.865 ;
        RECT 2414.000 191.015 2534.000 192.615 ;
        RECT 2375.730 186.565 2572.270 191.015 ;
      LAYER met5 ;
        RECT 2573.870 184.965 2648.130 197.865 ;
      LAYER met5 ;
        RECT 2649.730 192.615 2846.270 197.865 ;
        RECT 2688.000 191.015 2808.000 192.615 ;
        RECT 2649.730 186.565 2846.270 191.015 ;
      LAYER met5 ;
        RECT 2847.870 184.965 2917.130 197.865 ;
      LAYER met5 ;
        RECT 2918.730 192.615 3115.270 197.865 ;
        RECT 2957.000 191.015 3077.000 192.615 ;
        RECT 2918.730 186.565 3115.270 191.015 ;
      LAYER met5 ;
        RECT 3116.870 184.965 3186.130 197.865 ;
      LAYER met5 ;
        RECT 3187.730 192.615 3385.270 197.865 ;
      LAYER met5 ;
        RECT 3386.870 196.050 3388.535 197.865 ;
      LAYER met5 ;
        RECT 3390.135 197.650 3395.385 501.270 ;
        RECT 3396.985 196.215 3401.435 501.270 ;
        RECT 3403.035 350.000 3406.285 501.030 ;
        RECT 3403.035 198.530 3406.285 345.000 ;
        RECT 3407.885 198.475 3412.335 501.270 ;
        RECT 3413.935 198.400 3418.385 501.270 ;
        RECT 3419.985 198.615 3423.235 501.270 ;
        RECT 3424.840 500.000 3428.085 501.270 ;
        RECT 3424.835 350.000 3428.085 500.000 ;
        RECT 3424.835 198.665 3428.085 345.000 ;
        RECT 3429.685 198.525 3434.135 501.270 ;
        RECT 3435.735 350.000 3444.735 501.270 ;
      LAYER met5 ;
        RECT 3424.835 197.015 3428.085 197.065 ;
        RECT 3403.035 196.875 3406.285 196.930 ;
        RECT 3419.985 196.925 3428.085 197.015 ;
        RECT 3403.035 196.800 3412.335 196.875 ;
        RECT 3419.985 196.800 3434.135 196.925 ;
        RECT 3386.870 194.615 3395.385 196.050 ;
        RECT 3403.035 194.615 3434.135 196.800 ;
      LAYER met5 ;
        RECT 3226.000 191.015 3346.000 192.615 ;
        RECT 3187.730 186.565 3385.270 191.015 ;
      LAYER met5 ;
        RECT 3386.870 184.965 3434.135 194.615 ;
        RECT 153.865 181.715 196.930 184.965 ;
      LAYER met5 ;
        RECT 198.530 181.715 394.965 184.965 ;
      LAYER met5 ;
        RECT 396.565 181.715 466.435 184.965 ;
      LAYER met5 ;
        RECT 468.035 181.715 663.965 184.965 ;
      LAYER met5 ;
        RECT 665.565 181.715 735.435 184.965 ;
      LAYER met5 ;
        RECT 737.035 181.715 933.030 184.965 ;
      LAYER met5 ;
        RECT 934.630 181.715 1009.435 184.965 ;
      LAYER met5 ;
        RECT 1011.035 181.715 1206.965 184.965 ;
      LAYER met5 ;
        RECT 1208.565 181.715 1278.435 184.965 ;
      LAYER met5 ;
        RECT 1280.035 181.715 1476.030 184.965 ;
      LAYER met5 ;
        RECT 1477.630 181.715 1552.435 184.965 ;
      LAYER met5 ;
        RECT 1554.035 181.715 1750.030 184.965 ;
      LAYER met5 ;
        RECT 1751.630 181.715 1826.435 184.965 ;
      LAYER met5 ;
        RECT 1828.035 181.715 2024.030 184.965 ;
      LAYER met5 ;
        RECT 2025.630 181.715 2100.435 184.965 ;
      LAYER met5 ;
        RECT 2102.035 181.715 2298.030 184.965 ;
      LAYER met5 ;
        RECT 2299.630 181.715 2374.435 184.965 ;
      LAYER met5 ;
        RECT 2376.035 181.715 2572.030 184.965 ;
      LAYER met5 ;
        RECT 2573.630 181.715 2648.435 184.965 ;
      LAYER met5 ;
        RECT 2650.035 181.715 2845.965 184.965 ;
      LAYER met5 ;
        RECT 2847.565 181.715 2917.435 184.965 ;
      LAYER met5 ;
        RECT 2919.035 181.715 3114.965 184.965 ;
      LAYER met5 ;
        RECT 3116.565 181.715 3186.435 184.965 ;
      LAYER met5 ;
        RECT 3188.035 181.715 3385.255 184.965 ;
      LAYER met5 ;
        RECT 3386.855 181.715 3434.135 184.965 ;
        RECT 153.865 175.665 196.875 181.715 ;
      LAYER met5 ;
        RECT 198.475 175.665 395.270 180.115 ;
      LAYER met5 ;
        RECT 153.865 175.245 196.800 175.665 ;
        RECT 0.000 168.015 196.800 175.245 ;
      LAYER met5 ;
        RECT 198.400 169.615 395.270 174.065 ;
      LAYER met5 ;
        RECT 0.000 163.165 197.015 168.015 ;
      LAYER met5 ;
        RECT 198.615 164.765 395.270 168.015 ;
      LAYER met5 ;
        RECT 396.870 163.165 466.130 181.715 ;
      LAYER met5 ;
        RECT 467.730 175.665 664.270 180.115 ;
        RECT 467.730 169.615 664.270 174.065 ;
        RECT 467.730 164.765 664.270 168.015 ;
      LAYER met5 ;
        RECT 0.000 159.915 197.065 163.165 ;
      LAYER met5 ;
        RECT 198.665 163.160 394.000 163.165 ;
      LAYER met5 ;
        RECT 394.000 163.160 469.000 163.165 ;
      LAYER met5 ;
        RECT 469.000 163.160 663.000 163.165 ;
        RECT 198.665 159.915 395.270 163.160 ;
      LAYER met5 ;
        RECT 0.000 153.865 196.925 159.915 ;
      LAYER met5 ;
        RECT 198.525 153.865 395.270 158.315 ;
      LAYER met5 ;
        RECT 0.000 141.665 175.245 153.865 ;
      LAYER met5 ;
        RECT 176.845 143.265 395.270 152.265 ;
      LAYER met5 ;
        RECT 0.000 135.815 196.775 141.665 ;
      LAYER met5 ;
        RECT 198.375 137.415 395.270 141.665 ;
      LAYER met5 ;
        RECT 0.000 131.565 196.920 135.815 ;
      LAYER met5 ;
        RECT 198.520 131.565 395.270 135.815 ;
      LAYER met5 ;
        RECT 0.000 103.415 195.755 131.565 ;
      LAYER met5 ;
        RECT 197.355 105.015 395.270 129.965 ;
      LAYER met5 ;
        RECT 396.870 103.415 466.130 163.160 ;
      LAYER met5 ;
        RECT 467.730 159.915 664.270 163.160 ;
        RECT 467.730 153.865 664.270 158.315 ;
        RECT 467.730 143.265 664.270 152.265 ;
        RECT 467.730 137.415 664.270 141.665 ;
        RECT 467.730 131.565 664.270 135.815 ;
        RECT 467.730 105.015 664.270 129.965 ;
      LAYER met5 ;
        RECT 665.870 103.415 735.130 181.715 ;
      LAYER met5 ;
        RECT 736.730 175.665 933.270 180.115 ;
        RECT 736.730 169.615 933.270 174.065 ;
        RECT 736.730 164.765 933.270 168.015 ;
        RECT 738.000 163.160 932.000 163.165 ;
        RECT 736.730 159.915 933.270 163.160 ;
        RECT 736.730 153.865 933.270 158.315 ;
        RECT 736.730 143.265 933.270 152.265 ;
        RECT 736.730 137.415 933.270 141.665 ;
        RECT 736.730 131.565 933.270 135.815 ;
        RECT 736.730 105.015 933.270 129.965 ;
      LAYER met5 ;
        RECT 934.870 103.415 1009.130 181.715 ;
      LAYER met5 ;
        RECT 1010.730 175.665 1207.270 180.115 ;
        RECT 1010.730 169.615 1207.270 174.065 ;
        RECT 1010.730 164.765 1207.270 168.015 ;
      LAYER met5 ;
        RECT 1208.870 163.165 1278.130 181.715 ;
      LAYER met5 ;
        RECT 1279.730 175.665 1476.270 180.115 ;
        RECT 1279.730 169.615 1476.270 174.065 ;
        RECT 1279.730 164.765 1476.270 168.015 ;
        RECT 1012.000 163.160 1206.000 163.165 ;
      LAYER met5 ;
        RECT 1206.000 163.160 1281.000 163.165 ;
      LAYER met5 ;
        RECT 1281.000 163.160 1475.000 163.165 ;
        RECT 1010.730 159.915 1207.270 163.160 ;
        RECT 1010.730 153.865 1207.270 158.315 ;
        RECT 1010.730 143.265 1207.270 152.265 ;
        RECT 1010.730 137.415 1207.270 141.665 ;
        RECT 1010.730 131.565 1207.270 135.815 ;
        RECT 1010.730 105.015 1207.270 129.965 ;
      LAYER met5 ;
        RECT 1208.870 103.415 1278.130 163.160 ;
      LAYER met5 ;
        RECT 1279.730 159.915 1476.270 163.160 ;
        RECT 1279.730 153.865 1476.270 158.315 ;
        RECT 1279.730 143.265 1476.270 152.265 ;
        RECT 1279.730 137.415 1476.270 141.665 ;
        RECT 1279.730 131.565 1476.270 135.815 ;
        RECT 1279.730 105.015 1476.270 129.965 ;
      LAYER met5 ;
        RECT 1477.870 103.415 1552.130 181.715 ;
      LAYER met5 ;
        RECT 1553.730 175.665 1750.270 180.115 ;
        RECT 1553.730 169.615 1750.270 174.065 ;
        RECT 1553.730 164.765 1750.270 168.015 ;
        RECT 1555.000 163.160 1749.000 163.165 ;
        RECT 1553.730 159.915 1750.270 163.160 ;
        RECT 1553.730 153.865 1750.270 158.315 ;
        RECT 1553.730 143.265 1750.270 152.265 ;
        RECT 1553.730 137.415 1750.270 141.665 ;
        RECT 1553.730 131.565 1750.270 135.815 ;
        RECT 1553.730 105.015 1750.270 129.965 ;
      LAYER met5 ;
        RECT 1751.870 103.415 1826.130 181.715 ;
      LAYER met5 ;
        RECT 1827.730 175.665 2024.270 180.115 ;
        RECT 1827.730 169.615 2024.270 174.065 ;
        RECT 1827.730 164.765 2024.270 168.015 ;
        RECT 1829.000 163.160 2023.000 163.165 ;
        RECT 1827.730 159.915 2024.270 163.160 ;
        RECT 1827.730 153.865 2024.270 158.315 ;
        RECT 1827.730 143.265 2024.270 152.265 ;
        RECT 1827.730 137.415 2024.270 141.665 ;
        RECT 1827.730 131.565 2024.270 135.815 ;
        RECT 1827.730 105.015 2024.270 129.965 ;
      LAYER met5 ;
        RECT 2025.870 103.415 2100.130 181.715 ;
      LAYER met5 ;
        RECT 2101.730 175.665 2298.270 180.115 ;
        RECT 2101.730 169.615 2298.270 174.065 ;
        RECT 2101.730 164.765 2298.270 168.015 ;
        RECT 2103.000 163.160 2297.000 163.165 ;
        RECT 2101.730 159.915 2298.270 163.160 ;
        RECT 2101.730 153.865 2298.270 158.315 ;
        RECT 2101.730 143.265 2298.270 152.265 ;
        RECT 2101.730 137.415 2298.270 141.665 ;
        RECT 2101.730 131.565 2298.270 135.815 ;
        RECT 2101.730 105.015 2298.270 129.965 ;
      LAYER met5 ;
        RECT 2299.870 103.415 2374.130 181.715 ;
      LAYER met5 ;
        RECT 2375.730 175.665 2572.270 180.115 ;
        RECT 2375.730 169.615 2572.270 174.065 ;
        RECT 2375.730 164.765 2572.270 168.015 ;
        RECT 2377.000 163.160 2571.000 163.165 ;
        RECT 2375.730 159.915 2572.270 163.160 ;
        RECT 2375.730 153.865 2572.270 158.315 ;
        RECT 2375.730 143.265 2572.270 152.265 ;
        RECT 2375.730 137.415 2572.270 141.665 ;
        RECT 2375.730 131.565 2572.270 135.815 ;
        RECT 2375.730 105.015 2572.270 129.965 ;
      LAYER met5 ;
        RECT 2573.870 103.415 2648.130 181.715 ;
      LAYER met5 ;
        RECT 2649.730 175.665 2846.270 180.115 ;
        RECT 2649.730 169.615 2846.270 174.065 ;
        RECT 2649.730 164.765 2846.270 168.015 ;
      LAYER met5 ;
        RECT 2847.870 163.165 2917.130 181.715 ;
      LAYER met5 ;
        RECT 2918.730 175.665 3115.270 180.115 ;
        RECT 2918.730 169.615 3115.270 174.065 ;
        RECT 2918.730 164.765 3115.270 168.015 ;
      LAYER met5 ;
        RECT 3116.870 163.165 3186.130 181.715 ;
      LAYER met5 ;
        RECT 3187.730 175.665 3385.270 180.115 ;
      LAYER met5 ;
        RECT 3386.870 175.245 3434.135 181.715 ;
      LAYER met5 ;
        RECT 3435.735 176.845 3444.735 345.000 ;
        RECT 3446.335 198.375 3450.585 501.270 ;
        RECT 3452.185 198.520 3456.435 501.270 ;
        RECT 3458.035 197.355 3482.985 501.270 ;
      LAYER met5 ;
        RECT 3484.585 500.000 3588.000 502.870 ;
      LAYER met5 ;
        RECT 3563.785 200.000 3588.000 500.000 ;
      LAYER met5 ;
        RECT 3452.185 196.775 3456.435 196.920 ;
        RECT 3446.335 195.755 3456.435 196.775 ;
        RECT 3484.585 195.755 3588.000 200.000 ;
        RECT 3446.335 175.245 3588.000 195.755 ;
      LAYER met5 ;
        RECT 3187.730 169.615 3385.270 174.065 ;
        RECT 3187.730 164.765 3385.270 168.015 ;
        RECT 2651.000 163.160 2845.000 163.165 ;
      LAYER met5 ;
        RECT 2845.000 163.160 2920.000 163.165 ;
      LAYER met5 ;
        RECT 2920.000 163.160 3114.000 163.165 ;
      LAYER met5 ;
        RECT 3114.000 163.160 3189.000 163.165 ;
      LAYER met5 ;
        RECT 3189.000 163.160 3384.000 163.165 ;
        RECT 2649.730 159.915 2846.270 163.160 ;
        RECT 2649.730 153.865 2846.270 158.315 ;
        RECT 2649.730 143.265 2846.270 152.265 ;
        RECT 2649.730 137.415 2846.270 141.665 ;
        RECT 2649.730 131.565 2846.270 135.815 ;
        RECT 2649.730 105.015 2846.270 129.965 ;
      LAYER met5 ;
        RECT 2847.870 103.415 2917.130 163.160 ;
      LAYER met5 ;
        RECT 2918.730 159.915 3115.270 163.160 ;
        RECT 2918.730 153.865 3115.270 158.315 ;
        RECT 2918.730 143.265 3115.270 152.265 ;
        RECT 2918.730 137.415 3115.270 141.665 ;
        RECT 2918.730 131.565 3115.270 135.815 ;
        RECT 2918.730 105.015 3115.270 129.965 ;
      LAYER met5 ;
        RECT 3116.870 103.415 3186.130 163.160 ;
      LAYER met5 ;
        RECT 3187.730 159.915 3385.270 163.160 ;
        RECT 3187.730 153.865 3385.270 158.315 ;
      LAYER met5 ;
        RECT 3386.870 153.865 3588.000 175.245 ;
      LAYER met5 ;
        RECT 3187.730 143.265 3411.155 152.265 ;
      LAYER met5 ;
        RECT 3412.755 141.665 3588.000 153.865 ;
      LAYER met5 ;
        RECT 3187.730 137.415 3385.270 141.665 ;
        RECT 3187.730 131.565 3385.270 135.815 ;
      LAYER met5 ;
        RECT 3386.870 131.565 3588.000 141.665 ;
      LAYER met5 ;
        RECT 3187.730 105.015 3385.855 129.965 ;
      LAYER met5 ;
        RECT 3387.455 103.415 3588.000 131.565 ;
        RECT 0.000 0.000 200.000 103.415 ;
        RECT 394.000 96.480 469.000 103.415 ;
        RECT 394.000 32.455 399.510 96.480 ;
        RECT 463.550 32.455 469.000 96.480 ;
      LAYER met5 ;
        RECT 200.000 0.000 394.000 24.215 ;
      LAYER met5 ;
        RECT 394.000 0.000 469.000 32.455 ;
        RECT 663.000 93.145 738.000 103.415 ;
        RECT 663.000 34.115 681.965 93.145 ;
        RECT 722.350 34.115 738.000 93.145 ;
        RECT 663.000 25.815 738.000 34.115 ;
        RECT 932.000 97.040 1012.000 103.415 ;
        RECT 932.000 31.390 936.600 97.040 ;
        RECT 1002.400 31.390 1012.000 97.040 ;
      LAYER met5 ;
        RECT 469.000 0.000 664.270 24.215 ;
      LAYER met5 ;
        RECT 665.870 0.000 735.130 25.815 ;
      LAYER met5 ;
        RECT 736.730 0.000 932.000 24.215 ;
      LAYER met5 ;
        RECT 932.000 0.000 1012.000 31.390 ;
        RECT 1206.000 99.700 1281.000 103.415 ;
        RECT 1206.000 29.235 1214.730 99.700 ;
        RECT 1272.330 29.235 1281.000 99.700 ;
      LAYER met5 ;
        RECT 1012.000 0.000 1206.000 24.215 ;
      LAYER met5 ;
        RECT 1206.000 0.000 1281.000 29.235 ;
        RECT 1475.000 97.040 1555.000 103.415 ;
        RECT 1475.000 31.390 1479.600 97.040 ;
        RECT 1545.400 31.390 1555.000 97.040 ;
      LAYER met5 ;
        RECT 1281.000 0.000 1475.000 24.215 ;
      LAYER met5 ;
        RECT 1475.000 0.000 1555.000 31.390 ;
        RECT 1749.000 97.040 1829.000 103.415 ;
        RECT 1749.000 31.390 1753.600 97.040 ;
        RECT 1819.400 31.390 1829.000 97.040 ;
      LAYER met5 ;
        RECT 1555.000 0.000 1749.000 24.215 ;
      LAYER met5 ;
        RECT 1749.000 0.000 1829.000 31.390 ;
        RECT 2023.000 97.040 2103.000 103.415 ;
        RECT 2023.000 31.390 2027.600 97.040 ;
        RECT 2093.400 31.390 2103.000 97.040 ;
      LAYER met5 ;
        RECT 1829.000 0.000 2023.000 24.215 ;
      LAYER met5 ;
        RECT 2023.000 0.000 2103.000 31.390 ;
        RECT 2297.000 97.040 2377.000 103.415 ;
        RECT 2297.000 31.390 2301.600 97.040 ;
        RECT 2367.400 31.390 2377.000 97.040 ;
      LAYER met5 ;
        RECT 2103.000 0.000 2297.000 24.215 ;
      LAYER met5 ;
        RECT 2297.000 0.000 2377.000 31.390 ;
        RECT 2571.000 97.040 2651.000 103.415 ;
        RECT 2571.000 31.390 2575.600 97.040 ;
        RECT 2641.400 31.390 2651.000 97.040 ;
      LAYER met5 ;
        RECT 2377.000 0.000 2571.000 24.215 ;
      LAYER met5 ;
        RECT 2571.000 0.000 2651.000 31.390 ;
        RECT 2845.000 96.480 2920.000 103.415 ;
        RECT 2845.000 32.455 2850.510 96.480 ;
        RECT 2914.550 32.455 2920.000 96.480 ;
      LAYER met5 ;
        RECT 2651.000 0.000 2845.000 24.215 ;
      LAYER met5 ;
        RECT 2845.000 0.000 2920.000 32.455 ;
        RECT 3114.000 96.480 3189.000 103.415 ;
        RECT 3114.000 32.455 3119.510 96.480 ;
        RECT 3183.550 32.455 3189.000 96.480 ;
      LAYER met5 ;
        RECT 2920.000 0.000 3114.000 24.215 ;
      LAYER met5 ;
        RECT 3114.000 0.000 3189.000 32.455 ;
      LAYER met5 ;
        RECT 3189.000 0.000 3384.000 24.215 ;
      LAYER met5 ;
        RECT 3384.000 0.000 3588.000 103.415 ;
  END
END chip_io_alt
END LIBRARY

