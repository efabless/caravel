// This is the unpowered netlist.
module mgmt_protect (caravel_clk,
    caravel_clk2,
    caravel_rstn,
    mprj_ack_i_core,
    mprj_ack_i_user,
    mprj_cyc_o_core,
    mprj_cyc_o_user,
    mprj_iena_wb,
    mprj_stb_o_core,
    mprj_stb_o_user,
    mprj_we_o_core,
    mprj_we_o_user,
    user1_vcc_powergood,
    user1_vdd_powergood,
    user2_vcc_powergood,
    user2_vdd_powergood,
    user_clock,
    user_clock2,
    user_reset,
    la_data_in_core,
    la_data_in_mprj,
    la_data_out_core,
    la_data_out_mprj,
    la_iena_mprj,
    la_oenb_core,
    la_oenb_mprj,
    mprj_adr_o_core,
    mprj_adr_o_user,
    mprj_dat_i_core,
    mprj_dat_i_user,
    mprj_dat_o_core,
    mprj_dat_o_user,
    mprj_sel_o_core,
    mprj_sel_o_user,
    user_irq,
    user_irq_core,
    user_irq_ena);
 input caravel_clk;
 input caravel_clk2;
 input caravel_rstn;
 output mprj_ack_i_core;
 input mprj_ack_i_user;
 input mprj_cyc_o_core;
 output mprj_cyc_o_user;
 input mprj_iena_wb;
 input mprj_stb_o_core;
 output mprj_stb_o_user;
 input mprj_we_o_core;
 output mprj_we_o_user;
 output user1_vcc_powergood;
 output user1_vdd_powergood;
 output user2_vcc_powergood;
 output user2_vdd_powergood;
 output user_clock;
 output user_clock2;
 output user_reset;
 output [127:0] la_data_in_core;
 output [127:0] la_data_in_mprj;
 input [127:0] la_data_out_core;
 input [127:0] la_data_out_mprj;
 input [127:0] la_iena_mprj;
 output [127:0] la_oenb_core;
 input [127:0] la_oenb_mprj;
 input [31:0] mprj_adr_o_core;
 output [31:0] mprj_adr_o_user;
 output [31:0] mprj_dat_i_core;
 input [31:0] mprj_dat_i_user;
 input [31:0] mprj_dat_o_core;
 output [31:0] mprj_dat_o_user;
 input [3:0] mprj_sel_o_core;
 output [3:0] mprj_sel_o_user;
 output [2:0] user_irq;
 input [2:0] user_irq_core;
 input [2:0] user_irq_ena;

 wire \la_data_in_enable[0] ;
 wire \la_data_in_enable[100] ;
 wire \la_data_in_enable[101] ;
 wire \la_data_in_enable[102] ;
 wire \la_data_in_enable[103] ;
 wire \la_data_in_enable[104] ;
 wire \la_data_in_enable[105] ;
 wire \la_data_in_enable[106] ;
 wire \la_data_in_enable[107] ;
 wire \la_data_in_enable[108] ;
 wire \la_data_in_enable[109] ;
 wire \la_data_in_enable[10] ;
 wire \la_data_in_enable[110] ;
 wire \la_data_in_enable[111] ;
 wire \la_data_in_enable[112] ;
 wire \la_data_in_enable[113] ;
 wire \la_data_in_enable[114] ;
 wire \la_data_in_enable[115] ;
 wire \la_data_in_enable[116] ;
 wire \la_data_in_enable[117] ;
 wire \la_data_in_enable[118] ;
 wire \la_data_in_enable[119] ;
 wire \la_data_in_enable[11] ;
 wire \la_data_in_enable[120] ;
 wire \la_data_in_enable[121] ;
 wire \la_data_in_enable[122] ;
 wire \la_data_in_enable[123] ;
 wire \la_data_in_enable[124] ;
 wire \la_data_in_enable[125] ;
 wire \la_data_in_enable[126] ;
 wire \la_data_in_enable[127] ;
 wire \la_data_in_enable[12] ;
 wire \la_data_in_enable[13] ;
 wire \la_data_in_enable[14] ;
 wire \la_data_in_enable[15] ;
 wire \la_data_in_enable[16] ;
 wire \la_data_in_enable[17] ;
 wire \la_data_in_enable[18] ;
 wire \la_data_in_enable[19] ;
 wire \la_data_in_enable[1] ;
 wire \la_data_in_enable[20] ;
 wire \la_data_in_enable[21] ;
 wire \la_data_in_enable[22] ;
 wire \la_data_in_enable[23] ;
 wire \la_data_in_enable[24] ;
 wire \la_data_in_enable[25] ;
 wire \la_data_in_enable[26] ;
 wire \la_data_in_enable[27] ;
 wire \la_data_in_enable[28] ;
 wire \la_data_in_enable[29] ;
 wire \la_data_in_enable[2] ;
 wire \la_data_in_enable[30] ;
 wire \la_data_in_enable[31] ;
 wire \la_data_in_enable[32] ;
 wire \la_data_in_enable[33] ;
 wire \la_data_in_enable[34] ;
 wire \la_data_in_enable[35] ;
 wire \la_data_in_enable[36] ;
 wire \la_data_in_enable[37] ;
 wire \la_data_in_enable[38] ;
 wire \la_data_in_enable[39] ;
 wire \la_data_in_enable[3] ;
 wire \la_data_in_enable[40] ;
 wire \la_data_in_enable[41] ;
 wire \la_data_in_enable[42] ;
 wire \la_data_in_enable[43] ;
 wire \la_data_in_enable[44] ;
 wire \la_data_in_enable[45] ;
 wire \la_data_in_enable[46] ;
 wire \la_data_in_enable[47] ;
 wire \la_data_in_enable[48] ;
 wire \la_data_in_enable[49] ;
 wire \la_data_in_enable[4] ;
 wire \la_data_in_enable[50] ;
 wire \la_data_in_enable[51] ;
 wire \la_data_in_enable[52] ;
 wire \la_data_in_enable[53] ;
 wire \la_data_in_enable[54] ;
 wire \la_data_in_enable[55] ;
 wire \la_data_in_enable[56] ;
 wire \la_data_in_enable[57] ;
 wire \la_data_in_enable[58] ;
 wire \la_data_in_enable[59] ;
 wire \la_data_in_enable[5] ;
 wire \la_data_in_enable[60] ;
 wire \la_data_in_enable[61] ;
 wire \la_data_in_enable[62] ;
 wire \la_data_in_enable[63] ;
 wire \la_data_in_enable[64] ;
 wire \la_data_in_enable[65] ;
 wire \la_data_in_enable[66] ;
 wire \la_data_in_enable[67] ;
 wire \la_data_in_enable[68] ;
 wire \la_data_in_enable[69] ;
 wire \la_data_in_enable[6] ;
 wire \la_data_in_enable[70] ;
 wire \la_data_in_enable[71] ;
 wire \la_data_in_enable[72] ;
 wire \la_data_in_enable[73] ;
 wire \la_data_in_enable[74] ;
 wire \la_data_in_enable[75] ;
 wire \la_data_in_enable[76] ;
 wire \la_data_in_enable[77] ;
 wire \la_data_in_enable[78] ;
 wire \la_data_in_enable[79] ;
 wire \la_data_in_enable[7] ;
 wire \la_data_in_enable[80] ;
 wire \la_data_in_enable[81] ;
 wire \la_data_in_enable[82] ;
 wire \la_data_in_enable[83] ;
 wire \la_data_in_enable[84] ;
 wire \la_data_in_enable[85] ;
 wire \la_data_in_enable[86] ;
 wire \la_data_in_enable[87] ;
 wire \la_data_in_enable[88] ;
 wire \la_data_in_enable[89] ;
 wire \la_data_in_enable[8] ;
 wire \la_data_in_enable[90] ;
 wire \la_data_in_enable[91] ;
 wire \la_data_in_enable[92] ;
 wire \la_data_in_enable[93] ;
 wire \la_data_in_enable[94] ;
 wire \la_data_in_enable[95] ;
 wire \la_data_in_enable[96] ;
 wire \la_data_in_enable[97] ;
 wire \la_data_in_enable[98] ;
 wire \la_data_in_enable[99] ;
 wire \la_data_in_enable[9] ;
 wire \la_data_in_mprj_bar[0] ;
 wire \la_data_in_mprj_bar[100] ;
 wire \la_data_in_mprj_bar[101] ;
 wire \la_data_in_mprj_bar[102] ;
 wire \la_data_in_mprj_bar[103] ;
 wire \la_data_in_mprj_bar[104] ;
 wire \la_data_in_mprj_bar[105] ;
 wire \la_data_in_mprj_bar[106] ;
 wire \la_data_in_mprj_bar[107] ;
 wire \la_data_in_mprj_bar[108] ;
 wire \la_data_in_mprj_bar[109] ;
 wire \la_data_in_mprj_bar[10] ;
 wire \la_data_in_mprj_bar[110] ;
 wire \la_data_in_mprj_bar[111] ;
 wire \la_data_in_mprj_bar[112] ;
 wire \la_data_in_mprj_bar[113] ;
 wire \la_data_in_mprj_bar[114] ;
 wire \la_data_in_mprj_bar[115] ;
 wire \la_data_in_mprj_bar[116] ;
 wire \la_data_in_mprj_bar[117] ;
 wire \la_data_in_mprj_bar[118] ;
 wire \la_data_in_mprj_bar[119] ;
 wire \la_data_in_mprj_bar[11] ;
 wire \la_data_in_mprj_bar[120] ;
 wire \la_data_in_mprj_bar[121] ;
 wire \la_data_in_mprj_bar[122] ;
 wire \la_data_in_mprj_bar[123] ;
 wire \la_data_in_mprj_bar[124] ;
 wire \la_data_in_mprj_bar[125] ;
 wire \la_data_in_mprj_bar[126] ;
 wire \la_data_in_mprj_bar[127] ;
 wire \la_data_in_mprj_bar[12] ;
 wire \la_data_in_mprj_bar[13] ;
 wire \la_data_in_mprj_bar[14] ;
 wire \la_data_in_mprj_bar[15] ;
 wire \la_data_in_mprj_bar[16] ;
 wire \la_data_in_mprj_bar[17] ;
 wire \la_data_in_mprj_bar[18] ;
 wire \la_data_in_mprj_bar[19] ;
 wire \la_data_in_mprj_bar[1] ;
 wire \la_data_in_mprj_bar[20] ;
 wire \la_data_in_mprj_bar[21] ;
 wire \la_data_in_mprj_bar[22] ;
 wire \la_data_in_mprj_bar[23] ;
 wire \la_data_in_mprj_bar[24] ;
 wire \la_data_in_mprj_bar[25] ;
 wire \la_data_in_mprj_bar[26] ;
 wire \la_data_in_mprj_bar[27] ;
 wire \la_data_in_mprj_bar[28] ;
 wire \la_data_in_mprj_bar[29] ;
 wire \la_data_in_mprj_bar[2] ;
 wire \la_data_in_mprj_bar[30] ;
 wire \la_data_in_mprj_bar[31] ;
 wire \la_data_in_mprj_bar[32] ;
 wire \la_data_in_mprj_bar[33] ;
 wire \la_data_in_mprj_bar[34] ;
 wire \la_data_in_mprj_bar[35] ;
 wire \la_data_in_mprj_bar[36] ;
 wire \la_data_in_mprj_bar[37] ;
 wire \la_data_in_mprj_bar[38] ;
 wire \la_data_in_mprj_bar[39] ;
 wire \la_data_in_mprj_bar[3] ;
 wire \la_data_in_mprj_bar[40] ;
 wire \la_data_in_mprj_bar[41] ;
 wire \la_data_in_mprj_bar[42] ;
 wire \la_data_in_mprj_bar[43] ;
 wire \la_data_in_mprj_bar[44] ;
 wire \la_data_in_mprj_bar[45] ;
 wire \la_data_in_mprj_bar[46] ;
 wire \la_data_in_mprj_bar[47] ;
 wire \la_data_in_mprj_bar[48] ;
 wire \la_data_in_mprj_bar[49] ;
 wire \la_data_in_mprj_bar[4] ;
 wire \la_data_in_mprj_bar[50] ;
 wire \la_data_in_mprj_bar[51] ;
 wire \la_data_in_mprj_bar[52] ;
 wire \la_data_in_mprj_bar[53] ;
 wire \la_data_in_mprj_bar[54] ;
 wire \la_data_in_mprj_bar[55] ;
 wire \la_data_in_mprj_bar[56] ;
 wire \la_data_in_mprj_bar[57] ;
 wire \la_data_in_mprj_bar[58] ;
 wire \la_data_in_mprj_bar[59] ;
 wire \la_data_in_mprj_bar[5] ;
 wire \la_data_in_mprj_bar[60] ;
 wire \la_data_in_mprj_bar[61] ;
 wire \la_data_in_mprj_bar[62] ;
 wire \la_data_in_mprj_bar[63] ;
 wire \la_data_in_mprj_bar[64] ;
 wire \la_data_in_mprj_bar[65] ;
 wire \la_data_in_mprj_bar[66] ;
 wire \la_data_in_mprj_bar[67] ;
 wire \la_data_in_mprj_bar[68] ;
 wire \la_data_in_mprj_bar[69] ;
 wire \la_data_in_mprj_bar[6] ;
 wire \la_data_in_mprj_bar[70] ;
 wire \la_data_in_mprj_bar[71] ;
 wire \la_data_in_mprj_bar[72] ;
 wire \la_data_in_mprj_bar[73] ;
 wire \la_data_in_mprj_bar[74] ;
 wire \la_data_in_mprj_bar[75] ;
 wire \la_data_in_mprj_bar[76] ;
 wire \la_data_in_mprj_bar[77] ;
 wire \la_data_in_mprj_bar[78] ;
 wire \la_data_in_mprj_bar[79] ;
 wire \la_data_in_mprj_bar[7] ;
 wire \la_data_in_mprj_bar[80] ;
 wire \la_data_in_mprj_bar[81] ;
 wire \la_data_in_mprj_bar[82] ;
 wire \la_data_in_mprj_bar[83] ;
 wire \la_data_in_mprj_bar[84] ;
 wire \la_data_in_mprj_bar[85] ;
 wire \la_data_in_mprj_bar[86] ;
 wire \la_data_in_mprj_bar[87] ;
 wire \la_data_in_mprj_bar[88] ;
 wire \la_data_in_mprj_bar[89] ;
 wire \la_data_in_mprj_bar[8] ;
 wire \la_data_in_mprj_bar[90] ;
 wire \la_data_in_mprj_bar[91] ;
 wire \la_data_in_mprj_bar[92] ;
 wire \la_data_in_mprj_bar[93] ;
 wire \la_data_in_mprj_bar[94] ;
 wire \la_data_in_mprj_bar[95] ;
 wire \la_data_in_mprj_bar[96] ;
 wire \la_data_in_mprj_bar[97] ;
 wire \la_data_in_mprj_bar[98] ;
 wire \la_data_in_mprj_bar[99] ;
 wire \la_data_in_mprj_bar[9] ;
 wire mprj_ack_i_core_bar;
 wire \mprj_dat_i_core_bar[0] ;
 wire \mprj_dat_i_core_bar[10] ;
 wire \mprj_dat_i_core_bar[11] ;
 wire \mprj_dat_i_core_bar[12] ;
 wire \mprj_dat_i_core_bar[13] ;
 wire \mprj_dat_i_core_bar[14] ;
 wire \mprj_dat_i_core_bar[15] ;
 wire \mprj_dat_i_core_bar[16] ;
 wire \mprj_dat_i_core_bar[17] ;
 wire \mprj_dat_i_core_bar[18] ;
 wire \mprj_dat_i_core_bar[19] ;
 wire \mprj_dat_i_core_bar[1] ;
 wire \mprj_dat_i_core_bar[20] ;
 wire \mprj_dat_i_core_bar[21] ;
 wire \mprj_dat_i_core_bar[22] ;
 wire \mprj_dat_i_core_bar[23] ;
 wire \mprj_dat_i_core_bar[24] ;
 wire \mprj_dat_i_core_bar[25] ;
 wire \mprj_dat_i_core_bar[26] ;
 wire \mprj_dat_i_core_bar[27] ;
 wire \mprj_dat_i_core_bar[28] ;
 wire \mprj_dat_i_core_bar[29] ;
 wire \mprj_dat_i_core_bar[2] ;
 wire \mprj_dat_i_core_bar[30] ;
 wire \mprj_dat_i_core_bar[31] ;
 wire \mprj_dat_i_core_bar[3] ;
 wire \mprj_dat_i_core_bar[4] ;
 wire \mprj_dat_i_core_bar[5] ;
 wire \mprj_dat_i_core_bar[6] ;
 wire \mprj_dat_i_core_bar[7] ;
 wire \mprj_dat_i_core_bar[8] ;
 wire \mprj_dat_i_core_bar[9] ;
 wire \mprj_logic1[0] ;
 wire \mprj_logic1[100] ;
 wire \mprj_logic1[101] ;
 wire \mprj_logic1[102] ;
 wire \mprj_logic1[103] ;
 wire \mprj_logic1[104] ;
 wire \mprj_logic1[105] ;
 wire \mprj_logic1[106] ;
 wire \mprj_logic1[107] ;
 wire \mprj_logic1[108] ;
 wire \mprj_logic1[109] ;
 wire \mprj_logic1[10] ;
 wire \mprj_logic1[110] ;
 wire \mprj_logic1[111] ;
 wire \mprj_logic1[112] ;
 wire \mprj_logic1[113] ;
 wire \mprj_logic1[114] ;
 wire \mprj_logic1[115] ;
 wire \mprj_logic1[116] ;
 wire \mprj_logic1[117] ;
 wire \mprj_logic1[118] ;
 wire \mprj_logic1[119] ;
 wire \mprj_logic1[11] ;
 wire \mprj_logic1[120] ;
 wire \mprj_logic1[121] ;
 wire \mprj_logic1[122] ;
 wire \mprj_logic1[123] ;
 wire \mprj_logic1[124] ;
 wire \mprj_logic1[125] ;
 wire \mprj_logic1[126] ;
 wire \mprj_logic1[127] ;
 wire \mprj_logic1[128] ;
 wire \mprj_logic1[129] ;
 wire \mprj_logic1[12] ;
 wire \mprj_logic1[130] ;
 wire \mprj_logic1[131] ;
 wire \mprj_logic1[132] ;
 wire \mprj_logic1[133] ;
 wire \mprj_logic1[134] ;
 wire \mprj_logic1[135] ;
 wire \mprj_logic1[136] ;
 wire \mprj_logic1[137] ;
 wire \mprj_logic1[138] ;
 wire \mprj_logic1[139] ;
 wire \mprj_logic1[13] ;
 wire \mprj_logic1[140] ;
 wire \mprj_logic1[141] ;
 wire \mprj_logic1[142] ;
 wire \mprj_logic1[143] ;
 wire \mprj_logic1[144] ;
 wire \mprj_logic1[145] ;
 wire \mprj_logic1[146] ;
 wire \mprj_logic1[147] ;
 wire \mprj_logic1[148] ;
 wire \mprj_logic1[149] ;
 wire \mprj_logic1[14] ;
 wire \mprj_logic1[150] ;
 wire \mprj_logic1[151] ;
 wire \mprj_logic1[152] ;
 wire \mprj_logic1[153] ;
 wire \mprj_logic1[154] ;
 wire \mprj_logic1[155] ;
 wire \mprj_logic1[156] ;
 wire \mprj_logic1[157] ;
 wire \mprj_logic1[158] ;
 wire \mprj_logic1[159] ;
 wire \mprj_logic1[15] ;
 wire \mprj_logic1[160] ;
 wire \mprj_logic1[161] ;
 wire \mprj_logic1[162] ;
 wire \mprj_logic1[163] ;
 wire \mprj_logic1[164] ;
 wire \mprj_logic1[165] ;
 wire \mprj_logic1[166] ;
 wire \mprj_logic1[167] ;
 wire \mprj_logic1[168] ;
 wire \mprj_logic1[169] ;
 wire \mprj_logic1[16] ;
 wire \mprj_logic1[170] ;
 wire \mprj_logic1[171] ;
 wire \mprj_logic1[172] ;
 wire \mprj_logic1[173] ;
 wire \mprj_logic1[174] ;
 wire \mprj_logic1[175] ;
 wire \mprj_logic1[176] ;
 wire \mprj_logic1[177] ;
 wire \mprj_logic1[178] ;
 wire \mprj_logic1[179] ;
 wire \mprj_logic1[17] ;
 wire \mprj_logic1[180] ;
 wire \mprj_logic1[181] ;
 wire \mprj_logic1[182] ;
 wire \mprj_logic1[183] ;
 wire \mprj_logic1[184] ;
 wire \mprj_logic1[185] ;
 wire \mprj_logic1[186] ;
 wire \mprj_logic1[187] ;
 wire \mprj_logic1[188] ;
 wire \mprj_logic1[189] ;
 wire \mprj_logic1[18] ;
 wire \mprj_logic1[190] ;
 wire \mprj_logic1[191] ;
 wire \mprj_logic1[192] ;
 wire \mprj_logic1[193] ;
 wire \mprj_logic1[194] ;
 wire \mprj_logic1[195] ;
 wire \mprj_logic1[196] ;
 wire \mprj_logic1[197] ;
 wire \mprj_logic1[198] ;
 wire \mprj_logic1[199] ;
 wire \mprj_logic1[19] ;
 wire \mprj_logic1[1] ;
 wire \mprj_logic1[200] ;
 wire \mprj_logic1[201] ;
 wire \mprj_logic1[202] ;
 wire \mprj_logic1[203] ;
 wire \mprj_logic1[204] ;
 wire \mprj_logic1[205] ;
 wire \mprj_logic1[206] ;
 wire \mprj_logic1[207] ;
 wire \mprj_logic1[208] ;
 wire \mprj_logic1[209] ;
 wire \mprj_logic1[20] ;
 wire \mprj_logic1[210] ;
 wire \mprj_logic1[211] ;
 wire \mprj_logic1[212] ;
 wire \mprj_logic1[213] ;
 wire \mprj_logic1[214] ;
 wire \mprj_logic1[215] ;
 wire \mprj_logic1[216] ;
 wire \mprj_logic1[217] ;
 wire \mprj_logic1[218] ;
 wire \mprj_logic1[219] ;
 wire \mprj_logic1[21] ;
 wire \mprj_logic1[220] ;
 wire \mprj_logic1[221] ;
 wire \mprj_logic1[222] ;
 wire \mprj_logic1[223] ;
 wire \mprj_logic1[224] ;
 wire \mprj_logic1[225] ;
 wire \mprj_logic1[226] ;
 wire \mprj_logic1[227] ;
 wire \mprj_logic1[228] ;
 wire \mprj_logic1[229] ;
 wire \mprj_logic1[22] ;
 wire \mprj_logic1[230] ;
 wire \mprj_logic1[231] ;
 wire \mprj_logic1[232] ;
 wire \mprj_logic1[233] ;
 wire \mprj_logic1[234] ;
 wire \mprj_logic1[235] ;
 wire \mprj_logic1[236] ;
 wire \mprj_logic1[237] ;
 wire \mprj_logic1[238] ;
 wire \mprj_logic1[239] ;
 wire \mprj_logic1[23] ;
 wire \mprj_logic1[240] ;
 wire \mprj_logic1[241] ;
 wire \mprj_logic1[242] ;
 wire \mprj_logic1[243] ;
 wire \mprj_logic1[244] ;
 wire \mprj_logic1[245] ;
 wire \mprj_logic1[246] ;
 wire \mprj_logic1[247] ;
 wire \mprj_logic1[248] ;
 wire \mprj_logic1[249] ;
 wire \mprj_logic1[24] ;
 wire \mprj_logic1[250] ;
 wire \mprj_logic1[251] ;
 wire \mprj_logic1[252] ;
 wire \mprj_logic1[253] ;
 wire \mprj_logic1[254] ;
 wire \mprj_logic1[255] ;
 wire \mprj_logic1[256] ;
 wire \mprj_logic1[257] ;
 wire \mprj_logic1[258] ;
 wire \mprj_logic1[259] ;
 wire \mprj_logic1[25] ;
 wire \mprj_logic1[260] ;
 wire \mprj_logic1[261] ;
 wire \mprj_logic1[262] ;
 wire \mprj_logic1[263] ;
 wire \mprj_logic1[264] ;
 wire \mprj_logic1[265] ;
 wire \mprj_logic1[266] ;
 wire \mprj_logic1[267] ;
 wire \mprj_logic1[268] ;
 wire \mprj_logic1[269] ;
 wire \mprj_logic1[26] ;
 wire \mprj_logic1[270] ;
 wire \mprj_logic1[271] ;
 wire \mprj_logic1[272] ;
 wire \mprj_logic1[273] ;
 wire \mprj_logic1[274] ;
 wire \mprj_logic1[275] ;
 wire \mprj_logic1[276] ;
 wire \mprj_logic1[277] ;
 wire \mprj_logic1[278] ;
 wire \mprj_logic1[279] ;
 wire \mprj_logic1[27] ;
 wire \mprj_logic1[280] ;
 wire \mprj_logic1[281] ;
 wire \mprj_logic1[282] ;
 wire \mprj_logic1[283] ;
 wire \mprj_logic1[284] ;
 wire \mprj_logic1[285] ;
 wire \mprj_logic1[286] ;
 wire \mprj_logic1[287] ;
 wire \mprj_logic1[288] ;
 wire \mprj_logic1[289] ;
 wire \mprj_logic1[28] ;
 wire \mprj_logic1[290] ;
 wire \mprj_logic1[291] ;
 wire \mprj_logic1[292] ;
 wire \mprj_logic1[293] ;
 wire \mprj_logic1[294] ;
 wire \mprj_logic1[295] ;
 wire \mprj_logic1[296] ;
 wire \mprj_logic1[297] ;
 wire \mprj_logic1[298] ;
 wire \mprj_logic1[299] ;
 wire \mprj_logic1[29] ;
 wire \mprj_logic1[2] ;
 wire \mprj_logic1[300] ;
 wire \mprj_logic1[301] ;
 wire \mprj_logic1[302] ;
 wire \mprj_logic1[303] ;
 wire \mprj_logic1[304] ;
 wire \mprj_logic1[305] ;
 wire \mprj_logic1[306] ;
 wire \mprj_logic1[307] ;
 wire \mprj_logic1[308] ;
 wire \mprj_logic1[309] ;
 wire \mprj_logic1[30] ;
 wire \mprj_logic1[310] ;
 wire \mprj_logic1[311] ;
 wire \mprj_logic1[312] ;
 wire \mprj_logic1[313] ;
 wire \mprj_logic1[314] ;
 wire \mprj_logic1[315] ;
 wire \mprj_logic1[316] ;
 wire \mprj_logic1[317] ;
 wire \mprj_logic1[318] ;
 wire \mprj_logic1[319] ;
 wire \mprj_logic1[31] ;
 wire \mprj_logic1[320] ;
 wire \mprj_logic1[321] ;
 wire \mprj_logic1[322] ;
 wire \mprj_logic1[323] ;
 wire \mprj_logic1[324] ;
 wire \mprj_logic1[325] ;
 wire \mprj_logic1[326] ;
 wire \mprj_logic1[327] ;
 wire \mprj_logic1[328] ;
 wire \mprj_logic1[329] ;
 wire \mprj_logic1[32] ;
 wire \mprj_logic1[330] ;
 wire \mprj_logic1[331] ;
 wire \mprj_logic1[332] ;
 wire \mprj_logic1[333] ;
 wire \mprj_logic1[334] ;
 wire \mprj_logic1[335] ;
 wire \mprj_logic1[336] ;
 wire \mprj_logic1[337] ;
 wire \mprj_logic1[338] ;
 wire \mprj_logic1[339] ;
 wire \mprj_logic1[33] ;
 wire \mprj_logic1[340] ;
 wire \mprj_logic1[341] ;
 wire \mprj_logic1[342] ;
 wire \mprj_logic1[343] ;
 wire \mprj_logic1[344] ;
 wire \mprj_logic1[345] ;
 wire \mprj_logic1[346] ;
 wire \mprj_logic1[347] ;
 wire \mprj_logic1[348] ;
 wire \mprj_logic1[349] ;
 wire \mprj_logic1[34] ;
 wire \mprj_logic1[350] ;
 wire \mprj_logic1[351] ;
 wire \mprj_logic1[352] ;
 wire \mprj_logic1[353] ;
 wire \mprj_logic1[354] ;
 wire \mprj_logic1[355] ;
 wire \mprj_logic1[356] ;
 wire \mprj_logic1[357] ;
 wire \mprj_logic1[358] ;
 wire \mprj_logic1[359] ;
 wire \mprj_logic1[35] ;
 wire \mprj_logic1[360] ;
 wire \mprj_logic1[361] ;
 wire \mprj_logic1[362] ;
 wire \mprj_logic1[363] ;
 wire \mprj_logic1[364] ;
 wire \mprj_logic1[365] ;
 wire \mprj_logic1[366] ;
 wire \mprj_logic1[367] ;
 wire \mprj_logic1[368] ;
 wire \mprj_logic1[369] ;
 wire \mprj_logic1[36] ;
 wire \mprj_logic1[370] ;
 wire \mprj_logic1[371] ;
 wire \mprj_logic1[372] ;
 wire \mprj_logic1[373] ;
 wire \mprj_logic1[374] ;
 wire \mprj_logic1[375] ;
 wire \mprj_logic1[376] ;
 wire \mprj_logic1[377] ;
 wire \mprj_logic1[378] ;
 wire \mprj_logic1[379] ;
 wire \mprj_logic1[37] ;
 wire \mprj_logic1[380] ;
 wire \mprj_logic1[381] ;
 wire \mprj_logic1[382] ;
 wire \mprj_logic1[383] ;
 wire \mprj_logic1[384] ;
 wire \mprj_logic1[385] ;
 wire \mprj_logic1[386] ;
 wire \mprj_logic1[387] ;
 wire \mprj_logic1[388] ;
 wire \mprj_logic1[389] ;
 wire \mprj_logic1[38] ;
 wire \mprj_logic1[390] ;
 wire \mprj_logic1[391] ;
 wire \mprj_logic1[392] ;
 wire \mprj_logic1[393] ;
 wire \mprj_logic1[394] ;
 wire \mprj_logic1[395] ;
 wire \mprj_logic1[396] ;
 wire \mprj_logic1[397] ;
 wire \mprj_logic1[398] ;
 wire \mprj_logic1[399] ;
 wire \mprj_logic1[39] ;
 wire \mprj_logic1[3] ;
 wire \mprj_logic1[400] ;
 wire \mprj_logic1[401] ;
 wire \mprj_logic1[402] ;
 wire \mprj_logic1[403] ;
 wire \mprj_logic1[404] ;
 wire \mprj_logic1[405] ;
 wire \mprj_logic1[406] ;
 wire \mprj_logic1[407] ;
 wire \mprj_logic1[408] ;
 wire \mprj_logic1[409] ;
 wire \mprj_logic1[40] ;
 wire \mprj_logic1[410] ;
 wire \mprj_logic1[411] ;
 wire \mprj_logic1[412] ;
 wire \mprj_logic1[413] ;
 wire \mprj_logic1[414] ;
 wire \mprj_logic1[415] ;
 wire \mprj_logic1[416] ;
 wire \mprj_logic1[417] ;
 wire \mprj_logic1[418] ;
 wire \mprj_logic1[419] ;
 wire \mprj_logic1[41] ;
 wire \mprj_logic1[420] ;
 wire \mprj_logic1[421] ;
 wire \mprj_logic1[422] ;
 wire \mprj_logic1[423] ;
 wire \mprj_logic1[424] ;
 wire \mprj_logic1[425] ;
 wire \mprj_logic1[426] ;
 wire \mprj_logic1[427] ;
 wire \mprj_logic1[428] ;
 wire \mprj_logic1[429] ;
 wire \mprj_logic1[42] ;
 wire \mprj_logic1[430] ;
 wire \mprj_logic1[431] ;
 wire \mprj_logic1[432] ;
 wire \mprj_logic1[433] ;
 wire \mprj_logic1[434] ;
 wire \mprj_logic1[435] ;
 wire \mprj_logic1[436] ;
 wire \mprj_logic1[437] ;
 wire \mprj_logic1[438] ;
 wire \mprj_logic1[439] ;
 wire \mprj_logic1[43] ;
 wire \mprj_logic1[440] ;
 wire \mprj_logic1[441] ;
 wire \mprj_logic1[442] ;
 wire \mprj_logic1[443] ;
 wire \mprj_logic1[444] ;
 wire \mprj_logic1[445] ;
 wire \mprj_logic1[446] ;
 wire \mprj_logic1[447] ;
 wire \mprj_logic1[448] ;
 wire \mprj_logic1[449] ;
 wire \mprj_logic1[44] ;
 wire \mprj_logic1[450] ;
 wire \mprj_logic1[451] ;
 wire \mprj_logic1[452] ;
 wire \mprj_logic1[453] ;
 wire \mprj_logic1[454] ;
 wire \mprj_logic1[455] ;
 wire \mprj_logic1[456] ;
 wire \mprj_logic1[457] ;
 wire \mprj_logic1[458] ;
 wire \mprj_logic1[459] ;
 wire \mprj_logic1[45] ;
 wire \mprj_logic1[460] ;
 wire \mprj_logic1[462] ;
 wire \mprj_logic1[46] ;
 wire \mprj_logic1[47] ;
 wire \mprj_logic1[48] ;
 wire \mprj_logic1[49] ;
 wire \mprj_logic1[4] ;
 wire \mprj_logic1[50] ;
 wire \mprj_logic1[51] ;
 wire \mprj_logic1[52] ;
 wire \mprj_logic1[53] ;
 wire \mprj_logic1[54] ;
 wire \mprj_logic1[55] ;
 wire \mprj_logic1[56] ;
 wire \mprj_logic1[57] ;
 wire \mprj_logic1[58] ;
 wire \mprj_logic1[59] ;
 wire \mprj_logic1[5] ;
 wire \mprj_logic1[60] ;
 wire \mprj_logic1[61] ;
 wire \mprj_logic1[62] ;
 wire \mprj_logic1[63] ;
 wire \mprj_logic1[64] ;
 wire \mprj_logic1[65] ;
 wire \mprj_logic1[66] ;
 wire \mprj_logic1[67] ;
 wire \mprj_logic1[68] ;
 wire \mprj_logic1[69] ;
 wire \mprj_logic1[6] ;
 wire \mprj_logic1[70] ;
 wire \mprj_logic1[71] ;
 wire \mprj_logic1[72] ;
 wire \mprj_logic1[73] ;
 wire \mprj_logic1[74] ;
 wire \mprj_logic1[75] ;
 wire \mprj_logic1[76] ;
 wire \mprj_logic1[77] ;
 wire \mprj_logic1[78] ;
 wire \mprj_logic1[79] ;
 wire \mprj_logic1[7] ;
 wire \mprj_logic1[80] ;
 wire \mprj_logic1[81] ;
 wire \mprj_logic1[82] ;
 wire \mprj_logic1[83] ;
 wire \mprj_logic1[84] ;
 wire \mprj_logic1[85] ;
 wire \mprj_logic1[86] ;
 wire \mprj_logic1[87] ;
 wire \mprj_logic1[88] ;
 wire \mprj_logic1[89] ;
 wire \mprj_logic1[8] ;
 wire \mprj_logic1[90] ;
 wire \mprj_logic1[91] ;
 wire \mprj_logic1[92] ;
 wire \mprj_logic1[93] ;
 wire \mprj_logic1[94] ;
 wire \mprj_logic1[95] ;
 wire \mprj_logic1[96] ;
 wire \mprj_logic1[97] ;
 wire \mprj_logic1[98] ;
 wire \mprj_logic1[99] ;
 wire \mprj_logic1[9] ;
 wire \user_irq_bar[0] ;
 wire \user_irq_bar[1] ;
 wire \user_irq_bar[2] ;
 wire \user_irq_enable[0] ;
 wire \user_irq_enable[1] ;
 wire \user_irq_enable[2] ;
 wire wb_in_enable;
 wire net2;
 wire net1;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;

 sky130_fd_sc_hd__clkinv_2 _000_ (.A(\la_data_in_mprj_bar[17] ),
    .Y(net627));
 sky130_fd_sc_hd__clkinv_2 _001_ (.A(\la_data_in_mprj_bar[18] ),
    .Y(net628));
 sky130_fd_sc_hd__inv_2 _002_ (.A(\la_data_in_mprj_bar[19] ),
    .Y(net629));
 sky130_fd_sc_hd__inv_2 _003_ (.A(\la_data_in_mprj_bar[20] ),
    .Y(net631));
 sky130_fd_sc_hd__inv_2 _004_ (.A(\la_data_in_mprj_bar[21] ),
    .Y(net632));
 sky130_fd_sc_hd__inv_2 _005_ (.A(\la_data_in_mprj_bar[22] ),
    .Y(net633));
 sky130_fd_sc_hd__inv_2 _006_ (.A(\la_data_in_mprj_bar[23] ),
    .Y(net634));
 sky130_fd_sc_hd__inv_2 _007_ (.A(\la_data_in_mprj_bar[24] ),
    .Y(net635));
 sky130_fd_sc_hd__inv_2 _008_ (.A(\la_data_in_mprj_bar[25] ),
    .Y(net636));
 sky130_fd_sc_hd__inv_2 _009_ (.A(\la_data_in_mprj_bar[26] ),
    .Y(net637));
 sky130_fd_sc_hd__inv_2 _010_ (.A(\la_data_in_mprj_bar[27] ),
    .Y(net638));
 sky130_fd_sc_hd__inv_2 _011_ (.A(\la_data_in_mprj_bar[28] ),
    .Y(net639));
 sky130_fd_sc_hd__inv_2 _012_ (.A(\la_data_in_mprj_bar[29] ),
    .Y(net640));
 sky130_fd_sc_hd__inv_2 _013_ (.A(\la_data_in_mprj_bar[30] ),
    .Y(net642));
 sky130_fd_sc_hd__clkinv_2 _014_ (.A(\la_data_in_mprj_bar[31] ),
    .Y(net643));
 sky130_fd_sc_hd__inv_2 _015_ (.A(\la_data_in_mprj_bar[32] ),
    .Y(net644));
 sky130_fd_sc_hd__inv_2 _016_ (.A(\la_data_in_mprj_bar[33] ),
    .Y(net645));
 sky130_fd_sc_hd__clkinv_2 _017_ (.A(\la_data_in_mprj_bar[34] ),
    .Y(net646));
 sky130_fd_sc_hd__clkinv_2 _018_ (.A(\la_data_in_mprj_bar[35] ),
    .Y(net647));
 sky130_fd_sc_hd__clkinv_2 _019_ (.A(\la_data_in_mprj_bar[36] ),
    .Y(net648));
 sky130_fd_sc_hd__inv_2 _020_ (.A(\la_data_in_mprj_bar[37] ),
    .Y(net649));
 sky130_fd_sc_hd__inv_2 _021_ (.A(\la_data_in_mprj_bar[38] ),
    .Y(net650));
 sky130_fd_sc_hd__inv_2 _022_ (.A(\la_data_in_mprj_bar[39] ),
    .Y(net651));
 sky130_fd_sc_hd__inv_2 _023_ (.A(\la_data_in_mprj_bar[40] ),
    .Y(net653));
 sky130_fd_sc_hd__inv_2 _024_ (.A(\la_data_in_mprj_bar[41] ),
    .Y(net654));
 sky130_fd_sc_hd__inv_2 _025_ (.A(\la_data_in_mprj_bar[42] ),
    .Y(net655));
 sky130_fd_sc_hd__inv_2 _026_ (.A(\la_data_in_mprj_bar[43] ),
    .Y(net656));
 sky130_fd_sc_hd__inv_2 _027_ (.A(\la_data_in_mprj_bar[44] ),
    .Y(net657));
 sky130_fd_sc_hd__inv_2 _028_ (.A(\la_data_in_mprj_bar[45] ),
    .Y(net658));
 sky130_fd_sc_hd__inv_2 _029_ (.A(\la_data_in_mprj_bar[46] ),
    .Y(net659));
 sky130_fd_sc_hd__inv_2 _030_ (.A(\la_data_in_mprj_bar[47] ),
    .Y(net660));
 sky130_fd_sc_hd__inv_2 _031_ (.A(\la_data_in_mprj_bar[48] ),
    .Y(net661));
 sky130_fd_sc_hd__clkinv_2 _032_ (.A(\la_data_in_mprj_bar[49] ),
    .Y(net662));
 sky130_fd_sc_hd__clkinv_2 _033_ (.A(\la_data_in_mprj_bar[50] ),
    .Y(net664));
 sky130_fd_sc_hd__clkinv_2 _034_ (.A(\la_data_in_mprj_bar[51] ),
    .Y(net665));
 sky130_fd_sc_hd__inv_2 _035_ (.A(\la_data_in_mprj_bar[52] ),
    .Y(net666));
 sky130_fd_sc_hd__inv_2 _036_ (.A(\la_data_in_mprj_bar[53] ),
    .Y(net667));
 sky130_fd_sc_hd__inv_2 _037_ (.A(\la_data_in_mprj_bar[54] ),
    .Y(net668));
 sky130_fd_sc_hd__inv_2 _038_ (.A(\la_data_in_mprj_bar[55] ),
    .Y(net669));
 sky130_fd_sc_hd__inv_2 _039_ (.A(\la_data_in_mprj_bar[56] ),
    .Y(net670));
 sky130_fd_sc_hd__inv_2 _040_ (.A(\la_data_in_mprj_bar[57] ),
    .Y(net671));
 sky130_fd_sc_hd__inv_2 _041_ (.A(\la_data_in_mprj_bar[58] ),
    .Y(net672));
 sky130_fd_sc_hd__inv_2 _042_ (.A(\la_data_in_mprj_bar[59] ),
    .Y(net673));
 sky130_fd_sc_hd__inv_2 _043_ (.A(\la_data_in_mprj_bar[60] ),
    .Y(net675));
 sky130_fd_sc_hd__clkinv_2 _044_ (.A(\la_data_in_mprj_bar[61] ),
    .Y(net676));
 sky130_fd_sc_hd__clkinv_2 _045_ (.A(\la_data_in_mprj_bar[62] ),
    .Y(net677));
 sky130_fd_sc_hd__clkinv_2 _046_ (.A(\la_data_in_mprj_bar[63] ),
    .Y(net678));
 sky130_fd_sc_hd__clkinv_2 _047_ (.A(\la_data_in_mprj_bar[64] ),
    .Y(net679));
 sky130_fd_sc_hd__inv_2 _048_ (.A(\la_data_in_mprj_bar[65] ),
    .Y(net680));
 sky130_fd_sc_hd__clkinv_4 _049_ (.A(\la_data_in_mprj_bar[66] ),
    .Y(net681));
 sky130_fd_sc_hd__clkinv_4 _050_ (.A(\la_data_in_mprj_bar[67] ),
    .Y(net682));
 sky130_fd_sc_hd__inv_4 _051_ (.A(\la_data_in_mprj_bar[68] ),
    .Y(net683));
 sky130_fd_sc_hd__clkinv_4 _052_ (.A(\la_data_in_mprj_bar[69] ),
    .Y(net684));
 sky130_fd_sc_hd__clkinv_4 _053_ (.A(\la_data_in_mprj_bar[70] ),
    .Y(net686));
 sky130_fd_sc_hd__clkinv_4 _054_ (.A(\la_data_in_mprj_bar[71] ),
    .Y(net687));
 sky130_fd_sc_hd__clkinv_4 _055_ (.A(\la_data_in_mprj_bar[72] ),
    .Y(net688));
 sky130_fd_sc_hd__clkinv_4 _056_ (.A(\la_data_in_mprj_bar[73] ),
    .Y(net689));
 sky130_fd_sc_hd__inv_2 _057_ (.A(\la_data_in_mprj_bar[74] ),
    .Y(net690));
 sky130_fd_sc_hd__inv_2 _058_ (.A(\la_data_in_mprj_bar[75] ),
    .Y(net691));
 sky130_fd_sc_hd__inv_2 _059_ (.A(\la_data_in_mprj_bar[76] ),
    .Y(net692));
 sky130_fd_sc_hd__inv_2 _060_ (.A(\la_data_in_mprj_bar[77] ),
    .Y(net693));
 sky130_fd_sc_hd__clkinv_2 _061_ (.A(\la_data_in_mprj_bar[78] ),
    .Y(net694));
 sky130_fd_sc_hd__inv_2 _062_ (.A(\la_data_in_mprj_bar[79] ),
    .Y(net695));
 sky130_fd_sc_hd__inv_2 _063_ (.A(\la_data_in_mprj_bar[80] ),
    .Y(net697));
 sky130_fd_sc_hd__clkinv_2 _064_ (.A(\la_data_in_mprj_bar[81] ),
    .Y(net698));
 sky130_fd_sc_hd__clkinv_2 _065_ (.A(\la_data_in_mprj_bar[82] ),
    .Y(net699));
 sky130_fd_sc_hd__clkinv_2 _066_ (.A(\la_data_in_mprj_bar[83] ),
    .Y(net700));
 sky130_fd_sc_hd__clkinv_2 _067_ (.A(\la_data_in_mprj_bar[84] ),
    .Y(net701));
 sky130_fd_sc_hd__clkinv_2 _068_ (.A(\la_data_in_mprj_bar[85] ),
    .Y(net702));
 sky130_fd_sc_hd__clkinv_2 _069_ (.A(\la_data_in_mprj_bar[86] ),
    .Y(net703));
 sky130_fd_sc_hd__clkinv_2 _070_ (.A(\la_data_in_mprj_bar[87] ),
    .Y(net704));
 sky130_fd_sc_hd__inv_2 _071_ (.A(\la_data_in_mprj_bar[88] ),
    .Y(net705));
 sky130_fd_sc_hd__clkinv_2 _072_ (.A(\la_data_in_mprj_bar[89] ),
    .Y(net706));
 sky130_fd_sc_hd__clkinv_2 _073_ (.A(\la_data_in_mprj_bar[90] ),
    .Y(net708));
 sky130_fd_sc_hd__inv_2 _074_ (.A(\la_data_in_mprj_bar[91] ),
    .Y(net709));
 sky130_fd_sc_hd__clkinv_2 _075_ (.A(\la_data_in_mprj_bar[92] ),
    .Y(net710));
 sky130_fd_sc_hd__inv_2 _076_ (.A(\la_data_in_mprj_bar[93] ),
    .Y(net711));
 sky130_fd_sc_hd__clkinv_4 _077_ (.A(\la_data_in_mprj_bar[94] ),
    .Y(net712));
 sky130_fd_sc_hd__clkinv_4 _078_ (.A(\la_data_in_mprj_bar[95] ),
    .Y(net713));
 sky130_fd_sc_hd__clkinv_4 _079_ (.A(\la_data_in_mprj_bar[96] ),
    .Y(net714));
 sky130_fd_sc_hd__inv_2 _080_ (.A(\la_data_in_mprj_bar[97] ),
    .Y(net715));
 sky130_fd_sc_hd__inv_2 _081_ (.A(\la_data_in_mprj_bar[98] ),
    .Y(net716));
 sky130_fd_sc_hd__inv_2 _082_ (.A(\la_data_in_mprj_bar[99] ),
    .Y(net717));
 sky130_fd_sc_hd__clkinv_2 _083_ (.A(\la_data_in_mprj_bar[100] ),
    .Y(net592));
 sky130_fd_sc_hd__clkinv_2 _084_ (.A(\la_data_in_mprj_bar[101] ),
    .Y(net593));
 sky130_fd_sc_hd__clkinv_2 _085_ (.A(\la_data_in_mprj_bar[102] ),
    .Y(net594));
 sky130_fd_sc_hd__inv_2 _086_ (.A(\la_data_in_mprj_bar[103] ),
    .Y(net595));
 sky130_fd_sc_hd__inv_2 _087_ (.A(\la_data_in_mprj_bar[104] ),
    .Y(net596));
 sky130_fd_sc_hd__inv_2 _088_ (.A(\la_data_in_mprj_bar[105] ),
    .Y(net597));
 sky130_fd_sc_hd__inv_2 _089_ (.A(\la_data_in_mprj_bar[106] ),
    .Y(net598));
 sky130_fd_sc_hd__inv_2 _090_ (.A(\la_data_in_mprj_bar[107] ),
    .Y(net599));
 sky130_fd_sc_hd__clkinv_2 _091_ (.A(\la_data_in_mprj_bar[108] ),
    .Y(net600));
 sky130_fd_sc_hd__clkinv_2 _092_ (.A(\la_data_in_mprj_bar[109] ),
    .Y(net601));
 sky130_fd_sc_hd__inv_2 _093_ (.A(\la_data_in_mprj_bar[110] ),
    .Y(net603));
 sky130_fd_sc_hd__inv_2 _094_ (.A(\la_data_in_mprj_bar[111] ),
    .Y(net604));
 sky130_fd_sc_hd__inv_2 _095_ (.A(\la_data_in_mprj_bar[112] ),
    .Y(net605));
 sky130_fd_sc_hd__inv_2 _096_ (.A(\la_data_in_mprj_bar[113] ),
    .Y(net606));
 sky130_fd_sc_hd__inv_2 _097_ (.A(\la_data_in_mprj_bar[114] ),
    .Y(net607));
 sky130_fd_sc_hd__inv_2 _098_ (.A(\la_data_in_mprj_bar[115] ),
    .Y(net608));
 sky130_fd_sc_hd__inv_2 _099_ (.A(\la_data_in_mprj_bar[116] ),
    .Y(net609));
 sky130_fd_sc_hd__inv_2 _100_ (.A(\la_data_in_mprj_bar[117] ),
    .Y(net610));
 sky130_fd_sc_hd__inv_2 _101_ (.A(\la_data_in_mprj_bar[118] ),
    .Y(net611));
 sky130_fd_sc_hd__clkinv_2 _102_ (.A(\la_data_in_mprj_bar[119] ),
    .Y(net612));
 sky130_fd_sc_hd__clkinv_2 _103_ (.A(\la_data_in_mprj_bar[120] ),
    .Y(net614));
 sky130_fd_sc_hd__clkinv_2 _104_ (.A(\la_data_in_mprj_bar[121] ),
    .Y(net615));
 sky130_fd_sc_hd__clkinv_2 _105_ (.A(\la_data_in_mprj_bar[122] ),
    .Y(net616));
 sky130_fd_sc_hd__inv_2 _106_ (.A(\la_data_in_mprj_bar[123] ),
    .Y(net617));
 sky130_fd_sc_hd__inv_2 _107_ (.A(\la_data_in_mprj_bar[124] ),
    .Y(net618));
 sky130_fd_sc_hd__clkinv_2 _108_ (.A(\la_data_in_mprj_bar[125] ),
    .Y(net619));
 sky130_fd_sc_hd__clkinv_2 _109_ (.A(\la_data_in_mprj_bar[126] ),
    .Y(net620));
 sky130_fd_sc_hd__inv_2 _110_ (.A(\la_data_in_mprj_bar[127] ),
    .Y(net621));
 sky130_fd_sc_hd__clkinv_2 _111_ (.A(\user_irq_bar[0] ),
    .Y(net957));
 sky130_fd_sc_hd__inv_2 _112_ (.A(\user_irq_bar[1] ),
    .Y(net958));
 sky130_fd_sc_hd__inv_2 _113_ (.A(\user_irq_bar[2] ),
    .Y(net959));
 sky130_fd_sc_hd__inv_2 _114_ (.A(\mprj_dat_i_core_bar[0] ),
    .Y(net881));
 sky130_fd_sc_hd__inv_2 _115_ (.A(\mprj_dat_i_core_bar[1] ),
    .Y(net892));
 sky130_fd_sc_hd__inv_2 _116_ (.A(\mprj_dat_i_core_bar[2] ),
    .Y(net903));
 sky130_fd_sc_hd__inv_2 _117_ (.A(\mprj_dat_i_core_bar[3] ),
    .Y(net906));
 sky130_fd_sc_hd__inv_2 _118_ (.A(\mprj_dat_i_core_bar[4] ),
    .Y(net907));
 sky130_fd_sc_hd__inv_2 _119_ (.A(\mprj_dat_i_core_bar[5] ),
    .Y(net908));
 sky130_fd_sc_hd__inv_2 _120_ (.A(\mprj_dat_i_core_bar[6] ),
    .Y(net909));
 sky130_fd_sc_hd__inv_2 _121_ (.A(\mprj_dat_i_core_bar[7] ),
    .Y(net910));
 sky130_fd_sc_hd__inv_2 _122_ (.A(\mprj_dat_i_core_bar[8] ),
    .Y(net911));
 sky130_fd_sc_hd__clkinv_2 _123_ (.A(\mprj_dat_i_core_bar[9] ),
    .Y(net912));
 sky130_fd_sc_hd__inv_2 _124_ (.A(\mprj_dat_i_core_bar[10] ),
    .Y(net882));
 sky130_fd_sc_hd__inv_2 _125_ (.A(\mprj_dat_i_core_bar[11] ),
    .Y(net883));
 sky130_fd_sc_hd__inv_2 _126_ (.A(\mprj_dat_i_core_bar[12] ),
    .Y(net884));
 sky130_fd_sc_hd__inv_2 _127_ (.A(\mprj_dat_i_core_bar[13] ),
    .Y(net885));
 sky130_fd_sc_hd__inv_2 _128_ (.A(\mprj_dat_i_core_bar[14] ),
    .Y(net886));
 sky130_fd_sc_hd__inv_2 _129_ (.A(\mprj_dat_i_core_bar[15] ),
    .Y(net887));
 sky130_fd_sc_hd__inv_2 _130_ (.A(\mprj_dat_i_core_bar[16] ),
    .Y(net888));
 sky130_fd_sc_hd__inv_2 _131_ (.A(\mprj_dat_i_core_bar[17] ),
    .Y(net889));
 sky130_fd_sc_hd__inv_2 _132_ (.A(\mprj_dat_i_core_bar[18] ),
    .Y(net890));
 sky130_fd_sc_hd__inv_2 _133_ (.A(\mprj_dat_i_core_bar[19] ),
    .Y(net891));
 sky130_fd_sc_hd__inv_2 _134_ (.A(\mprj_dat_i_core_bar[20] ),
    .Y(net893));
 sky130_fd_sc_hd__inv_2 _135_ (.A(\mprj_dat_i_core_bar[21] ),
    .Y(net894));
 sky130_fd_sc_hd__clkinv_2 _136_ (.A(\mprj_dat_i_core_bar[22] ),
    .Y(net895));
 sky130_fd_sc_hd__clkinv_2 _137_ (.A(\mprj_dat_i_core_bar[23] ),
    .Y(net896));
 sky130_fd_sc_hd__clkinv_2 _138_ (.A(\mprj_dat_i_core_bar[24] ),
    .Y(net897));
 sky130_fd_sc_hd__clkinv_2 _139_ (.A(\mprj_dat_i_core_bar[25] ),
    .Y(net898));
 sky130_fd_sc_hd__clkinv_2 _140_ (.A(\mprj_dat_i_core_bar[26] ),
    .Y(net899));
 sky130_fd_sc_hd__clkinv_2 _141_ (.A(\mprj_dat_i_core_bar[27] ),
    .Y(net900));
 sky130_fd_sc_hd__clkinv_2 _142_ (.A(\mprj_dat_i_core_bar[28] ),
    .Y(net901));
 sky130_fd_sc_hd__clkinv_2 _143_ (.A(\mprj_dat_i_core_bar[29] ),
    .Y(net902));
 sky130_fd_sc_hd__clkinv_2 _144_ (.A(\mprj_dat_i_core_bar[30] ),
    .Y(net904));
 sky130_fd_sc_hd__clkinv_2 _145_ (.A(\mprj_dat_i_core_bar[31] ),
    .Y(net905));
 sky130_fd_sc_hd__clkinv_2 _146_ (.A(mprj_ack_i_core_bar),
    .Y(net847));
 sky130_fd_sc_hd__inv_2 _147_ (.A(\la_data_in_mprj_bar[0] ),
    .Y(net591));
 sky130_fd_sc_hd__clkinv_2 _148_ (.A(\la_data_in_mprj_bar[1] ),
    .Y(net630));
 sky130_fd_sc_hd__clkinv_2 _149_ (.A(\la_data_in_mprj_bar[2] ),
    .Y(net641));
 sky130_fd_sc_hd__clkinv_2 _150_ (.A(\la_data_in_mprj_bar[3] ),
    .Y(net652));
 sky130_fd_sc_hd__inv_2 _151_ (.A(\la_data_in_mprj_bar[4] ),
    .Y(net663));
 sky130_fd_sc_hd__clkinv_2 _152_ (.A(\la_data_in_mprj_bar[5] ),
    .Y(net674));
 sky130_fd_sc_hd__clkinv_2 _153_ (.A(\la_data_in_mprj_bar[6] ),
    .Y(net685));
 sky130_fd_sc_hd__clkinv_2 _154_ (.A(\la_data_in_mprj_bar[7] ),
    .Y(net696));
 sky130_fd_sc_hd__clkinv_2 _155_ (.A(\la_data_in_mprj_bar[8] ),
    .Y(net707));
 sky130_fd_sc_hd__clkinv_2 _156_ (.A(\la_data_in_mprj_bar[9] ),
    .Y(net718));
 sky130_fd_sc_hd__clkinv_2 _157_ (.A(\la_data_in_mprj_bar[10] ),
    .Y(net602));
 sky130_fd_sc_hd__inv_2 _158_ (.A(\la_data_in_mprj_bar[11] ),
    .Y(net613));
 sky130_fd_sc_hd__inv_2 _159_ (.A(\la_data_in_mprj_bar[12] ),
    .Y(net622));
 sky130_fd_sc_hd__inv_2 _160_ (.A(\la_data_in_mprj_bar[13] ),
    .Y(net623));
 sky130_fd_sc_hd__clkinv_2 _161_ (.A(\la_data_in_mprj_bar[14] ),
    .Y(net624));
 sky130_fd_sc_hd__clkinv_2 _162_ (.A(\la_data_in_mprj_bar[15] ),
    .Y(net625));
 sky130_fd_sc_hd__clkinv_2 _163_ (.A(\la_data_in_mprj_bar[16] ),
    .Y(net626));
 sky130_fd_sc_hd__and2_1 _164_ (.A(\mprj_logic1[331] ),
    .B(net171),
    .X(\la_data_in_enable[1] ));
 sky130_fd_sc_hd__and2_1 _165_ (.A(\mprj_logic1[332] ),
    .B(net182),
    .X(\la_data_in_enable[2] ));
 sky130_fd_sc_hd__and2_1 _166_ (.A(\mprj_logic1[333] ),
    .B(net193),
    .X(\la_data_in_enable[3] ));
 sky130_fd_sc_hd__and2_1 _167_ (.A(\mprj_logic1[334] ),
    .B(net204),
    .X(\la_data_in_enable[4] ));
 sky130_fd_sc_hd__and2_4 _168_ (.A(\mprj_logic1[335] ),
    .B(net215),
    .X(\la_data_in_enable[5] ));
 sky130_fd_sc_hd__and2_4 _169_ (.A(\mprj_logic1[336] ),
    .B(net226),
    .X(\la_data_in_enable[6] ));
 sky130_fd_sc_hd__and2_4 _170_ (.A(\mprj_logic1[337] ),
    .B(net237),
    .X(\la_data_in_enable[7] ));
 sky130_fd_sc_hd__and2_4 _171_ (.A(\mprj_logic1[338] ),
    .B(net248),
    .X(\la_data_in_enable[8] ));
 sky130_fd_sc_hd__and2_4 _172_ (.A(\mprj_logic1[339] ),
    .B(net259),
    .X(\la_data_in_enable[9] ));
 sky130_fd_sc_hd__and2_4 _173_ (.A(\mprj_logic1[340] ),
    .B(net143),
    .X(\la_data_in_enable[10] ));
 sky130_fd_sc_hd__and2_4 _174_ (.A(\mprj_logic1[341] ),
    .B(net154),
    .X(\la_data_in_enable[11] ));
 sky130_fd_sc_hd__and2_4 _175_ (.A(\mprj_logic1[342] ),
    .B(net163),
    .X(\la_data_in_enable[12] ));
 sky130_fd_sc_hd__and2_4 _176_ (.A(\mprj_logic1[343] ),
    .B(net164),
    .X(\la_data_in_enable[13] ));
 sky130_fd_sc_hd__and2_4 _177_ (.A(\mprj_logic1[344] ),
    .B(net165),
    .X(\la_data_in_enable[14] ));
 sky130_fd_sc_hd__and2_2 _178_ (.A(\mprj_logic1[345] ),
    .B(net166),
    .X(\la_data_in_enable[15] ));
 sky130_fd_sc_hd__and2_2 _179_ (.A(\mprj_logic1[346] ),
    .B(net167),
    .X(\la_data_in_enable[16] ));
 sky130_fd_sc_hd__and2_1 _180_ (.A(\mprj_logic1[347] ),
    .B(net168),
    .X(\la_data_in_enable[17] ));
 sky130_fd_sc_hd__and2_2 _181_ (.A(\mprj_logic1[348] ),
    .B(net169),
    .X(\la_data_in_enable[18] ));
 sky130_fd_sc_hd__and2_2 _182_ (.A(\mprj_logic1[349] ),
    .B(net170),
    .X(\la_data_in_enable[19] ));
 sky130_fd_sc_hd__and2_2 _183_ (.A(\mprj_logic1[350] ),
    .B(net172),
    .X(\la_data_in_enable[20] ));
 sky130_fd_sc_hd__and2_2 _184_ (.A(\mprj_logic1[351] ),
    .B(net173),
    .X(\la_data_in_enable[21] ));
 sky130_fd_sc_hd__and2_2 _185_ (.A(\mprj_logic1[352] ),
    .B(net174),
    .X(\la_data_in_enable[22] ));
 sky130_fd_sc_hd__and2_1 _186_ (.A(\mprj_logic1[353] ),
    .B(net175),
    .X(\la_data_in_enable[23] ));
 sky130_fd_sc_hd__and2_2 _187_ (.A(\mprj_logic1[354] ),
    .B(net176),
    .X(\la_data_in_enable[24] ));
 sky130_fd_sc_hd__and2_2 _188_ (.A(\mprj_logic1[355] ),
    .B(net177),
    .X(\la_data_in_enable[25] ));
 sky130_fd_sc_hd__and2_2 _189_ (.A(\mprj_logic1[356] ),
    .B(net178),
    .X(\la_data_in_enable[26] ));
 sky130_fd_sc_hd__and2_2 _190_ (.A(\mprj_logic1[357] ),
    .B(net179),
    .X(\la_data_in_enable[27] ));
 sky130_fd_sc_hd__and2_2 _191_ (.A(\mprj_logic1[358] ),
    .B(net180),
    .X(\la_data_in_enable[28] ));
 sky130_fd_sc_hd__and2_2 _192_ (.A(\mprj_logic1[359] ),
    .B(net181),
    .X(\la_data_in_enable[29] ));
 sky130_fd_sc_hd__and2_2 _193_ (.A(\mprj_logic1[360] ),
    .B(net183),
    .X(\la_data_in_enable[30] ));
 sky130_fd_sc_hd__and2_1 _194_ (.A(\mprj_logic1[361] ),
    .B(net184),
    .X(\la_data_in_enable[31] ));
 sky130_fd_sc_hd__and2_2 _195_ (.A(\mprj_logic1[362] ),
    .B(net185),
    .X(\la_data_in_enable[32] ));
 sky130_fd_sc_hd__and2_2 _196_ (.A(\mprj_logic1[363] ),
    .B(net186),
    .X(\la_data_in_enable[33] ));
 sky130_fd_sc_hd__and2_1 _197_ (.A(\mprj_logic1[364] ),
    .B(net187),
    .X(\la_data_in_enable[34] ));
 sky130_fd_sc_hd__and2_2 _198_ (.A(\mprj_logic1[365] ),
    .B(net188),
    .X(\la_data_in_enable[35] ));
 sky130_fd_sc_hd__and2_2 _199_ (.A(\mprj_logic1[366] ),
    .B(net189),
    .X(\la_data_in_enable[36] ));
 sky130_fd_sc_hd__and2_2 _200_ (.A(\mprj_logic1[367] ),
    .B(net190),
    .X(\la_data_in_enable[37] ));
 sky130_fd_sc_hd__and2_2 _201_ (.A(\mprj_logic1[368] ),
    .B(net191),
    .X(\la_data_in_enable[38] ));
 sky130_fd_sc_hd__and2_4 _202_ (.A(\mprj_logic1[369] ),
    .B(net192),
    .X(\la_data_in_enable[39] ));
 sky130_fd_sc_hd__and2_4 _203_ (.A(\mprj_logic1[370] ),
    .B(net194),
    .X(\la_data_in_enable[40] ));
 sky130_fd_sc_hd__and2_2 _204_ (.A(\mprj_logic1[371] ),
    .B(net195),
    .X(\la_data_in_enable[41] ));
 sky130_fd_sc_hd__and2_2 _205_ (.A(\mprj_logic1[372] ),
    .B(net196),
    .X(\la_data_in_enable[42] ));
 sky130_fd_sc_hd__and2_1 _206_ (.A(\mprj_logic1[373] ),
    .B(net197),
    .X(\la_data_in_enable[43] ));
 sky130_fd_sc_hd__and2_1 _207_ (.A(\mprj_logic1[374] ),
    .B(net198),
    .X(\la_data_in_enable[44] ));
 sky130_fd_sc_hd__and2_1 _208_ (.A(\mprj_logic1[375] ),
    .B(net199),
    .X(\la_data_in_enable[45] ));
 sky130_fd_sc_hd__and2_1 _209_ (.A(\mprj_logic1[376] ),
    .B(net200),
    .X(\la_data_in_enable[46] ));
 sky130_fd_sc_hd__and2_1 _210_ (.A(\mprj_logic1[377] ),
    .B(net201),
    .X(\la_data_in_enable[47] ));
 sky130_fd_sc_hd__and2_1 _211_ (.A(\mprj_logic1[378] ),
    .B(net202),
    .X(\la_data_in_enable[48] ));
 sky130_fd_sc_hd__and2_2 _212_ (.A(\mprj_logic1[379] ),
    .B(net203),
    .X(\la_data_in_enable[49] ));
 sky130_fd_sc_hd__and2_2 _213_ (.A(\mprj_logic1[380] ),
    .B(net205),
    .X(\la_data_in_enable[50] ));
 sky130_fd_sc_hd__and2_2 _214_ (.A(\mprj_logic1[381] ),
    .B(net206),
    .X(\la_data_in_enable[51] ));
 sky130_fd_sc_hd__and2_2 _215_ (.A(\mprj_logic1[382] ),
    .B(net207),
    .X(\la_data_in_enable[52] ));
 sky130_fd_sc_hd__and2_4 _216_ (.A(\mprj_logic1[383] ),
    .B(net208),
    .X(\la_data_in_enable[53] ));
 sky130_fd_sc_hd__and2_2 _217_ (.A(\mprj_logic1[384] ),
    .B(net209),
    .X(\la_data_in_enable[54] ));
 sky130_fd_sc_hd__and2_2 _218_ (.A(\mprj_logic1[385] ),
    .B(net210),
    .X(\la_data_in_enable[55] ));
 sky130_fd_sc_hd__and2_2 _219_ (.A(\mprj_logic1[386] ),
    .B(net211),
    .X(\la_data_in_enable[56] ));
 sky130_fd_sc_hd__and2_2 _220_ (.A(\mprj_logic1[387] ),
    .B(net212),
    .X(\la_data_in_enable[57] ));
 sky130_fd_sc_hd__and2_2 _221_ (.A(\mprj_logic1[388] ),
    .B(net213),
    .X(\la_data_in_enable[58] ));
 sky130_fd_sc_hd__and2_2 _222_ (.A(\mprj_logic1[389] ),
    .B(net214),
    .X(\la_data_in_enable[59] ));
 sky130_fd_sc_hd__and2_2 _223_ (.A(\mprj_logic1[390] ),
    .B(net216),
    .X(\la_data_in_enable[60] ));
 sky130_fd_sc_hd__and2_2 _224_ (.A(\mprj_logic1[391] ),
    .B(net217),
    .X(\la_data_in_enable[61] ));
 sky130_fd_sc_hd__and2_4 _225_ (.A(\mprj_logic1[392] ),
    .B(net218),
    .X(\la_data_in_enable[62] ));
 sky130_fd_sc_hd__and2_2 _226_ (.A(\mprj_logic1[393] ),
    .B(net219),
    .X(\la_data_in_enable[63] ));
 sky130_fd_sc_hd__and2_2 _227_ (.A(\mprj_logic1[394] ),
    .B(net220),
    .X(\la_data_in_enable[64] ));
 sky130_fd_sc_hd__and2_2 _228_ (.A(\mprj_logic1[395] ),
    .B(net221),
    .X(\la_data_in_enable[65] ));
 sky130_fd_sc_hd__and2_2 _229_ (.A(\mprj_logic1[396] ),
    .B(net222),
    .X(\la_data_in_enable[66] ));
 sky130_fd_sc_hd__and2_4 _230_ (.A(\mprj_logic1[397] ),
    .B(net223),
    .X(\la_data_in_enable[67] ));
 sky130_fd_sc_hd__and2_2 _231_ (.A(\mprj_logic1[398] ),
    .B(net224),
    .X(\la_data_in_enable[68] ));
 sky130_fd_sc_hd__and2_2 _232_ (.A(\mprj_logic1[399] ),
    .B(net225),
    .X(\la_data_in_enable[69] ));
 sky130_fd_sc_hd__and2_2 _233_ (.A(\mprj_logic1[400] ),
    .B(net227),
    .X(\la_data_in_enable[70] ));
 sky130_fd_sc_hd__and2_4 _234_ (.A(\mprj_logic1[401] ),
    .B(net228),
    .X(\la_data_in_enable[71] ));
 sky130_fd_sc_hd__and2_4 _235_ (.A(\mprj_logic1[402] ),
    .B(net229),
    .X(\la_data_in_enable[72] ));
 sky130_fd_sc_hd__and2_4 _236_ (.A(\mprj_logic1[403] ),
    .B(net230),
    .X(\la_data_in_enable[73] ));
 sky130_fd_sc_hd__and2_4 _237_ (.A(\mprj_logic1[404] ),
    .B(net231),
    .X(\la_data_in_enable[74] ));
 sky130_fd_sc_hd__and2_4 _238_ (.A(\mprj_logic1[405] ),
    .B(net232),
    .X(\la_data_in_enable[75] ));
 sky130_fd_sc_hd__and2_4 _239_ (.A(\mprj_logic1[406] ),
    .B(net233),
    .X(\la_data_in_enable[76] ));
 sky130_fd_sc_hd__and2_4 _240_ (.A(\mprj_logic1[407] ),
    .B(net234),
    .X(\la_data_in_enable[77] ));
 sky130_fd_sc_hd__and2_4 _241_ (.A(\mprj_logic1[408] ),
    .B(net235),
    .X(\la_data_in_enable[78] ));
 sky130_fd_sc_hd__and2_4 _242_ (.A(\mprj_logic1[409] ),
    .B(net236),
    .X(\la_data_in_enable[79] ));
 sky130_fd_sc_hd__and2_4 _243_ (.A(\mprj_logic1[410] ),
    .B(net238),
    .X(\la_data_in_enable[80] ));
 sky130_fd_sc_hd__and2_4 _244_ (.A(\mprj_logic1[411] ),
    .B(net239),
    .X(\la_data_in_enable[81] ));
 sky130_fd_sc_hd__and2_4 _245_ (.A(\mprj_logic1[412] ),
    .B(net240),
    .X(\la_data_in_enable[82] ));
 sky130_fd_sc_hd__and2_4 _246_ (.A(\mprj_logic1[413] ),
    .B(net241),
    .X(\la_data_in_enable[83] ));
 sky130_fd_sc_hd__and2_4 _247_ (.A(\mprj_logic1[414] ),
    .B(net242),
    .X(\la_data_in_enable[84] ));
 sky130_fd_sc_hd__and2_4 _248_ (.A(\mprj_logic1[415] ),
    .B(net243),
    .X(\la_data_in_enable[85] ));
 sky130_fd_sc_hd__and2_4 _249_ (.A(\mprj_logic1[416] ),
    .B(net244),
    .X(\la_data_in_enable[86] ));
 sky130_fd_sc_hd__and2_4 _250_ (.A(\mprj_logic1[417] ),
    .B(net245),
    .X(\la_data_in_enable[87] ));
 sky130_fd_sc_hd__and2_4 _251_ (.A(\mprj_logic1[418] ),
    .B(net246),
    .X(\la_data_in_enable[88] ));
 sky130_fd_sc_hd__and2_4 _252_ (.A(\mprj_logic1[419] ),
    .B(net247),
    .X(\la_data_in_enable[89] ));
 sky130_fd_sc_hd__and2_4 _253_ (.A(\mprj_logic1[420] ),
    .B(net249),
    .X(\la_data_in_enable[90] ));
 sky130_fd_sc_hd__and2_4 _254_ (.A(\mprj_logic1[421] ),
    .B(net250),
    .X(\la_data_in_enable[91] ));
 sky130_fd_sc_hd__and2_4 _255_ (.A(\mprj_logic1[422] ),
    .B(net251),
    .X(\la_data_in_enable[92] ));
 sky130_fd_sc_hd__and2_4 _256_ (.A(\mprj_logic1[423] ),
    .B(net252),
    .X(\la_data_in_enable[93] ));
 sky130_fd_sc_hd__and2_4 _257_ (.A(\mprj_logic1[424] ),
    .B(net253),
    .X(\la_data_in_enable[94] ));
 sky130_fd_sc_hd__and2_4 _258_ (.A(\mprj_logic1[425] ),
    .B(net254),
    .X(\la_data_in_enable[95] ));
 sky130_fd_sc_hd__and2_4 _259_ (.A(\mprj_logic1[426] ),
    .B(net255),
    .X(\la_data_in_enable[96] ));
 sky130_fd_sc_hd__and2_4 _260_ (.A(\mprj_logic1[427] ),
    .B(net256),
    .X(\la_data_in_enable[97] ));
 sky130_fd_sc_hd__and2_4 _261_ (.A(\mprj_logic1[428] ),
    .B(net257),
    .X(\la_data_in_enable[98] ));
 sky130_fd_sc_hd__and2_4 _262_ (.A(\mprj_logic1[429] ),
    .B(net258),
    .X(\la_data_in_enable[99] ));
 sky130_fd_sc_hd__and2_4 _263_ (.A(\mprj_logic1[430] ),
    .B(net133),
    .X(\la_data_in_enable[100] ));
 sky130_fd_sc_hd__and2_4 _264_ (.A(\mprj_logic1[431] ),
    .B(net134),
    .X(\la_data_in_enable[101] ));
 sky130_fd_sc_hd__and2_4 _265_ (.A(\mprj_logic1[432] ),
    .B(net135),
    .X(\la_data_in_enable[102] ));
 sky130_fd_sc_hd__and2_4 _266_ (.A(\mprj_logic1[433] ),
    .B(net136),
    .X(\la_data_in_enable[103] ));
 sky130_fd_sc_hd__and2_4 _267_ (.A(\mprj_logic1[434] ),
    .B(net137),
    .X(\la_data_in_enable[104] ));
 sky130_fd_sc_hd__and2_4 _268_ (.A(\mprj_logic1[435] ),
    .B(net138),
    .X(\la_data_in_enable[105] ));
 sky130_fd_sc_hd__and2_4 _269_ (.A(\mprj_logic1[436] ),
    .B(net139),
    .X(\la_data_in_enable[106] ));
 sky130_fd_sc_hd__and2_4 _270_ (.A(\mprj_logic1[437] ),
    .B(net140),
    .X(\la_data_in_enable[107] ));
 sky130_fd_sc_hd__and2_4 _271_ (.A(\mprj_logic1[438] ),
    .B(net141),
    .X(\la_data_in_enable[108] ));
 sky130_fd_sc_hd__and2_4 _272_ (.A(\mprj_logic1[439] ),
    .B(net142),
    .X(\la_data_in_enable[109] ));
 sky130_fd_sc_hd__and2_4 _273_ (.A(\mprj_logic1[440] ),
    .B(net144),
    .X(\la_data_in_enable[110] ));
 sky130_fd_sc_hd__and2_4 _274_ (.A(\mprj_logic1[441] ),
    .B(net145),
    .X(\la_data_in_enable[111] ));
 sky130_fd_sc_hd__and2_4 _275_ (.A(\mprj_logic1[442] ),
    .B(net146),
    .X(\la_data_in_enable[112] ));
 sky130_fd_sc_hd__and2_4 _276_ (.A(\mprj_logic1[443] ),
    .B(net147),
    .X(\la_data_in_enable[113] ));
 sky130_fd_sc_hd__and2_4 _277_ (.A(\mprj_logic1[444] ),
    .B(net148),
    .X(\la_data_in_enable[114] ));
 sky130_fd_sc_hd__and2_4 _278_ (.A(\mprj_logic1[445] ),
    .B(net149),
    .X(\la_data_in_enable[115] ));
 sky130_fd_sc_hd__and2_4 _279_ (.A(\mprj_logic1[446] ),
    .B(net150),
    .X(\la_data_in_enable[116] ));
 sky130_fd_sc_hd__and2_4 _280_ (.A(\mprj_logic1[447] ),
    .B(net151),
    .X(\la_data_in_enable[117] ));
 sky130_fd_sc_hd__and2_4 _281_ (.A(\mprj_logic1[448] ),
    .B(net152),
    .X(\la_data_in_enable[118] ));
 sky130_fd_sc_hd__and2_2 _282_ (.A(\mprj_logic1[449] ),
    .B(net153),
    .X(\la_data_in_enable[119] ));
 sky130_fd_sc_hd__and2_4 _283_ (.A(\mprj_logic1[450] ),
    .B(net155),
    .X(\la_data_in_enable[120] ));
 sky130_fd_sc_hd__and2_4 _284_ (.A(\mprj_logic1[451] ),
    .B(net156),
    .X(\la_data_in_enable[121] ));
 sky130_fd_sc_hd__and2_4 _285_ (.A(\mprj_logic1[452] ),
    .B(net157),
    .X(\la_data_in_enable[122] ));
 sky130_fd_sc_hd__and2_4 _286_ (.A(\mprj_logic1[453] ),
    .B(net158),
    .X(\la_data_in_enable[123] ));
 sky130_fd_sc_hd__and2_4 _287_ (.A(\mprj_logic1[454] ),
    .B(net159),
    .X(\la_data_in_enable[124] ));
 sky130_fd_sc_hd__and2_4 _288_ (.A(\mprj_logic1[455] ),
    .B(net160),
    .X(\la_data_in_enable[125] ));
 sky130_fd_sc_hd__and2_4 _289_ (.A(\mprj_logic1[456] ),
    .B(net161),
    .X(\la_data_in_enable[126] ));
 sky130_fd_sc_hd__and2_4 _290_ (.A(\mprj_logic1[457] ),
    .B(net162),
    .X(\la_data_in_enable[127] ));
 sky130_fd_sc_hd__and2_1 _291_ (.A(\mprj_logic1[458] ),
    .B(net460),
    .X(\user_irq_enable[0] ));
 sky130_fd_sc_hd__and2_1 _292_ (.A(\mprj_logic1[459] ),
    .B(net461),
    .X(\user_irq_enable[1] ));
 sky130_fd_sc_hd__and2_1 _293_ (.A(\mprj_logic1[460] ),
    .B(net462),
    .X(\user_irq_enable[2] ));
 sky130_fd_sc_hd__and2_4 _294_ (.A(\mprj_logic1[462] ),
    .B(net453),
    .X(wb_in_enable));
 sky130_fd_sc_hd__and2b_4 _295_ (.A_N(net3),
    .B(\mprj_logic1[0] ),
    .X(net960));
 sky130_fd_sc_hd__and2_4 _296_ (.A(\mprj_logic1[1] ),
    .B(net1),
    .X(net955));
 sky130_fd_sc_hd__and2_2 _297_ (.A(\mprj_logic1[2] ),
    .B(net2),
    .X(net956));
 sky130_fd_sc_hd__and2_4 _298_ (.A(\mprj_logic1[3] ),
    .B(net420),
    .X(net880));
 sky130_fd_sc_hd__and2_4 _299_ (.A(\mprj_logic1[4] ),
    .B(net458),
    .X(net949));
 sky130_fd_sc_hd__and2_4 _300_ (.A(\mprj_logic1[5] ),
    .B(net459),
    .X(net950));
 sky130_fd_sc_hd__and2_4 _301_ (.A(\mprj_logic1[6] ),
    .B(net454),
    .X(net945));
 sky130_fd_sc_hd__and2_4 _302_ (.A(\mprj_logic1[7] ),
    .B(net455),
    .X(net946));
 sky130_fd_sc_hd__and2_4 _303_ (.A(\mprj_logic1[8] ),
    .B(net456),
    .X(net947));
 sky130_fd_sc_hd__and2_4 _304_ (.A(\mprj_logic1[9] ),
    .B(net457),
    .X(net948));
 sky130_fd_sc_hd__and2_4 _305_ (.A(\mprj_logic1[10] ),
    .B(net388),
    .X(net848));
 sky130_fd_sc_hd__and2_4 _306_ (.A(\mprj_logic1[11] ),
    .B(net399),
    .X(net859));
 sky130_fd_sc_hd__and2_2 _307_ (.A(\mprj_logic1[12] ),
    .B(net410),
    .X(net870));
 sky130_fd_sc_hd__and2_4 _308_ (.A(\mprj_logic1[13] ),
    .B(net413),
    .X(net873));
 sky130_fd_sc_hd__and2_2 _309_ (.A(\mprj_logic1[14] ),
    .B(net414),
    .X(net874));
 sky130_fd_sc_hd__and2_4 _310_ (.A(\mprj_logic1[15] ),
    .B(net415),
    .X(net875));
 sky130_fd_sc_hd__and2_4 _311_ (.A(\mprj_logic1[16] ),
    .B(net416),
    .X(net876));
 sky130_fd_sc_hd__and2_4 _312_ (.A(\mprj_logic1[17] ),
    .B(net417),
    .X(net877));
 sky130_fd_sc_hd__and2_4 _313_ (.A(\mprj_logic1[18] ),
    .B(net418),
    .X(net878));
 sky130_fd_sc_hd__and2_4 _314_ (.A(\mprj_logic1[19] ),
    .B(net419),
    .X(net879));
 sky130_fd_sc_hd__and2_4 _315_ (.A(\mprj_logic1[20] ),
    .B(net389),
    .X(net849));
 sky130_fd_sc_hd__and2_4 _316_ (.A(\mprj_logic1[21] ),
    .B(net390),
    .X(net850));
 sky130_fd_sc_hd__and2_4 _317_ (.A(\mprj_logic1[22] ),
    .B(net391),
    .X(net851));
 sky130_fd_sc_hd__and2_4 _318_ (.A(\mprj_logic1[23] ),
    .B(net392),
    .X(net852));
 sky130_fd_sc_hd__and2_4 _319_ (.A(\mprj_logic1[24] ),
    .B(net393),
    .X(net853));
 sky130_fd_sc_hd__and2_4 _320_ (.A(\mprj_logic1[25] ),
    .B(net394),
    .X(net854));
 sky130_fd_sc_hd__and2_4 _321_ (.A(\mprj_logic1[26] ),
    .B(net395),
    .X(net855));
 sky130_fd_sc_hd__and2_4 _322_ (.A(\mprj_logic1[27] ),
    .B(net396),
    .X(net856));
 sky130_fd_sc_hd__and2_4 _323_ (.A(\mprj_logic1[28] ),
    .B(net397),
    .X(net857));
 sky130_fd_sc_hd__and2_4 _324_ (.A(\mprj_logic1[29] ),
    .B(net398),
    .X(net858));
 sky130_fd_sc_hd__and2_4 _325_ (.A(\mprj_logic1[30] ),
    .B(net400),
    .X(net860));
 sky130_fd_sc_hd__and2_4 _326_ (.A(\mprj_logic1[31] ),
    .B(net401),
    .X(net861));
 sky130_fd_sc_hd__and2_4 _327_ (.A(\mprj_logic1[32] ),
    .B(net402),
    .X(net862));
 sky130_fd_sc_hd__and2_4 _328_ (.A(\mprj_logic1[33] ),
    .B(net403),
    .X(net863));
 sky130_fd_sc_hd__and2_4 _329_ (.A(\mprj_logic1[34] ),
    .B(net404),
    .X(net864));
 sky130_fd_sc_hd__and2_4 _330_ (.A(\mprj_logic1[35] ),
    .B(net405),
    .X(net865));
 sky130_fd_sc_hd__and2_4 _331_ (.A(\mprj_logic1[36] ),
    .B(net406),
    .X(net866));
 sky130_fd_sc_hd__and2_4 _332_ (.A(\mprj_logic1[37] ),
    .B(net407),
    .X(net867));
 sky130_fd_sc_hd__and2_4 _333_ (.A(\mprj_logic1[38] ),
    .B(net408),
    .X(net868));
 sky130_fd_sc_hd__and2_4 _334_ (.A(\mprj_logic1[39] ),
    .B(net409),
    .X(net869));
 sky130_fd_sc_hd__and2_2 _335_ (.A(\mprj_logic1[40] ),
    .B(net411),
    .X(net871));
 sky130_fd_sc_hd__and2_4 _336_ (.A(\mprj_logic1[41] ),
    .B(net412),
    .X(net872));
 sky130_fd_sc_hd__and2_4 _337_ (.A(\mprj_logic1[42] ),
    .B(net421),
    .X(net913));
 sky130_fd_sc_hd__and2_4 _338_ (.A(\mprj_logic1[43] ),
    .B(net432),
    .X(net924));
 sky130_fd_sc_hd__and2_4 _339_ (.A(\mprj_logic1[44] ),
    .B(net443),
    .X(net935));
 sky130_fd_sc_hd__and2_4 _340_ (.A(\mprj_logic1[45] ),
    .B(net446),
    .X(net938));
 sky130_fd_sc_hd__and2_4 _341_ (.A(\mprj_logic1[46] ),
    .B(net447),
    .X(net939));
 sky130_fd_sc_hd__and2_4 _342_ (.A(\mprj_logic1[47] ),
    .B(net448),
    .X(net940));
 sky130_fd_sc_hd__and2_4 _343_ (.A(\mprj_logic1[48] ),
    .B(net449),
    .X(net941));
 sky130_fd_sc_hd__and2_4 _344_ (.A(\mprj_logic1[49] ),
    .B(net450),
    .X(net942));
 sky130_fd_sc_hd__and2_4 _345_ (.A(\mprj_logic1[50] ),
    .B(net451),
    .X(net943));
 sky130_fd_sc_hd__and2_4 _346_ (.A(\mprj_logic1[51] ),
    .B(net452),
    .X(net944));
 sky130_fd_sc_hd__and2_4 _347_ (.A(\mprj_logic1[52] ),
    .B(net422),
    .X(net914));
 sky130_fd_sc_hd__and2_4 _348_ (.A(\mprj_logic1[53] ),
    .B(net423),
    .X(net915));
 sky130_fd_sc_hd__and2_4 _349_ (.A(\mprj_logic1[54] ),
    .B(net424),
    .X(net916));
 sky130_fd_sc_hd__and2_4 _350_ (.A(\mprj_logic1[55] ),
    .B(net425),
    .X(net917));
 sky130_fd_sc_hd__and2_4 _351_ (.A(\mprj_logic1[56] ),
    .B(net426),
    .X(net918));
 sky130_fd_sc_hd__and2_4 _352_ (.A(\mprj_logic1[57] ),
    .B(net427),
    .X(net919));
 sky130_fd_sc_hd__and2_4 _353_ (.A(\mprj_logic1[58] ),
    .B(net428),
    .X(net920));
 sky130_fd_sc_hd__and2_4 _354_ (.A(\mprj_logic1[59] ),
    .B(net429),
    .X(net921));
 sky130_fd_sc_hd__and2_4 _355_ (.A(\mprj_logic1[60] ),
    .B(net430),
    .X(net922));
 sky130_fd_sc_hd__and2_4 _356_ (.A(\mprj_logic1[61] ),
    .B(net431),
    .X(net923));
 sky130_fd_sc_hd__and2_4 _357_ (.A(\mprj_logic1[62] ),
    .B(net433),
    .X(net925));
 sky130_fd_sc_hd__and2_4 _358_ (.A(\mprj_logic1[63] ),
    .B(net434),
    .X(net926));
 sky130_fd_sc_hd__and2_4 _359_ (.A(\mprj_logic1[64] ),
    .B(net435),
    .X(net927));
 sky130_fd_sc_hd__and2_4 _360_ (.A(\mprj_logic1[65] ),
    .B(net436),
    .X(net928));
 sky130_fd_sc_hd__and2_4 _361_ (.A(\mprj_logic1[66] ),
    .B(net437),
    .X(net929));
 sky130_fd_sc_hd__and2_4 _362_ (.A(\mprj_logic1[67] ),
    .B(net438),
    .X(net930));
 sky130_fd_sc_hd__and2_4 _363_ (.A(\mprj_logic1[68] ),
    .B(net439),
    .X(net931));
 sky130_fd_sc_hd__and2_4 _364_ (.A(\mprj_logic1[69] ),
    .B(net440),
    .X(net932));
 sky130_fd_sc_hd__and2_4 _365_ (.A(\mprj_logic1[70] ),
    .B(net441),
    .X(net933));
 sky130_fd_sc_hd__and2_4 _366_ (.A(\mprj_logic1[71] ),
    .B(net442),
    .X(net934));
 sky130_fd_sc_hd__and2_4 _367_ (.A(\mprj_logic1[72] ),
    .B(net444),
    .X(net936));
 sky130_fd_sc_hd__and2_4 _368_ (.A(\mprj_logic1[73] ),
    .B(net445),
    .X(net937));
 sky130_fd_sc_hd__and3b_4 _369_ (.A_N(net260),
    .B(\mprj_logic1[74] ),
    .C(net4),
    .X(net463));
 sky130_fd_sc_hd__and3b_4 _370_ (.A_N(net299),
    .B(\mprj_logic1[75] ),
    .C(net43),
    .X(net502));
 sky130_fd_sc_hd__and3b_4 _371_ (.A_N(net310),
    .B(\mprj_logic1[76] ),
    .C(net54),
    .X(net513));
 sky130_fd_sc_hd__and3b_4 _372_ (.A_N(net321),
    .B(\mprj_logic1[77] ),
    .C(net65),
    .X(net524));
 sky130_fd_sc_hd__and3b_4 _373_ (.A_N(net332),
    .B(\mprj_logic1[78] ),
    .C(net76),
    .X(net535));
 sky130_fd_sc_hd__and3b_4 _374_ (.A_N(net343),
    .B(\mprj_logic1[79] ),
    .C(net87),
    .X(net546));
 sky130_fd_sc_hd__and3b_4 _375_ (.A_N(net354),
    .B(\mprj_logic1[80] ),
    .C(net98),
    .X(net557));
 sky130_fd_sc_hd__and3b_4 _376_ (.A_N(net365),
    .B(\mprj_logic1[81] ),
    .C(net109),
    .X(net568));
 sky130_fd_sc_hd__and3b_4 _377_ (.A_N(net376),
    .B(\mprj_logic1[82] ),
    .C(net120),
    .X(net579));
 sky130_fd_sc_hd__and3b_4 _378_ (.A_N(net387),
    .B(\mprj_logic1[83] ),
    .C(net131),
    .X(net590));
 sky130_fd_sc_hd__and3b_4 _379_ (.A_N(net271),
    .B(\mprj_logic1[84] ),
    .C(net15),
    .X(net474));
 sky130_fd_sc_hd__and3b_4 _380_ (.A_N(net282),
    .B(\mprj_logic1[85] ),
    .C(net26),
    .X(net485));
 sky130_fd_sc_hd__and3b_4 _381_ (.A_N(net291),
    .B(\mprj_logic1[86] ),
    .C(net35),
    .X(net494));
 sky130_fd_sc_hd__and3b_4 _382_ (.A_N(net292),
    .B(\mprj_logic1[87] ),
    .C(net36),
    .X(net495));
 sky130_fd_sc_hd__and3b_4 _383_ (.A_N(net293),
    .B(\mprj_logic1[88] ),
    .C(net37),
    .X(net496));
 sky130_fd_sc_hd__and3b_4 _384_ (.A_N(net294),
    .B(\mprj_logic1[89] ),
    .C(net38),
    .X(net497));
 sky130_fd_sc_hd__and3b_4 _385_ (.A_N(net295),
    .B(\mprj_logic1[90] ),
    .C(net39),
    .X(net498));
 sky130_fd_sc_hd__and3b_4 _386_ (.A_N(net296),
    .B(\mprj_logic1[91] ),
    .C(net40),
    .X(net499));
 sky130_fd_sc_hd__and3b_4 _387_ (.A_N(net297),
    .B(\mprj_logic1[92] ),
    .C(net41),
    .X(net500));
 sky130_fd_sc_hd__and3b_4 _388_ (.A_N(net298),
    .B(\mprj_logic1[93] ),
    .C(net42),
    .X(net501));
 sky130_fd_sc_hd__and3b_4 _389_ (.A_N(net300),
    .B(\mprj_logic1[94] ),
    .C(net44),
    .X(net503));
 sky130_fd_sc_hd__and3b_4 _390_ (.A_N(net301),
    .B(\mprj_logic1[95] ),
    .C(net45),
    .X(net504));
 sky130_fd_sc_hd__and3b_4 _391_ (.A_N(net302),
    .B(\mprj_logic1[96] ),
    .C(net46),
    .X(net505));
 sky130_fd_sc_hd__and3b_4 _392_ (.A_N(net303),
    .B(\mprj_logic1[97] ),
    .C(net47),
    .X(net506));
 sky130_fd_sc_hd__and3b_4 _393_ (.A_N(net304),
    .B(\mprj_logic1[98] ),
    .C(net48),
    .X(net507));
 sky130_fd_sc_hd__and3b_4 _394_ (.A_N(net305),
    .B(\mprj_logic1[99] ),
    .C(net49),
    .X(net508));
 sky130_fd_sc_hd__and3b_4 _395_ (.A_N(net306),
    .B(\mprj_logic1[100] ),
    .C(net50),
    .X(net509));
 sky130_fd_sc_hd__and3b_4 _396_ (.A_N(net307),
    .B(\mprj_logic1[101] ),
    .C(net51),
    .X(net510));
 sky130_fd_sc_hd__and3b_4 _397_ (.A_N(net308),
    .B(\mprj_logic1[102] ),
    .C(net52),
    .X(net511));
 sky130_fd_sc_hd__and3b_4 _398_ (.A_N(net309),
    .B(\mprj_logic1[103] ),
    .C(net53),
    .X(net512));
 sky130_fd_sc_hd__and3b_4 _399_ (.A_N(net311),
    .B(\mprj_logic1[104] ),
    .C(net55),
    .X(net514));
 sky130_fd_sc_hd__and3b_4 _400_ (.A_N(net312),
    .B(\mprj_logic1[105] ),
    .C(net56),
    .X(net515));
 sky130_fd_sc_hd__and3b_4 _401_ (.A_N(net313),
    .B(\mprj_logic1[106] ),
    .C(net57),
    .X(net516));
 sky130_fd_sc_hd__and3b_4 _402_ (.A_N(net314),
    .B(\mprj_logic1[107] ),
    .C(net58),
    .X(net517));
 sky130_fd_sc_hd__and3b_4 _403_ (.A_N(net315),
    .B(\mprj_logic1[108] ),
    .C(net59),
    .X(net518));
 sky130_fd_sc_hd__and3b_4 _404_ (.A_N(net316),
    .B(\mprj_logic1[109] ),
    .C(net60),
    .X(net519));
 sky130_fd_sc_hd__and3b_4 _405_ (.A_N(net317),
    .B(\mprj_logic1[110] ),
    .C(net61),
    .X(net520));
 sky130_fd_sc_hd__and3b_4 _406_ (.A_N(net318),
    .B(\mprj_logic1[111] ),
    .C(net62),
    .X(net521));
 sky130_fd_sc_hd__and3b_4 _407_ (.A_N(net319),
    .B(\mprj_logic1[112] ),
    .C(net63),
    .X(net522));
 sky130_fd_sc_hd__and3b_4 _408_ (.A_N(net320),
    .B(\mprj_logic1[113] ),
    .C(net64),
    .X(net523));
 sky130_fd_sc_hd__and3b_4 _409_ (.A_N(net322),
    .B(\mprj_logic1[114] ),
    .C(net66),
    .X(net525));
 sky130_fd_sc_hd__and3b_4 _410_ (.A_N(net323),
    .B(\mprj_logic1[115] ),
    .C(net67),
    .X(net526));
 sky130_fd_sc_hd__and3b_4 _411_ (.A_N(net324),
    .B(\mprj_logic1[116] ),
    .C(net68),
    .X(net527));
 sky130_fd_sc_hd__and3b_4 _412_ (.A_N(net325),
    .B(\mprj_logic1[117] ),
    .C(net69),
    .X(net528));
 sky130_fd_sc_hd__and3b_4 _413_ (.A_N(net326),
    .B(\mprj_logic1[118] ),
    .C(net70),
    .X(net529));
 sky130_fd_sc_hd__and3b_4 _414_ (.A_N(net327),
    .B(\mprj_logic1[119] ),
    .C(net71),
    .X(net530));
 sky130_fd_sc_hd__and3b_4 _415_ (.A_N(net328),
    .B(\mprj_logic1[120] ),
    .C(net72),
    .X(net531));
 sky130_fd_sc_hd__and3b_4 _416_ (.A_N(net329),
    .B(\mprj_logic1[121] ),
    .C(net73),
    .X(net532));
 sky130_fd_sc_hd__and3b_4 _417_ (.A_N(net330),
    .B(\mprj_logic1[122] ),
    .C(net74),
    .X(net533));
 sky130_fd_sc_hd__and3b_4 _418_ (.A_N(net331),
    .B(\mprj_logic1[123] ),
    .C(net75),
    .X(net534));
 sky130_fd_sc_hd__and3b_4 _419_ (.A_N(net333),
    .B(\mprj_logic1[124] ),
    .C(net77),
    .X(net536));
 sky130_fd_sc_hd__and3b_4 _420_ (.A_N(net334),
    .B(\mprj_logic1[125] ),
    .C(net78),
    .X(net537));
 sky130_fd_sc_hd__and3b_4 _421_ (.A_N(net335),
    .B(\mprj_logic1[126] ),
    .C(net79),
    .X(net538));
 sky130_fd_sc_hd__and3b_4 _422_ (.A_N(net336),
    .B(\mprj_logic1[127] ),
    .C(net80),
    .X(net539));
 sky130_fd_sc_hd__and3b_4 _423_ (.A_N(net337),
    .B(\mprj_logic1[128] ),
    .C(net81),
    .X(net540));
 sky130_fd_sc_hd__and3b_4 _424_ (.A_N(net338),
    .B(\mprj_logic1[129] ),
    .C(net82),
    .X(net541));
 sky130_fd_sc_hd__and3b_4 _425_ (.A_N(net339),
    .B(\mprj_logic1[130] ),
    .C(net83),
    .X(net542));
 sky130_fd_sc_hd__and3b_4 _426_ (.A_N(net340),
    .B(\mprj_logic1[131] ),
    .C(net84),
    .X(net543));
 sky130_fd_sc_hd__and3b_4 _427_ (.A_N(net341),
    .B(\mprj_logic1[132] ),
    .C(net85),
    .X(net544));
 sky130_fd_sc_hd__and3b_4 _428_ (.A_N(net342),
    .B(\mprj_logic1[133] ),
    .C(net86),
    .X(net545));
 sky130_fd_sc_hd__and3b_4 _429_ (.A_N(net344),
    .B(\mprj_logic1[134] ),
    .C(net88),
    .X(net547));
 sky130_fd_sc_hd__and3b_4 _430_ (.A_N(net345),
    .B(\mprj_logic1[135] ),
    .C(net89),
    .X(net548));
 sky130_fd_sc_hd__and3b_4 _431_ (.A_N(net346),
    .B(\mprj_logic1[136] ),
    .C(net90),
    .X(net549));
 sky130_fd_sc_hd__and3b_4 _432_ (.A_N(net347),
    .B(\mprj_logic1[137] ),
    .C(net91),
    .X(net550));
 sky130_fd_sc_hd__and3b_4 _433_ (.A_N(net348),
    .B(\mprj_logic1[138] ),
    .C(net92),
    .X(net551));
 sky130_fd_sc_hd__and3b_4 _434_ (.A_N(net349),
    .B(\mprj_logic1[139] ),
    .C(net93),
    .X(net552));
 sky130_fd_sc_hd__and3b_4 _435_ (.A_N(net350),
    .B(\mprj_logic1[140] ),
    .C(net94),
    .X(net553));
 sky130_fd_sc_hd__and3b_4 _436_ (.A_N(net351),
    .B(\mprj_logic1[141] ),
    .C(net95),
    .X(net554));
 sky130_fd_sc_hd__and3b_4 _437_ (.A_N(net352),
    .B(\mprj_logic1[142] ),
    .C(net96),
    .X(net555));
 sky130_fd_sc_hd__and3b_4 _438_ (.A_N(net353),
    .B(\mprj_logic1[143] ),
    .C(net97),
    .X(net556));
 sky130_fd_sc_hd__and3b_4 _439_ (.A_N(net355),
    .B(\mprj_logic1[144] ),
    .C(net99),
    .X(net558));
 sky130_fd_sc_hd__and3b_4 _440_ (.A_N(net356),
    .B(\mprj_logic1[145] ),
    .C(net100),
    .X(net559));
 sky130_fd_sc_hd__and3b_4 _441_ (.A_N(net357),
    .B(\mprj_logic1[146] ),
    .C(net101),
    .X(net560));
 sky130_fd_sc_hd__and3b_4 _442_ (.A_N(net358),
    .B(\mprj_logic1[147] ),
    .C(net102),
    .X(net561));
 sky130_fd_sc_hd__and3b_4 _443_ (.A_N(net359),
    .B(\mprj_logic1[148] ),
    .C(net103),
    .X(net562));
 sky130_fd_sc_hd__and3b_4 _444_ (.A_N(net360),
    .B(\mprj_logic1[149] ),
    .C(net104),
    .X(net563));
 sky130_fd_sc_hd__and3b_4 _445_ (.A_N(net361),
    .B(\mprj_logic1[150] ),
    .C(net105),
    .X(net564));
 sky130_fd_sc_hd__and3b_4 _446_ (.A_N(net362),
    .B(\mprj_logic1[151] ),
    .C(net106),
    .X(net565));
 sky130_fd_sc_hd__and3b_4 _447_ (.A_N(net363),
    .B(\mprj_logic1[152] ),
    .C(net107),
    .X(net566));
 sky130_fd_sc_hd__and3b_4 _448_ (.A_N(net364),
    .B(\mprj_logic1[153] ),
    .C(net108),
    .X(net567));
 sky130_fd_sc_hd__and3b_4 _449_ (.A_N(net366),
    .B(\mprj_logic1[154] ),
    .C(net110),
    .X(net569));
 sky130_fd_sc_hd__and3b_4 _450_ (.A_N(net367),
    .B(\mprj_logic1[155] ),
    .C(net111),
    .X(net570));
 sky130_fd_sc_hd__and3b_4 _451_ (.A_N(net368),
    .B(\mprj_logic1[156] ),
    .C(net112),
    .X(net571));
 sky130_fd_sc_hd__and3b_4 _452_ (.A_N(net369),
    .B(\mprj_logic1[157] ),
    .C(net113),
    .X(net572));
 sky130_fd_sc_hd__and3b_4 _453_ (.A_N(net370),
    .B(\mprj_logic1[158] ),
    .C(net114),
    .X(net573));
 sky130_fd_sc_hd__and3b_4 _454_ (.A_N(net371),
    .B(\mprj_logic1[159] ),
    .C(net115),
    .X(net574));
 sky130_fd_sc_hd__and3b_4 _455_ (.A_N(net372),
    .B(\mprj_logic1[160] ),
    .C(net116),
    .X(net575));
 sky130_fd_sc_hd__and3b_4 _456_ (.A_N(net373),
    .B(\mprj_logic1[161] ),
    .C(net117),
    .X(net576));
 sky130_fd_sc_hd__and3b_4 _457_ (.A_N(net374),
    .B(\mprj_logic1[162] ),
    .C(net118),
    .X(net577));
 sky130_fd_sc_hd__and3b_4 _458_ (.A_N(net375),
    .B(\mprj_logic1[163] ),
    .C(net119),
    .X(net578));
 sky130_fd_sc_hd__and3b_4 _459_ (.A_N(net377),
    .B(\mprj_logic1[164] ),
    .C(net121),
    .X(net580));
 sky130_fd_sc_hd__and3b_4 _460_ (.A_N(net378),
    .B(\mprj_logic1[165] ),
    .C(net122),
    .X(net581));
 sky130_fd_sc_hd__and3b_4 _461_ (.A_N(net379),
    .B(\mprj_logic1[166] ),
    .C(net123),
    .X(net582));
 sky130_fd_sc_hd__and3b_4 _462_ (.A_N(net380),
    .B(\mprj_logic1[167] ),
    .C(net124),
    .X(net583));
 sky130_fd_sc_hd__and3b_4 _463_ (.A_N(net381),
    .B(\mprj_logic1[168] ),
    .C(net125),
    .X(net584));
 sky130_fd_sc_hd__and3b_4 _464_ (.A_N(net382),
    .B(\mprj_logic1[169] ),
    .C(net126),
    .X(net585));
 sky130_fd_sc_hd__and3b_4 _465_ (.A_N(net383),
    .B(\mprj_logic1[170] ),
    .C(net127),
    .X(net586));
 sky130_fd_sc_hd__and3b_4 _466_ (.A_N(net384),
    .B(\mprj_logic1[171] ),
    .C(net128),
    .X(net587));
 sky130_fd_sc_hd__and3b_4 _467_ (.A_N(net385),
    .B(\mprj_logic1[172] ),
    .C(net129),
    .X(net588));
 sky130_fd_sc_hd__and3b_4 _468_ (.A_N(net386),
    .B(\mprj_logic1[173] ),
    .C(net130),
    .X(net589));
 sky130_fd_sc_hd__and3b_4 _469_ (.A_N(net261),
    .B(\mprj_logic1[174] ),
    .C(net5),
    .X(net464));
 sky130_fd_sc_hd__and3b_4 _470_ (.A_N(net262),
    .B(\mprj_logic1[175] ),
    .C(net6),
    .X(net465));
 sky130_fd_sc_hd__and3b_4 _471_ (.A_N(net263),
    .B(\mprj_logic1[176] ),
    .C(net7),
    .X(net466));
 sky130_fd_sc_hd__and3b_4 _472_ (.A_N(net264),
    .B(\mprj_logic1[177] ),
    .C(net8),
    .X(net467));
 sky130_fd_sc_hd__and3b_4 _473_ (.A_N(net265),
    .B(\mprj_logic1[178] ),
    .C(net9),
    .X(net468));
 sky130_fd_sc_hd__and3b_4 _474_ (.A_N(net266),
    .B(\mprj_logic1[179] ),
    .C(net10),
    .X(net469));
 sky130_fd_sc_hd__and3b_4 _475_ (.A_N(net267),
    .B(\mprj_logic1[180] ),
    .C(net11),
    .X(net470));
 sky130_fd_sc_hd__and3b_4 _476_ (.A_N(net268),
    .B(\mprj_logic1[181] ),
    .C(net12),
    .X(net471));
 sky130_fd_sc_hd__and3b_4 _477_ (.A_N(net269),
    .B(\mprj_logic1[182] ),
    .C(net13),
    .X(net472));
 sky130_fd_sc_hd__and3b_4 _478_ (.A_N(net270),
    .B(\mprj_logic1[183] ),
    .C(net14),
    .X(net473));
 sky130_fd_sc_hd__and3b_4 _479_ (.A_N(net272),
    .B(\mprj_logic1[184] ),
    .C(net16),
    .X(net475));
 sky130_fd_sc_hd__and3b_4 _480_ (.A_N(net273),
    .B(\mprj_logic1[185] ),
    .C(net17),
    .X(net476));
 sky130_fd_sc_hd__and3b_4 _481_ (.A_N(net274),
    .B(\mprj_logic1[186] ),
    .C(net18),
    .X(net477));
 sky130_fd_sc_hd__and3b_4 _482_ (.A_N(net275),
    .B(\mprj_logic1[187] ),
    .C(net19),
    .X(net478));
 sky130_fd_sc_hd__and3b_4 _483_ (.A_N(net276),
    .B(\mprj_logic1[188] ),
    .C(net20),
    .X(net479));
 sky130_fd_sc_hd__and3b_4 _484_ (.A_N(net277),
    .B(\mprj_logic1[189] ),
    .C(net21),
    .X(net480));
 sky130_fd_sc_hd__and3b_4 _485_ (.A_N(net278),
    .B(\mprj_logic1[190] ),
    .C(net22),
    .X(net481));
 sky130_fd_sc_hd__and3b_4 _486_ (.A_N(net279),
    .B(\mprj_logic1[191] ),
    .C(net23),
    .X(net482));
 sky130_fd_sc_hd__and3b_4 _487_ (.A_N(net280),
    .B(\mprj_logic1[192] ),
    .C(net24),
    .X(net483));
 sky130_fd_sc_hd__and3b_4 _488_ (.A_N(net281),
    .B(\mprj_logic1[193] ),
    .C(net25),
    .X(net484));
 sky130_fd_sc_hd__and3b_4 _489_ (.A_N(net283),
    .B(\mprj_logic1[194] ),
    .C(net27),
    .X(net486));
 sky130_fd_sc_hd__and3b_4 _490_ (.A_N(net284),
    .B(\mprj_logic1[195] ),
    .C(net28),
    .X(net487));
 sky130_fd_sc_hd__and3b_4 _491_ (.A_N(net285),
    .B(\mprj_logic1[196] ),
    .C(net29),
    .X(net488));
 sky130_fd_sc_hd__and3b_4 _492_ (.A_N(net286),
    .B(\mprj_logic1[197] ),
    .C(net30),
    .X(net489));
 sky130_fd_sc_hd__and3b_4 _493_ (.A_N(net287),
    .B(\mprj_logic1[198] ),
    .C(net31),
    .X(net490));
 sky130_fd_sc_hd__and3b_4 _494_ (.A_N(net288),
    .B(\mprj_logic1[199] ),
    .C(net32),
    .X(net491));
 sky130_fd_sc_hd__and3b_4 _495_ (.A_N(net289),
    .B(\mprj_logic1[200] ),
    .C(net33),
    .X(net492));
 sky130_fd_sc_hd__and3b_4 _496_ (.A_N(net290),
    .B(\mprj_logic1[201] ),
    .C(net34),
    .X(net493));
 sky130_fd_sc_hd__and2_4 _497_ (.A(net260),
    .B(\mprj_logic1[202] ),
    .X(net719));
 sky130_fd_sc_hd__and2_4 _498_ (.A(net299),
    .B(\mprj_logic1[203] ),
    .X(net758));
 sky130_fd_sc_hd__and2_4 _499_ (.A(net310),
    .B(\mprj_logic1[204] ),
    .X(net769));
 sky130_fd_sc_hd__and2_4 _500_ (.A(net321),
    .B(\mprj_logic1[205] ),
    .X(net780));
 sky130_fd_sc_hd__and2_4 _501_ (.A(net332),
    .B(\mprj_logic1[206] ),
    .X(net791));
 sky130_fd_sc_hd__and2_4 _502_ (.A(net343),
    .B(\mprj_logic1[207] ),
    .X(net802));
 sky130_fd_sc_hd__and2_4 _503_ (.A(net354),
    .B(\mprj_logic1[208] ),
    .X(net813));
 sky130_fd_sc_hd__and2_4 _504_ (.A(net365),
    .B(\mprj_logic1[209] ),
    .X(net824));
 sky130_fd_sc_hd__and2_4 _505_ (.A(net376),
    .B(\mprj_logic1[210] ),
    .X(net835));
 sky130_fd_sc_hd__and2_4 _506_ (.A(net387),
    .B(\mprj_logic1[211] ),
    .X(net846));
 sky130_fd_sc_hd__and2_4 _507_ (.A(net271),
    .B(\mprj_logic1[212] ),
    .X(net730));
 sky130_fd_sc_hd__and2_4 _508_ (.A(net282),
    .B(\mprj_logic1[213] ),
    .X(net741));
 sky130_fd_sc_hd__and2_4 _509_ (.A(net291),
    .B(\mprj_logic1[214] ),
    .X(net750));
 sky130_fd_sc_hd__and2_4 _510_ (.A(net292),
    .B(\mprj_logic1[215] ),
    .X(net751));
 sky130_fd_sc_hd__and2_4 _511_ (.A(net293),
    .B(\mprj_logic1[216] ),
    .X(net752));
 sky130_fd_sc_hd__and2_4 _512_ (.A(net294),
    .B(\mprj_logic1[217] ),
    .X(net753));
 sky130_fd_sc_hd__and2_4 _513_ (.A(net295),
    .B(\mprj_logic1[218] ),
    .X(net754));
 sky130_fd_sc_hd__and2_4 _514_ (.A(net296),
    .B(\mprj_logic1[219] ),
    .X(net755));
 sky130_fd_sc_hd__and2_4 _515_ (.A(net297),
    .B(\mprj_logic1[220] ),
    .X(net756));
 sky130_fd_sc_hd__and2_4 _516_ (.A(net298),
    .B(\mprj_logic1[221] ),
    .X(net757));
 sky130_fd_sc_hd__and2_4 _517_ (.A(net300),
    .B(\mprj_logic1[222] ),
    .X(net759));
 sky130_fd_sc_hd__and2_4 _518_ (.A(net301),
    .B(\mprj_logic1[223] ),
    .X(net760));
 sky130_fd_sc_hd__and2_4 _519_ (.A(net302),
    .B(\mprj_logic1[224] ),
    .X(net761));
 sky130_fd_sc_hd__and2_4 _520_ (.A(net303),
    .B(\mprj_logic1[225] ),
    .X(net762));
 sky130_fd_sc_hd__and2_4 _521_ (.A(net304),
    .B(\mprj_logic1[226] ),
    .X(net763));
 sky130_fd_sc_hd__and2_4 _522_ (.A(net305),
    .B(\mprj_logic1[227] ),
    .X(net764));
 sky130_fd_sc_hd__and2_4 _523_ (.A(net306),
    .B(\mprj_logic1[228] ),
    .X(net765));
 sky130_fd_sc_hd__and2_4 _524_ (.A(net307),
    .B(\mprj_logic1[229] ),
    .X(net766));
 sky130_fd_sc_hd__and2_4 _525_ (.A(net308),
    .B(\mprj_logic1[230] ),
    .X(net767));
 sky130_fd_sc_hd__and2_4 _526_ (.A(net309),
    .B(\mprj_logic1[231] ),
    .X(net768));
 sky130_fd_sc_hd__and2_4 _527_ (.A(net311),
    .B(\mprj_logic1[232] ),
    .X(net770));
 sky130_fd_sc_hd__and2_4 _528_ (.A(net312),
    .B(\mprj_logic1[233] ),
    .X(net771));
 sky130_fd_sc_hd__and2_4 _529_ (.A(net313),
    .B(\mprj_logic1[234] ),
    .X(net772));
 sky130_fd_sc_hd__and2_4 _530_ (.A(net314),
    .B(\mprj_logic1[235] ),
    .X(net773));
 sky130_fd_sc_hd__and2_4 _531_ (.A(net315),
    .B(\mprj_logic1[236] ),
    .X(net774));
 sky130_fd_sc_hd__and2_4 _532_ (.A(net316),
    .B(\mprj_logic1[237] ),
    .X(net775));
 sky130_fd_sc_hd__and2_4 _533_ (.A(net317),
    .B(\mprj_logic1[238] ),
    .X(net776));
 sky130_fd_sc_hd__and2_4 _534_ (.A(net318),
    .B(\mprj_logic1[239] ),
    .X(net777));
 sky130_fd_sc_hd__and2_4 _535_ (.A(net319),
    .B(\mprj_logic1[240] ),
    .X(net778));
 sky130_fd_sc_hd__and2_4 _536_ (.A(net320),
    .B(\mprj_logic1[241] ),
    .X(net779));
 sky130_fd_sc_hd__and2_4 _537_ (.A(net322),
    .B(\mprj_logic1[242] ),
    .X(net781));
 sky130_fd_sc_hd__and2_4 _538_ (.A(net323),
    .B(\mprj_logic1[243] ),
    .X(net782));
 sky130_fd_sc_hd__and2_4 _539_ (.A(net324),
    .B(\mprj_logic1[244] ),
    .X(net783));
 sky130_fd_sc_hd__and2_4 _540_ (.A(net325),
    .B(\mprj_logic1[245] ),
    .X(net784));
 sky130_fd_sc_hd__and2_4 _541_ (.A(net326),
    .B(\mprj_logic1[246] ),
    .X(net785));
 sky130_fd_sc_hd__and2_4 _542_ (.A(net327),
    .B(\mprj_logic1[247] ),
    .X(net786));
 sky130_fd_sc_hd__and2_4 _543_ (.A(net328),
    .B(\mprj_logic1[248] ),
    .X(net787));
 sky130_fd_sc_hd__and2_4 _544_ (.A(net329),
    .B(\mprj_logic1[249] ),
    .X(net788));
 sky130_fd_sc_hd__and2_4 _545_ (.A(net330),
    .B(\mprj_logic1[250] ),
    .X(net789));
 sky130_fd_sc_hd__and2_4 _546_ (.A(net331),
    .B(\mprj_logic1[251] ),
    .X(net790));
 sky130_fd_sc_hd__and2_4 _547_ (.A(net333),
    .B(\mprj_logic1[252] ),
    .X(net792));
 sky130_fd_sc_hd__and2_4 _548_ (.A(net334),
    .B(\mprj_logic1[253] ),
    .X(net793));
 sky130_fd_sc_hd__and2_4 _549_ (.A(net335),
    .B(\mprj_logic1[254] ),
    .X(net794));
 sky130_fd_sc_hd__and2_4 _550_ (.A(net336),
    .B(\mprj_logic1[255] ),
    .X(net795));
 sky130_fd_sc_hd__and2_4 _551_ (.A(net337),
    .B(\mprj_logic1[256] ),
    .X(net796));
 sky130_fd_sc_hd__and2_4 _552_ (.A(net338),
    .B(\mprj_logic1[257] ),
    .X(net797));
 sky130_fd_sc_hd__and2_4 _553_ (.A(net339),
    .B(\mprj_logic1[258] ),
    .X(net798));
 sky130_fd_sc_hd__and2_4 _554_ (.A(net340),
    .B(\mprj_logic1[259] ),
    .X(net799));
 sky130_fd_sc_hd__and2_4 _555_ (.A(net341),
    .B(\mprj_logic1[260] ),
    .X(net800));
 sky130_fd_sc_hd__and2_4 _556_ (.A(net342),
    .B(\mprj_logic1[261] ),
    .X(net801));
 sky130_fd_sc_hd__and2_4 _557_ (.A(net344),
    .B(\mprj_logic1[262] ),
    .X(net803));
 sky130_fd_sc_hd__and2_4 _558_ (.A(net345),
    .B(\mprj_logic1[263] ),
    .X(net804));
 sky130_fd_sc_hd__and2_4 _559_ (.A(net346),
    .B(\mprj_logic1[264] ),
    .X(net805));
 sky130_fd_sc_hd__and2_4 _560_ (.A(net347),
    .B(\mprj_logic1[265] ),
    .X(net806));
 sky130_fd_sc_hd__and2_4 _561_ (.A(net348),
    .B(\mprj_logic1[266] ),
    .X(net807));
 sky130_fd_sc_hd__and2_2 _562_ (.A(net349),
    .B(\mprj_logic1[267] ),
    .X(net808));
 sky130_fd_sc_hd__and2_4 _563_ (.A(net350),
    .B(\mprj_logic1[268] ),
    .X(net809));
 sky130_fd_sc_hd__and2_2 _564_ (.A(net351),
    .B(\mprj_logic1[269] ),
    .X(net810));
 sky130_fd_sc_hd__and2_4 _565_ (.A(net352),
    .B(\mprj_logic1[270] ),
    .X(net811));
 sky130_fd_sc_hd__and2_4 _566_ (.A(net353),
    .B(\mprj_logic1[271] ),
    .X(net812));
 sky130_fd_sc_hd__and2_4 _567_ (.A(net355),
    .B(\mprj_logic1[272] ),
    .X(net814));
 sky130_fd_sc_hd__and2_4 _568_ (.A(net356),
    .B(\mprj_logic1[273] ),
    .X(net815));
 sky130_fd_sc_hd__and2_4 _569_ (.A(net357),
    .B(\mprj_logic1[274] ),
    .X(net816));
 sky130_fd_sc_hd__and2_4 _570_ (.A(net358),
    .B(\mprj_logic1[275] ),
    .X(net817));
 sky130_fd_sc_hd__and2_4 _571_ (.A(net359),
    .B(\mprj_logic1[276] ),
    .X(net818));
 sky130_fd_sc_hd__and2_4 _572_ (.A(net360),
    .B(\mprj_logic1[277] ),
    .X(net819));
 sky130_fd_sc_hd__and2_4 _573_ (.A(net361),
    .B(\mprj_logic1[278] ),
    .X(net820));
 sky130_fd_sc_hd__and2_4 _574_ (.A(net362),
    .B(\mprj_logic1[279] ),
    .X(net821));
 sky130_fd_sc_hd__and2_4 _575_ (.A(net363),
    .B(\mprj_logic1[280] ),
    .X(net822));
 sky130_fd_sc_hd__and2_4 _576_ (.A(net364),
    .B(\mprj_logic1[281] ),
    .X(net823));
 sky130_fd_sc_hd__and2_4 _577_ (.A(net366),
    .B(\mprj_logic1[282] ),
    .X(net825));
 sky130_fd_sc_hd__and2_4 _578_ (.A(net367),
    .B(\mprj_logic1[283] ),
    .X(net826));
 sky130_fd_sc_hd__and2_4 _579_ (.A(net368),
    .B(\mprj_logic1[284] ),
    .X(net827));
 sky130_fd_sc_hd__and2_4 _580_ (.A(net369),
    .B(\mprj_logic1[285] ),
    .X(net828));
 sky130_fd_sc_hd__and2_4 _581_ (.A(net370),
    .B(\mprj_logic1[286] ),
    .X(net829));
 sky130_fd_sc_hd__and2_4 _582_ (.A(net371),
    .B(\mprj_logic1[287] ),
    .X(net830));
 sky130_fd_sc_hd__and2_4 _583_ (.A(net372),
    .B(\mprj_logic1[288] ),
    .X(net831));
 sky130_fd_sc_hd__and2_4 _584_ (.A(net373),
    .B(\mprj_logic1[289] ),
    .X(net832));
 sky130_fd_sc_hd__and2_4 _585_ (.A(net374),
    .B(\mprj_logic1[290] ),
    .X(net833));
 sky130_fd_sc_hd__and2_4 _586_ (.A(net375),
    .B(\mprj_logic1[291] ),
    .X(net834));
 sky130_fd_sc_hd__and2_4 _587_ (.A(net377),
    .B(\mprj_logic1[292] ),
    .X(net836));
 sky130_fd_sc_hd__and2_4 _588_ (.A(net378),
    .B(\mprj_logic1[293] ),
    .X(net837));
 sky130_fd_sc_hd__and2_4 _589_ (.A(net379),
    .B(\mprj_logic1[294] ),
    .X(net838));
 sky130_fd_sc_hd__and2_4 _590_ (.A(net380),
    .B(\mprj_logic1[295] ),
    .X(net839));
 sky130_fd_sc_hd__and2_4 _591_ (.A(net381),
    .B(\mprj_logic1[296] ),
    .X(net840));
 sky130_fd_sc_hd__and2_4 _592_ (.A(net382),
    .B(\mprj_logic1[297] ),
    .X(net841));
 sky130_fd_sc_hd__and2_4 _593_ (.A(net383),
    .B(\mprj_logic1[298] ),
    .X(net842));
 sky130_fd_sc_hd__and2_4 _594_ (.A(net384),
    .B(\mprj_logic1[299] ),
    .X(net843));
 sky130_fd_sc_hd__and2_2 _595_ (.A(net385),
    .B(\mprj_logic1[300] ),
    .X(net844));
 sky130_fd_sc_hd__and2_4 _596_ (.A(net386),
    .B(\mprj_logic1[301] ),
    .X(net845));
 sky130_fd_sc_hd__and2_4 _597_ (.A(net261),
    .B(\mprj_logic1[302] ),
    .X(net720));
 sky130_fd_sc_hd__and2_4 _598_ (.A(net262),
    .B(\mprj_logic1[303] ),
    .X(net721));
 sky130_fd_sc_hd__and2_4 _599_ (.A(net263),
    .B(\mprj_logic1[304] ),
    .X(net722));
 sky130_fd_sc_hd__and2_4 _600_ (.A(net264),
    .B(\mprj_logic1[305] ),
    .X(net723));
 sky130_fd_sc_hd__and2_4 _601_ (.A(net265),
    .B(\mprj_logic1[306] ),
    .X(net724));
 sky130_fd_sc_hd__and2_4 _602_ (.A(net266),
    .B(\mprj_logic1[307] ),
    .X(net725));
 sky130_fd_sc_hd__and2_4 _603_ (.A(net267),
    .B(\mprj_logic1[308] ),
    .X(net726));
 sky130_fd_sc_hd__and2_4 _604_ (.A(net268),
    .B(\mprj_logic1[309] ),
    .X(net727));
 sky130_fd_sc_hd__and2_4 _605_ (.A(net269),
    .B(\mprj_logic1[310] ),
    .X(net728));
 sky130_fd_sc_hd__and2_4 _606_ (.A(net270),
    .B(\mprj_logic1[311] ),
    .X(net729));
 sky130_fd_sc_hd__and2_4 _607_ (.A(net272),
    .B(\mprj_logic1[312] ),
    .X(net731));
 sky130_fd_sc_hd__and2_4 _608_ (.A(net273),
    .B(\mprj_logic1[313] ),
    .X(net732));
 sky130_fd_sc_hd__and2_4 _609_ (.A(net274),
    .B(\mprj_logic1[314] ),
    .X(net733));
 sky130_fd_sc_hd__and2_4 _610_ (.A(net275),
    .B(\mprj_logic1[315] ),
    .X(net734));
 sky130_fd_sc_hd__and2_4 _611_ (.A(net276),
    .B(\mprj_logic1[316] ),
    .X(net735));
 sky130_fd_sc_hd__and2_4 _612_ (.A(net277),
    .B(\mprj_logic1[317] ),
    .X(net736));
 sky130_fd_sc_hd__and2_4 _613_ (.A(net278),
    .B(\mprj_logic1[318] ),
    .X(net737));
 sky130_fd_sc_hd__and2_4 _614_ (.A(net279),
    .B(\mprj_logic1[319] ),
    .X(net738));
 sky130_fd_sc_hd__and2_4 _615_ (.A(net280),
    .B(\mprj_logic1[320] ),
    .X(net739));
 sky130_fd_sc_hd__and2_4 _616_ (.A(net281),
    .B(\mprj_logic1[321] ),
    .X(net740));
 sky130_fd_sc_hd__and2_4 _617_ (.A(net283),
    .B(\mprj_logic1[322] ),
    .X(net742));
 sky130_fd_sc_hd__and2_4 _618_ (.A(net284),
    .B(\mprj_logic1[323] ),
    .X(net743));
 sky130_fd_sc_hd__and2_4 _619_ (.A(net285),
    .B(\mprj_logic1[324] ),
    .X(net744));
 sky130_fd_sc_hd__and2_4 _620_ (.A(net286),
    .B(\mprj_logic1[325] ),
    .X(net745));
 sky130_fd_sc_hd__and2_4 _621_ (.A(net287),
    .B(\mprj_logic1[326] ),
    .X(net746));
 sky130_fd_sc_hd__and2_4 _622_ (.A(net288),
    .B(\mprj_logic1[327] ),
    .X(net747));
 sky130_fd_sc_hd__and2_4 _623_ (.A(net289),
    .B(\mprj_logic1[328] ),
    .X(net748));
 sky130_fd_sc_hd__and2_4 _624_ (.A(net290),
    .B(\mprj_logic1[329] ),
    .X(net749));
 sky130_fd_sc_hd__and2_1 _625_ (.A(\mprj_logic1[330] ),
    .B(net132),
    .X(\la_data_in_enable[0] ));
 mprj2_logic_high mprj2_logic_high_inst (.HI(net953));
 mprj_logic_high mprj_logic_high_inst (.HI({\mprj_logic1[462] ,
    net951,
    \mprj_logic1[460] ,
    \mprj_logic1[459] ,
    \mprj_logic1[458] ,
    \mprj_logic1[457] ,
    \mprj_logic1[456] ,
    \mprj_logic1[455] ,
    \mprj_logic1[454] ,
    \mprj_logic1[453] ,
    \mprj_logic1[452] ,
    \mprj_logic1[451] ,
    \mprj_logic1[450] ,
    \mprj_logic1[449] ,
    \mprj_logic1[448] ,
    \mprj_logic1[447] ,
    \mprj_logic1[446] ,
    \mprj_logic1[445] ,
    \mprj_logic1[444] ,
    \mprj_logic1[443] ,
    \mprj_logic1[442] ,
    \mprj_logic1[441] ,
    \mprj_logic1[440] ,
    \mprj_logic1[439] ,
    \mprj_logic1[438] ,
    \mprj_logic1[437] ,
    \mprj_logic1[436] ,
    \mprj_logic1[435] ,
    \mprj_logic1[434] ,
    \mprj_logic1[433] ,
    \mprj_logic1[432] ,
    \mprj_logic1[431] ,
    \mprj_logic1[430] ,
    \mprj_logic1[429] ,
    \mprj_logic1[428] ,
    \mprj_logic1[427] ,
    \mprj_logic1[426] ,
    \mprj_logic1[425] ,
    \mprj_logic1[424] ,
    \mprj_logic1[423] ,
    \mprj_logic1[422] ,
    \mprj_logic1[421] ,
    \mprj_logic1[420] ,
    \mprj_logic1[419] ,
    \mprj_logic1[418] ,
    \mprj_logic1[417] ,
    \mprj_logic1[416] ,
    \mprj_logic1[415] ,
    \mprj_logic1[414] ,
    \mprj_logic1[413] ,
    \mprj_logic1[412] ,
    \mprj_logic1[411] ,
    \mprj_logic1[410] ,
    \mprj_logic1[409] ,
    \mprj_logic1[408] ,
    \mprj_logic1[407] ,
    \mprj_logic1[406] ,
    \mprj_logic1[405] ,
    \mprj_logic1[404] ,
    \mprj_logic1[403] ,
    \mprj_logic1[402] ,
    \mprj_logic1[401] ,
    \mprj_logic1[400] ,
    \mprj_logic1[399] ,
    \mprj_logic1[398] ,
    \mprj_logic1[397] ,
    \mprj_logic1[396] ,
    \mprj_logic1[395] ,
    \mprj_logic1[394] ,
    \mprj_logic1[393] ,
    \mprj_logic1[392] ,
    \mprj_logic1[391] ,
    \mprj_logic1[390] ,
    \mprj_logic1[389] ,
    \mprj_logic1[388] ,
    \mprj_logic1[387] ,
    \mprj_logic1[386] ,
    \mprj_logic1[385] ,
    \mprj_logic1[384] ,
    \mprj_logic1[383] ,
    \mprj_logic1[382] ,
    \mprj_logic1[381] ,
    \mprj_logic1[380] ,
    \mprj_logic1[379] ,
    \mprj_logic1[378] ,
    \mprj_logic1[377] ,
    \mprj_logic1[376] ,
    \mprj_logic1[375] ,
    \mprj_logic1[374] ,
    \mprj_logic1[373] ,
    \mprj_logic1[372] ,
    \mprj_logic1[371] ,
    \mprj_logic1[370] ,
    \mprj_logic1[369] ,
    \mprj_logic1[368] ,
    \mprj_logic1[367] ,
    \mprj_logic1[366] ,
    \mprj_logic1[365] ,
    \mprj_logic1[364] ,
    \mprj_logic1[363] ,
    \mprj_logic1[362] ,
    \mprj_logic1[361] ,
    \mprj_logic1[360] ,
    \mprj_logic1[359] ,
    \mprj_logic1[358] ,
    \mprj_logic1[357] ,
    \mprj_logic1[356] ,
    \mprj_logic1[355] ,
    \mprj_logic1[354] ,
    \mprj_logic1[353] ,
    \mprj_logic1[352] ,
    \mprj_logic1[351] ,
    \mprj_logic1[350] ,
    \mprj_logic1[349] ,
    \mprj_logic1[348] ,
    \mprj_logic1[347] ,
    \mprj_logic1[346] ,
    \mprj_logic1[345] ,
    \mprj_logic1[344] ,
    \mprj_logic1[343] ,
    \mprj_logic1[342] ,
    \mprj_logic1[341] ,
    \mprj_logic1[340] ,
    \mprj_logic1[339] ,
    \mprj_logic1[338] ,
    \mprj_logic1[337] ,
    \mprj_logic1[336] ,
    \mprj_logic1[335] ,
    \mprj_logic1[334] ,
    \mprj_logic1[333] ,
    \mprj_logic1[332] ,
    \mprj_logic1[331] ,
    \mprj_logic1[330] ,
    \mprj_logic1[329] ,
    \mprj_logic1[328] ,
    \mprj_logic1[327] ,
    \mprj_logic1[326] ,
    \mprj_logic1[325] ,
    \mprj_logic1[324] ,
    \mprj_logic1[323] ,
    \mprj_logic1[322] ,
    \mprj_logic1[321] ,
    \mprj_logic1[320] ,
    \mprj_logic1[319] ,
    \mprj_logic1[318] ,
    \mprj_logic1[317] ,
    \mprj_logic1[316] ,
    \mprj_logic1[315] ,
    \mprj_logic1[314] ,
    \mprj_logic1[313] ,
    \mprj_logic1[312] ,
    \mprj_logic1[311] ,
    \mprj_logic1[310] ,
    \mprj_logic1[309] ,
    \mprj_logic1[308] ,
    \mprj_logic1[307] ,
    \mprj_logic1[306] ,
    \mprj_logic1[305] ,
    \mprj_logic1[304] ,
    \mprj_logic1[303] ,
    \mprj_logic1[302] ,
    \mprj_logic1[301] ,
    \mprj_logic1[300] ,
    \mprj_logic1[299] ,
    \mprj_logic1[298] ,
    \mprj_logic1[297] ,
    \mprj_logic1[296] ,
    \mprj_logic1[295] ,
    \mprj_logic1[294] ,
    \mprj_logic1[293] ,
    \mprj_logic1[292] ,
    \mprj_logic1[291] ,
    \mprj_logic1[290] ,
    \mprj_logic1[289] ,
    \mprj_logic1[288] ,
    \mprj_logic1[287] ,
    \mprj_logic1[286] ,
    \mprj_logic1[285] ,
    \mprj_logic1[284] ,
    \mprj_logic1[283] ,
    \mprj_logic1[282] ,
    \mprj_logic1[281] ,
    \mprj_logic1[280] ,
    \mprj_logic1[279] ,
    \mprj_logic1[278] ,
    \mprj_logic1[277] ,
    \mprj_logic1[276] ,
    \mprj_logic1[275] ,
    \mprj_logic1[274] ,
    \mprj_logic1[273] ,
    \mprj_logic1[272] ,
    \mprj_logic1[271] ,
    \mprj_logic1[270] ,
    \mprj_logic1[269] ,
    \mprj_logic1[268] ,
    \mprj_logic1[267] ,
    \mprj_logic1[266] ,
    \mprj_logic1[265] ,
    \mprj_logic1[264] ,
    \mprj_logic1[263] ,
    \mprj_logic1[262] ,
    \mprj_logic1[261] ,
    \mprj_logic1[260] ,
    \mprj_logic1[259] ,
    \mprj_logic1[258] ,
    \mprj_logic1[257] ,
    \mprj_logic1[256] ,
    \mprj_logic1[255] ,
    \mprj_logic1[254] ,
    \mprj_logic1[253] ,
    \mprj_logic1[252] ,
    \mprj_logic1[251] ,
    \mprj_logic1[250] ,
    \mprj_logic1[249] ,
    \mprj_logic1[248] ,
    \mprj_logic1[247] ,
    \mprj_logic1[246] ,
    \mprj_logic1[245] ,
    \mprj_logic1[244] ,
    \mprj_logic1[243] ,
    \mprj_logic1[242] ,
    \mprj_logic1[241] ,
    \mprj_logic1[240] ,
    \mprj_logic1[239] ,
    \mprj_logic1[238] ,
    \mprj_logic1[237] ,
    \mprj_logic1[236] ,
    \mprj_logic1[235] ,
    \mprj_logic1[234] ,
    \mprj_logic1[233] ,
    \mprj_logic1[232] ,
    \mprj_logic1[231] ,
    \mprj_logic1[230] ,
    \mprj_logic1[229] ,
    \mprj_logic1[228] ,
    \mprj_logic1[227] ,
    \mprj_logic1[226] ,
    \mprj_logic1[225] ,
    \mprj_logic1[224] ,
    \mprj_logic1[223] ,
    \mprj_logic1[222] ,
    \mprj_logic1[221] ,
    \mprj_logic1[220] ,
    \mprj_logic1[219] ,
    \mprj_logic1[218] ,
    \mprj_logic1[217] ,
    \mprj_logic1[216] ,
    \mprj_logic1[215] ,
    \mprj_logic1[214] ,
    \mprj_logic1[213] ,
    \mprj_logic1[212] ,
    \mprj_logic1[211] ,
    \mprj_logic1[210] ,
    \mprj_logic1[209] ,
    \mprj_logic1[208] ,
    \mprj_logic1[207] ,
    \mprj_logic1[206] ,
    \mprj_logic1[205] ,
    \mprj_logic1[204] ,
    \mprj_logic1[203] ,
    \mprj_logic1[202] ,
    \mprj_logic1[201] ,
    \mprj_logic1[200] ,
    \mprj_logic1[199] ,
    \mprj_logic1[198] ,
    \mprj_logic1[197] ,
    \mprj_logic1[196] ,
    \mprj_logic1[195] ,
    \mprj_logic1[194] ,
    \mprj_logic1[193] ,
    \mprj_logic1[192] ,
    \mprj_logic1[191] ,
    \mprj_logic1[190] ,
    \mprj_logic1[189] ,
    \mprj_logic1[188] ,
    \mprj_logic1[187] ,
    \mprj_logic1[186] ,
    \mprj_logic1[185] ,
    \mprj_logic1[184] ,
    \mprj_logic1[183] ,
    \mprj_logic1[182] ,
    \mprj_logic1[181] ,
    \mprj_logic1[180] ,
    \mprj_logic1[179] ,
    \mprj_logic1[178] ,
    \mprj_logic1[177] ,
    \mprj_logic1[176] ,
    \mprj_logic1[175] ,
    \mprj_logic1[174] ,
    \mprj_logic1[173] ,
    \mprj_logic1[172] ,
    \mprj_logic1[171] ,
    \mprj_logic1[170] ,
    \mprj_logic1[169] ,
    \mprj_logic1[168] ,
    \mprj_logic1[167] ,
    \mprj_logic1[166] ,
    \mprj_logic1[165] ,
    \mprj_logic1[164] ,
    \mprj_logic1[163] ,
    \mprj_logic1[162] ,
    \mprj_logic1[161] ,
    \mprj_logic1[160] ,
    \mprj_logic1[159] ,
    \mprj_logic1[158] ,
    \mprj_logic1[157] ,
    \mprj_logic1[156] ,
    \mprj_logic1[155] ,
    \mprj_logic1[154] ,
    \mprj_logic1[153] ,
    \mprj_logic1[152] ,
    \mprj_logic1[151] ,
    \mprj_logic1[150] ,
    \mprj_logic1[149] ,
    \mprj_logic1[148] ,
    \mprj_logic1[147] ,
    \mprj_logic1[146] ,
    \mprj_logic1[145] ,
    \mprj_logic1[144] ,
    \mprj_logic1[143] ,
    \mprj_logic1[142] ,
    \mprj_logic1[141] ,
    \mprj_logic1[140] ,
    \mprj_logic1[139] ,
    \mprj_logic1[138] ,
    \mprj_logic1[137] ,
    \mprj_logic1[136] ,
    \mprj_logic1[135] ,
    \mprj_logic1[134] ,
    \mprj_logic1[133] ,
    \mprj_logic1[132] ,
    \mprj_logic1[131] ,
    \mprj_logic1[130] ,
    \mprj_logic1[129] ,
    \mprj_logic1[128] ,
    \mprj_logic1[127] ,
    \mprj_logic1[126] ,
    \mprj_logic1[125] ,
    \mprj_logic1[124] ,
    \mprj_logic1[123] ,
    \mprj_logic1[122] ,
    \mprj_logic1[121] ,
    \mprj_logic1[120] ,
    \mprj_logic1[119] ,
    \mprj_logic1[118] ,
    \mprj_logic1[117] ,
    \mprj_logic1[116] ,
    \mprj_logic1[115] ,
    \mprj_logic1[114] ,
    \mprj_logic1[113] ,
    \mprj_logic1[112] ,
    \mprj_logic1[111] ,
    \mprj_logic1[110] ,
    \mprj_logic1[109] ,
    \mprj_logic1[108] ,
    \mprj_logic1[107] ,
    \mprj_logic1[106] ,
    \mprj_logic1[105] ,
    \mprj_logic1[104] ,
    \mprj_logic1[103] ,
    \mprj_logic1[102] ,
    \mprj_logic1[101] ,
    \mprj_logic1[100] ,
    \mprj_logic1[99] ,
    \mprj_logic1[98] ,
    \mprj_logic1[97] ,
    \mprj_logic1[96] ,
    \mprj_logic1[95] ,
    \mprj_logic1[94] ,
    \mprj_logic1[93] ,
    \mprj_logic1[92] ,
    \mprj_logic1[91] ,
    \mprj_logic1[90] ,
    \mprj_logic1[89] ,
    \mprj_logic1[88] ,
    \mprj_logic1[87] ,
    \mprj_logic1[86] ,
    \mprj_logic1[85] ,
    \mprj_logic1[84] ,
    \mprj_logic1[83] ,
    \mprj_logic1[82] ,
    \mprj_logic1[81] ,
    \mprj_logic1[80] ,
    \mprj_logic1[79] ,
    \mprj_logic1[78] ,
    \mprj_logic1[77] ,
    \mprj_logic1[76] ,
    \mprj_logic1[75] ,
    \mprj_logic1[74] ,
    \mprj_logic1[73] ,
    \mprj_logic1[72] ,
    \mprj_logic1[71] ,
    \mprj_logic1[70] ,
    \mprj_logic1[69] ,
    \mprj_logic1[68] ,
    \mprj_logic1[67] ,
    \mprj_logic1[66] ,
    \mprj_logic1[65] ,
    \mprj_logic1[64] ,
    \mprj_logic1[63] ,
    \mprj_logic1[62] ,
    \mprj_logic1[61] ,
    \mprj_logic1[60] ,
    \mprj_logic1[59] ,
    \mprj_logic1[58] ,
    \mprj_logic1[57] ,
    \mprj_logic1[56] ,
    \mprj_logic1[55] ,
    \mprj_logic1[54] ,
    \mprj_logic1[53] ,
    \mprj_logic1[52] ,
    \mprj_logic1[51] ,
    \mprj_logic1[50] ,
    \mprj_logic1[49] ,
    \mprj_logic1[48] ,
    \mprj_logic1[47] ,
    \mprj_logic1[46] ,
    \mprj_logic1[45] ,
    \mprj_logic1[44] ,
    \mprj_logic1[43] ,
    \mprj_logic1[42] ,
    \mprj_logic1[41] ,
    \mprj_logic1[40] ,
    \mprj_logic1[39] ,
    \mprj_logic1[38] ,
    \mprj_logic1[37] ,
    \mprj_logic1[36] ,
    \mprj_logic1[35] ,
    \mprj_logic1[34] ,
    \mprj_logic1[33] ,
    \mprj_logic1[32] ,
    \mprj_logic1[31] ,
    \mprj_logic1[30] ,
    \mprj_logic1[29] ,
    \mprj_logic1[28] ,
    \mprj_logic1[27] ,
    \mprj_logic1[26] ,
    \mprj_logic1[25] ,
    \mprj_logic1[24] ,
    \mprj_logic1[23] ,
    \mprj_logic1[22] ,
    \mprj_logic1[21] ,
    \mprj_logic1[20] ,
    \mprj_logic1[19] ,
    \mprj_logic1[18] ,
    \mprj_logic1[17] ,
    \mprj_logic1[16] ,
    \mprj_logic1[15] ,
    \mprj_logic1[14] ,
    \mprj_logic1[13] ,
    \mprj_logic1[12] ,
    \mprj_logic1[11] ,
    \mprj_logic1[10] ,
    \mprj_logic1[9] ,
    \mprj_logic1[8] ,
    \mprj_logic1[7] ,
    \mprj_logic1[6] ,
    \mprj_logic1[5] ,
    \mprj_logic1[4] ,
    \mprj_logic1[3] ,
    \mprj_logic1[2] ,
    \mprj_logic1[1] ,
    \mprj_logic1[0] }));
 mgmt_protect_hv powergood_check (.mprj2_vdd_logic1(net954),
    .mprj_vdd_logic1(net952));
 sky130_fd_sc_hd__nand2_1 \user_irq_gates[0]  (.A(user_irq_core[0]),
    .B(\user_irq_enable[0] ),
    .Y(\user_irq_bar[0] ));
 sky130_fd_sc_hd__nand2_1 \user_irq_gates[1]  (.A(user_irq_core[1]),
    .B(\user_irq_enable[1] ),
    .Y(\user_irq_bar[1] ));
 sky130_fd_sc_hd__nand2_1 \user_irq_gates[2]  (.A(user_irq_core[2]),
    .B(\user_irq_enable[2] ),
    .Y(\user_irq_bar[2] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[0]  (.A(la_data_out_core[0]),
    .B(\la_data_in_enable[0] ),
    .Y(\la_data_in_mprj_bar[0] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[100]  (.A(la_data_out_core[100]),
    .B(\la_data_in_enable[100] ),
    .Y(\la_data_in_mprj_bar[100] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[101]  (.A(la_data_out_core[101]),
    .B(\la_data_in_enable[101] ),
    .Y(\la_data_in_mprj_bar[101] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[102]  (.A(la_data_out_core[102]),
    .B(\la_data_in_enable[102] ),
    .Y(\la_data_in_mprj_bar[102] ));
 sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[103]  (.A(la_data_out_core[103]),
    .B(\la_data_in_enable[103] ),
    .Y(\la_data_in_mprj_bar[103] ));
 sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[104]  (.A(la_data_out_core[104]),
    .B(\la_data_in_enable[104] ),
    .Y(\la_data_in_mprj_bar[104] ));
 sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[105]  (.A(la_data_out_core[105]),
    .B(\la_data_in_enable[105] ),
    .Y(\la_data_in_mprj_bar[105] ));
 sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[106]  (.A(la_data_out_core[106]),
    .B(\la_data_in_enable[106] ),
    .Y(\la_data_in_mprj_bar[106] ));
 sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[107]  (.A(la_data_out_core[107]),
    .B(\la_data_in_enable[107] ),
    .Y(\la_data_in_mprj_bar[107] ));
 sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[108]  (.A(la_data_out_core[108]),
    .B(\la_data_in_enable[108] ),
    .Y(\la_data_in_mprj_bar[108] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[109]  (.A(la_data_out_core[109]),
    .B(\la_data_in_enable[109] ),
    .Y(\la_data_in_mprj_bar[109] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[10]  (.A(la_data_out_core[10]),
    .B(\la_data_in_enable[10] ),
    .Y(\la_data_in_mprj_bar[10] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[110]  (.A(la_data_out_core[110]),
    .B(\la_data_in_enable[110] ),
    .Y(\la_data_in_mprj_bar[110] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[111]  (.A(la_data_out_core[111]),
    .B(\la_data_in_enable[111] ),
    .Y(\la_data_in_mprj_bar[111] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[112]  (.A(la_data_out_core[112]),
    .B(\la_data_in_enable[112] ),
    .Y(\la_data_in_mprj_bar[112] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[113]  (.A(la_data_out_core[113]),
    .B(\la_data_in_enable[113] ),
    .Y(\la_data_in_mprj_bar[113] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[114]  (.A(la_data_out_core[114]),
    .B(\la_data_in_enable[114] ),
    .Y(\la_data_in_mprj_bar[114] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[115]  (.A(la_data_out_core[115]),
    .B(\la_data_in_enable[115] ),
    .Y(\la_data_in_mprj_bar[115] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[116]  (.A(la_data_out_core[116]),
    .B(\la_data_in_enable[116] ),
    .Y(\la_data_in_mprj_bar[116] ));
 sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[117]  (.A(la_data_out_core[117]),
    .B(\la_data_in_enable[117] ),
    .Y(\la_data_in_mprj_bar[117] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[118]  (.A(la_data_out_core[118]),
    .B(\la_data_in_enable[118] ),
    .Y(\la_data_in_mprj_bar[118] ));
 sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[119]  (.A(la_data_out_core[119]),
    .B(\la_data_in_enable[119] ),
    .Y(\la_data_in_mprj_bar[119] ));
 sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[11]  (.A(la_data_out_core[11]),
    .B(\la_data_in_enable[11] ),
    .Y(\la_data_in_mprj_bar[11] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[120]  (.A(la_data_out_core[120]),
    .B(\la_data_in_enable[120] ),
    .Y(\la_data_in_mprj_bar[120] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[121]  (.A(la_data_out_core[121]),
    .B(\la_data_in_enable[121] ),
    .Y(\la_data_in_mprj_bar[121] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[122]  (.A(la_data_out_core[122]),
    .B(\la_data_in_enable[122] ),
    .Y(\la_data_in_mprj_bar[122] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[123]  (.A(la_data_out_core[123]),
    .B(\la_data_in_enable[123] ),
    .Y(\la_data_in_mprj_bar[123] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[124]  (.A(la_data_out_core[124]),
    .B(\la_data_in_enable[124] ),
    .Y(\la_data_in_mprj_bar[124] ));
 sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[125]  (.A(la_data_out_core[125]),
    .B(\la_data_in_enable[125] ),
    .Y(\la_data_in_mprj_bar[125] ));
 sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[126]  (.A(la_data_out_core[126]),
    .B(\la_data_in_enable[126] ),
    .Y(\la_data_in_mprj_bar[126] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[127]  (.A(la_data_out_core[127]),
    .B(\la_data_in_enable[127] ),
    .Y(\la_data_in_mprj_bar[127] ));
 sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[12]  (.A(la_data_out_core[12]),
    .B(\la_data_in_enable[12] ),
    .Y(\la_data_in_mprj_bar[12] ));
 sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[13]  (.A(la_data_out_core[13]),
    .B(\la_data_in_enable[13] ),
    .Y(\la_data_in_mprj_bar[13] ));
 sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[14]  (.A(la_data_out_core[14]),
    .B(\la_data_in_enable[14] ),
    .Y(\la_data_in_mprj_bar[14] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[15]  (.A(la_data_out_core[15]),
    .B(\la_data_in_enable[15] ),
    .Y(\la_data_in_mprj_bar[15] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[16]  (.A(la_data_out_core[16]),
    .B(\la_data_in_enable[16] ),
    .Y(\la_data_in_mprj_bar[16] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[17]  (.A(la_data_out_core[17]),
    .B(\la_data_in_enable[17] ),
    .Y(\la_data_in_mprj_bar[17] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[18]  (.A(la_data_out_core[18]),
    .B(\la_data_in_enable[18] ),
    .Y(\la_data_in_mprj_bar[18] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[19]  (.A(la_data_out_core[19]),
    .B(\la_data_in_enable[19] ),
    .Y(\la_data_in_mprj_bar[19] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[1]  (.A(la_data_out_core[1]),
    .B(\la_data_in_enable[1] ),
    .Y(\la_data_in_mprj_bar[1] ));
 sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[20]  (.A(la_data_out_core[20]),
    .B(\la_data_in_enable[20] ),
    .Y(\la_data_in_mprj_bar[20] ));
 sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[21]  (.A(la_data_out_core[21]),
    .B(\la_data_in_enable[21] ),
    .Y(\la_data_in_mprj_bar[21] ));
 sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[22]  (.A(la_data_out_core[22]),
    .B(\la_data_in_enable[22] ),
    .Y(\la_data_in_mprj_bar[22] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[23]  (.A(la_data_out_core[23]),
    .B(\la_data_in_enable[23] ),
    .Y(\la_data_in_mprj_bar[23] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[24]  (.A(la_data_out_core[24]),
    .B(\la_data_in_enable[24] ),
    .Y(\la_data_in_mprj_bar[24] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[25]  (.A(la_data_out_core[25]),
    .B(\la_data_in_enable[25] ),
    .Y(\la_data_in_mprj_bar[25] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[26]  (.A(la_data_out_core[26]),
    .B(\la_data_in_enable[26] ),
    .Y(\la_data_in_mprj_bar[26] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[27]  (.A(la_data_out_core[27]),
    .B(\la_data_in_enable[27] ),
    .Y(\la_data_in_mprj_bar[27] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[28]  (.A(la_data_out_core[28]),
    .B(\la_data_in_enable[28] ),
    .Y(\la_data_in_mprj_bar[28] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[29]  (.A(la_data_out_core[29]),
    .B(\la_data_in_enable[29] ),
    .Y(\la_data_in_mprj_bar[29] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[2]  (.A(la_data_out_core[2]),
    .B(\la_data_in_enable[2] ),
    .Y(\la_data_in_mprj_bar[2] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[30]  (.A(la_data_out_core[30]),
    .B(\la_data_in_enable[30] ),
    .Y(\la_data_in_mprj_bar[30] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[31]  (.A(la_data_out_core[31]),
    .B(\la_data_in_enable[31] ),
    .Y(\la_data_in_mprj_bar[31] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[32]  (.A(la_data_out_core[32]),
    .B(\la_data_in_enable[32] ),
    .Y(\la_data_in_mprj_bar[32] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[33]  (.A(la_data_out_core[33]),
    .B(\la_data_in_enable[33] ),
    .Y(\la_data_in_mprj_bar[33] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[34]  (.A(la_data_out_core[34]),
    .B(\la_data_in_enable[34] ),
    .Y(\la_data_in_mprj_bar[34] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[35]  (.A(la_data_out_core[35]),
    .B(\la_data_in_enable[35] ),
    .Y(\la_data_in_mprj_bar[35] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[36]  (.A(la_data_out_core[36]),
    .B(\la_data_in_enable[36] ),
    .Y(\la_data_in_mprj_bar[36] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[37]  (.A(la_data_out_core[37]),
    .B(\la_data_in_enable[37] ),
    .Y(\la_data_in_mprj_bar[37] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[38]  (.A(la_data_out_core[38]),
    .B(\la_data_in_enable[38] ),
    .Y(\la_data_in_mprj_bar[38] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[39]  (.A(la_data_out_core[39]),
    .B(\la_data_in_enable[39] ),
    .Y(\la_data_in_mprj_bar[39] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[3]  (.A(la_data_out_core[3]),
    .B(\la_data_in_enable[3] ),
    .Y(\la_data_in_mprj_bar[3] ));
 sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[40]  (.A(la_data_out_core[40]),
    .B(\la_data_in_enable[40] ),
    .Y(\la_data_in_mprj_bar[40] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[41]  (.A(la_data_out_core[41]),
    .B(\la_data_in_enable[41] ),
    .Y(\la_data_in_mprj_bar[41] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[42]  (.A(la_data_out_core[42]),
    .B(\la_data_in_enable[42] ),
    .Y(\la_data_in_mprj_bar[42] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[43]  (.A(la_data_out_core[43]),
    .B(\la_data_in_enable[43] ),
    .Y(\la_data_in_mprj_bar[43] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[44]  (.A(la_data_out_core[44]),
    .B(\la_data_in_enable[44] ),
    .Y(\la_data_in_mprj_bar[44] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[45]  (.A(la_data_out_core[45]),
    .B(\la_data_in_enable[45] ),
    .Y(\la_data_in_mprj_bar[45] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[46]  (.A(la_data_out_core[46]),
    .B(\la_data_in_enable[46] ),
    .Y(\la_data_in_mprj_bar[46] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[47]  (.A(la_data_out_core[47]),
    .B(\la_data_in_enable[47] ),
    .Y(\la_data_in_mprj_bar[47] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[48]  (.A(la_data_out_core[48]),
    .B(\la_data_in_enable[48] ),
    .Y(\la_data_in_mprj_bar[48] ));
 sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[49]  (.A(la_data_out_core[49]),
    .B(\la_data_in_enable[49] ),
    .Y(\la_data_in_mprj_bar[49] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[4]  (.A(la_data_out_core[4]),
    .B(\la_data_in_enable[4] ),
    .Y(\la_data_in_mprj_bar[4] ));
 sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[50]  (.A(la_data_out_core[50]),
    .B(\la_data_in_enable[50] ),
    .Y(\la_data_in_mprj_bar[50] ));
 sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[51]  (.A(la_data_out_core[51]),
    .B(\la_data_in_enable[51] ),
    .Y(\la_data_in_mprj_bar[51] ));
 sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[52]  (.A(la_data_out_core[52]),
    .B(\la_data_in_enable[52] ),
    .Y(\la_data_in_mprj_bar[52] ));
 sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[53]  (.A(la_data_out_core[53]),
    .B(\la_data_in_enable[53] ),
    .Y(\la_data_in_mprj_bar[53] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[54]  (.A(la_data_out_core[54]),
    .B(\la_data_in_enable[54] ),
    .Y(\la_data_in_mprj_bar[54] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[55]  (.A(la_data_out_core[55]),
    .B(\la_data_in_enable[55] ),
    .Y(\la_data_in_mprj_bar[55] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[56]  (.A(la_data_out_core[56]),
    .B(\la_data_in_enable[56] ),
    .Y(\la_data_in_mprj_bar[56] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[57]  (.A(la_data_out_core[57]),
    .B(\la_data_in_enable[57] ),
    .Y(\la_data_in_mprj_bar[57] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[58]  (.A(la_data_out_core[58]),
    .B(\la_data_in_enable[58] ),
    .Y(\la_data_in_mprj_bar[58] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[59]  (.A(la_data_out_core[59]),
    .B(\la_data_in_enable[59] ),
    .Y(\la_data_in_mprj_bar[59] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[5]  (.A(la_data_out_core[5]),
    .B(\la_data_in_enable[5] ),
    .Y(\la_data_in_mprj_bar[5] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[60]  (.A(la_data_out_core[60]),
    .B(\la_data_in_enable[60] ),
    .Y(\la_data_in_mprj_bar[60] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[61]  (.A(la_data_out_core[61]),
    .B(\la_data_in_enable[61] ),
    .Y(\la_data_in_mprj_bar[61] ));
 sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[62]  (.A(la_data_out_core[62]),
    .B(\la_data_in_enable[62] ),
    .Y(\la_data_in_mprj_bar[62] ));
 sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[63]  (.A(la_data_out_core[63]),
    .B(\la_data_in_enable[63] ),
    .Y(\la_data_in_mprj_bar[63] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[64]  (.A(la_data_out_core[64]),
    .B(\la_data_in_enable[64] ),
    .Y(\la_data_in_mprj_bar[64] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[65]  (.A(la_data_out_core[65]),
    .B(\la_data_in_enable[65] ),
    .Y(\la_data_in_mprj_bar[65] ));
 sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[66]  (.A(la_data_out_core[66]),
    .B(\la_data_in_enable[66] ),
    .Y(\la_data_in_mprj_bar[66] ));
 sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[67]  (.A(la_data_out_core[67]),
    .B(\la_data_in_enable[67] ),
    .Y(\la_data_in_mprj_bar[67] ));
 sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[68]  (.A(la_data_out_core[68]),
    .B(\la_data_in_enable[68] ),
    .Y(\la_data_in_mprj_bar[68] ));
 sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[69]  (.A(la_data_out_core[69]),
    .B(\la_data_in_enable[69] ),
    .Y(\la_data_in_mprj_bar[69] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[6]  (.A(la_data_out_core[6]),
    .B(\la_data_in_enable[6] ),
    .Y(\la_data_in_mprj_bar[6] ));
 sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[70]  (.A(la_data_out_core[70]),
    .B(\la_data_in_enable[70] ),
    .Y(\la_data_in_mprj_bar[70] ));
 sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[71]  (.A(la_data_out_core[71]),
    .B(\la_data_in_enable[71] ),
    .Y(\la_data_in_mprj_bar[71] ));
 sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[72]  (.A(la_data_out_core[72]),
    .B(\la_data_in_enable[72] ),
    .Y(\la_data_in_mprj_bar[72] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[73]  (.A(la_data_out_core[73]),
    .B(\la_data_in_enable[73] ),
    .Y(\la_data_in_mprj_bar[73] ));
 sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[74]  (.A(la_data_out_core[74]),
    .B(\la_data_in_enable[74] ),
    .Y(\la_data_in_mprj_bar[74] ));
 sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[75]  (.A(la_data_out_core[75]),
    .B(\la_data_in_enable[75] ),
    .Y(\la_data_in_mprj_bar[75] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[76]  (.A(la_data_out_core[76]),
    .B(\la_data_in_enable[76] ),
    .Y(\la_data_in_mprj_bar[76] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[77]  (.A(la_data_out_core[77]),
    .B(\la_data_in_enable[77] ),
    .Y(\la_data_in_mprj_bar[77] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[78]  (.A(la_data_out_core[78]),
    .B(\la_data_in_enable[78] ),
    .Y(\la_data_in_mprj_bar[78] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[79]  (.A(la_data_out_core[79]),
    .B(\la_data_in_enable[79] ),
    .Y(\la_data_in_mprj_bar[79] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[7]  (.A(la_data_out_core[7]),
    .B(\la_data_in_enable[7] ),
    .Y(\la_data_in_mprj_bar[7] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[80]  (.A(la_data_out_core[80]),
    .B(\la_data_in_enable[80] ),
    .Y(\la_data_in_mprj_bar[80] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[81]  (.A(la_data_out_core[81]),
    .B(\la_data_in_enable[81] ),
    .Y(\la_data_in_mprj_bar[81] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[82]  (.A(la_data_out_core[82]),
    .B(\la_data_in_enable[82] ),
    .Y(\la_data_in_mprj_bar[82] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[83]  (.A(la_data_out_core[83]),
    .B(\la_data_in_enable[83] ),
    .Y(\la_data_in_mprj_bar[83] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[84]  (.A(la_data_out_core[84]),
    .B(\la_data_in_enable[84] ),
    .Y(\la_data_in_mprj_bar[84] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[85]  (.A(la_data_out_core[85]),
    .B(\la_data_in_enable[85] ),
    .Y(\la_data_in_mprj_bar[85] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[86]  (.A(la_data_out_core[86]),
    .B(\la_data_in_enable[86] ),
    .Y(\la_data_in_mprj_bar[86] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[87]  (.A(la_data_out_core[87]),
    .B(\la_data_in_enable[87] ),
    .Y(\la_data_in_mprj_bar[87] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[88]  (.A(la_data_out_core[88]),
    .B(\la_data_in_enable[88] ),
    .Y(\la_data_in_mprj_bar[88] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[89]  (.A(la_data_out_core[89]),
    .B(\la_data_in_enable[89] ),
    .Y(\la_data_in_mprj_bar[89] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[8]  (.A(la_data_out_core[8]),
    .B(\la_data_in_enable[8] ),
    .Y(\la_data_in_mprj_bar[8] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[90]  (.A(la_data_out_core[90]),
    .B(\la_data_in_enable[90] ),
    .Y(\la_data_in_mprj_bar[90] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[91]  (.A(la_data_out_core[91]),
    .B(\la_data_in_enable[91] ),
    .Y(\la_data_in_mprj_bar[91] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[92]  (.A(la_data_out_core[92]),
    .B(\la_data_in_enable[92] ),
    .Y(\la_data_in_mprj_bar[92] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[93]  (.A(la_data_out_core[93]),
    .B(\la_data_in_enable[93] ),
    .Y(\la_data_in_mprj_bar[93] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[94]  (.A(la_data_out_core[94]),
    .B(\la_data_in_enable[94] ),
    .Y(\la_data_in_mprj_bar[94] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[95]  (.A(la_data_out_core[95]),
    .B(\la_data_in_enable[95] ),
    .Y(\la_data_in_mprj_bar[95] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[96]  (.A(la_data_out_core[96]),
    .B(\la_data_in_enable[96] ),
    .Y(\la_data_in_mprj_bar[96] ));
 sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[97]  (.A(la_data_out_core[97]),
    .B(\la_data_in_enable[97] ),
    .Y(\la_data_in_mprj_bar[97] ));
 sky130_fd_sc_hd__nand2_4 \user_to_mprj_in_gates[98]  (.A(la_data_out_core[98]),
    .B(\la_data_in_enable[98] ),
    .Y(\la_data_in_mprj_bar[98] ));
 sky130_fd_sc_hd__nand2_8 \user_to_mprj_in_gates[99]  (.A(la_data_out_core[99]),
    .B(\la_data_in_enable[99] ),
    .Y(\la_data_in_mprj_bar[99] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[9]  (.A(la_data_out_core[9]),
    .B(\la_data_in_enable[9] ),
    .Y(\la_data_in_mprj_bar[9] ));
 sky130_fd_sc_hd__nand2_1 user_wb_ack_gate (.A(mprj_ack_i_user),
    .B(wb_in_enable),
    .Y(mprj_ack_i_core_bar));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[0]  (.A(mprj_dat_i_user[0]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[0] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[10]  (.A(mprj_dat_i_user[10]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[10] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[11]  (.A(mprj_dat_i_user[11]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[11] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[12]  (.A(mprj_dat_i_user[12]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[12] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[13]  (.A(mprj_dat_i_user[13]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[13] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[14]  (.A(mprj_dat_i_user[14]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[14] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[15]  (.A(mprj_dat_i_user[15]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[15] ));
 sky130_fd_sc_hd__nand2_2 \user_wb_dat_gates[16]  (.A(mprj_dat_i_user[16]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[16] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[17]  (.A(mprj_dat_i_user[17]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[17] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[18]  (.A(mprj_dat_i_user[18]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[18] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[19]  (.A(mprj_dat_i_user[19]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[19] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[1]  (.A(mprj_dat_i_user[1]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[1] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[20]  (.A(mprj_dat_i_user[20]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[20] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[21]  (.A(mprj_dat_i_user[21]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[21] ));
 sky130_fd_sc_hd__nand2_2 \user_wb_dat_gates[22]  (.A(mprj_dat_i_user[22]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[22] ));
 sky130_fd_sc_hd__nand2_2 \user_wb_dat_gates[23]  (.A(mprj_dat_i_user[23]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[23] ));
 sky130_fd_sc_hd__nand2_2 \user_wb_dat_gates[24]  (.A(mprj_dat_i_user[24]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[24] ));
 sky130_fd_sc_hd__nand2_2 \user_wb_dat_gates[25]  (.A(mprj_dat_i_user[25]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[25] ));
 sky130_fd_sc_hd__nand2_2 \user_wb_dat_gates[26]  (.A(mprj_dat_i_user[26]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[26] ));
 sky130_fd_sc_hd__nand2_2 \user_wb_dat_gates[27]  (.A(mprj_dat_i_user[27]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[27] ));
 sky130_fd_sc_hd__nand2_2 \user_wb_dat_gates[28]  (.A(mprj_dat_i_user[28]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[28] ));
 sky130_fd_sc_hd__nand2_2 \user_wb_dat_gates[29]  (.A(mprj_dat_i_user[29]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[29] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[2]  (.A(mprj_dat_i_user[2]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[2] ));
 sky130_fd_sc_hd__nand2_2 \user_wb_dat_gates[30]  (.A(mprj_dat_i_user[30]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[30] ));
 sky130_fd_sc_hd__nand2_2 \user_wb_dat_gates[31]  (.A(mprj_dat_i_user[31]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[31] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[3]  (.A(mprj_dat_i_user[3]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[3] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[4]  (.A(mprj_dat_i_user[4]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[4] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[5]  (.A(mprj_dat_i_user[5]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[5] ));
 sky130_fd_sc_hd__nand2_2 \user_wb_dat_gates[6]  (.A(mprj_dat_i_user[6]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[6] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[7]  (.A(mprj_dat_i_user[7]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[7] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[8]  (.A(mprj_dat_i_user[8]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[8] ));
 sky130_fd_sc_hd__nand2_2 \user_wb_dat_gates[9]  (.A(mprj_dat_i_user[9]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[9] ));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__clkbuf_4 input2 (.A(caravel_clk2),
    .X(net2));
 sky130_fd_sc_hd__buf_8 input1 (.A(caravel_clk),
    .X(net1));
 sky130_fd_sc_hd__buf_8 input3 (.A(caravel_rstn),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_4 input4 (.A(la_data_out_mprj[0]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_4 input5 (.A(la_data_out_mprj[100]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(la_data_out_mprj[101]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_4 input7 (.A(la_data_out_mprj[102]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_4 input8 (.A(la_data_out_mprj[103]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_4 input9 (.A(la_data_out_mprj[104]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_4 input10 (.A(la_data_out_mprj[105]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 input11 (.A(la_data_out_mprj[106]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 input12 (.A(la_data_out_mprj[107]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 input13 (.A(la_data_out_mprj[108]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_4 input14 (.A(la_data_out_mprj[109]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_4 input15 (.A(la_data_out_mprj[10]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_4 input16 (.A(la_data_out_mprj[110]),
    .X(net16));
 sky130_fd_sc_hd__buf_4 input17 (.A(la_data_out_mprj[111]),
    .X(net17));
 sky130_fd_sc_hd__buf_6 input18 (.A(la_data_out_mprj[112]),
    .X(net18));
 sky130_fd_sc_hd__buf_4 input19 (.A(la_data_out_mprj[113]),
    .X(net19));
 sky130_fd_sc_hd__buf_6 input20 (.A(la_data_out_mprj[114]),
    .X(net20));
 sky130_fd_sc_hd__buf_4 input21 (.A(la_data_out_mprj[115]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_4 input22 (.A(la_data_out_mprj[116]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_4 input23 (.A(la_data_out_mprj[117]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_4 input24 (.A(la_data_out_mprj[118]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_4 input25 (.A(la_data_out_mprj[119]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_4 input26 (.A(la_data_out_mprj[11]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_4 input27 (.A(la_data_out_mprj[120]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_4 input28 (.A(la_data_out_mprj[121]),
    .X(net28));
 sky130_fd_sc_hd__buf_4 input29 (.A(la_data_out_mprj[122]),
    .X(net29));
 sky130_fd_sc_hd__buf_4 input30 (.A(la_data_out_mprj[123]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_8 input31 (.A(la_data_out_mprj[124]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_8 input32 (.A(la_data_out_mprj[125]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_8 input33 (.A(la_data_out_mprj[126]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_8 input34 (.A(la_data_out_mprj[127]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_4 input35 (.A(la_data_out_mprj[12]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_4 input36 (.A(la_data_out_mprj[13]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_4 input37 (.A(la_data_out_mprj[14]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_4 input38 (.A(la_data_out_mprj[15]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_4 input39 (.A(la_data_out_mprj[16]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_4 input40 (.A(la_data_out_mprj[17]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_4 input41 (.A(la_data_out_mprj[18]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_4 input42 (.A(la_data_out_mprj[19]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_4 input43 (.A(la_data_out_mprj[1]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_4 input44 (.A(la_data_out_mprj[20]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_4 input45 (.A(la_data_out_mprj[21]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_4 input46 (.A(la_data_out_mprj[22]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_4 input47 (.A(la_data_out_mprj[23]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_4 input48 (.A(la_data_out_mprj[24]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_4 input49 (.A(la_data_out_mprj[25]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_4 input50 (.A(la_data_out_mprj[26]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_4 input51 (.A(la_data_out_mprj[27]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_4 input52 (.A(la_data_out_mprj[28]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_4 input53 (.A(la_data_out_mprj[29]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_4 input54 (.A(la_data_out_mprj[2]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_4 input55 (.A(la_data_out_mprj[30]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_4 input56 (.A(la_data_out_mprj[31]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_4 input57 (.A(la_data_out_mprj[32]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_4 input58 (.A(la_data_out_mprj[33]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_4 input59 (.A(la_data_out_mprj[34]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_4 input60 (.A(la_data_out_mprj[35]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_4 input61 (.A(la_data_out_mprj[36]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_4 input62 (.A(la_data_out_mprj[37]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_4 input63 (.A(la_data_out_mprj[38]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_4 input64 (.A(la_data_out_mprj[39]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_4 input65 (.A(la_data_out_mprj[3]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_4 input66 (.A(la_data_out_mprj[40]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_4 input67 (.A(la_data_out_mprj[41]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_4 input68 (.A(la_data_out_mprj[42]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_4 input69 (.A(la_data_out_mprj[43]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_4 input70 (.A(la_data_out_mprj[44]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_4 input71 (.A(la_data_out_mprj[45]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_4 input72 (.A(la_data_out_mprj[46]),
    .X(net72));
 sky130_fd_sc_hd__buf_4 input73 (.A(la_data_out_mprj[47]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_4 input74 (.A(la_data_out_mprj[48]),
    .X(net74));
 sky130_fd_sc_hd__buf_4 input75 (.A(la_data_out_mprj[49]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_4 input76 (.A(la_data_out_mprj[4]),
    .X(net76));
 sky130_fd_sc_hd__buf_4 input77 (.A(la_data_out_mprj[50]),
    .X(net77));
 sky130_fd_sc_hd__buf_4 input78 (.A(la_data_out_mprj[51]),
    .X(net78));
 sky130_fd_sc_hd__buf_4 input79 (.A(la_data_out_mprj[52]),
    .X(net79));
 sky130_fd_sc_hd__buf_4 input80 (.A(la_data_out_mprj[53]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_4 input81 (.A(la_data_out_mprj[54]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_4 input82 (.A(la_data_out_mprj[55]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_4 input83 (.A(la_data_out_mprj[56]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_4 input84 (.A(la_data_out_mprj[57]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_4 input85 (.A(la_data_out_mprj[58]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_4 input86 (.A(la_data_out_mprj[59]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_4 input87 (.A(la_data_out_mprj[5]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_4 input88 (.A(la_data_out_mprj[60]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_4 input89 (.A(la_data_out_mprj[61]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_4 input90 (.A(la_data_out_mprj[62]),
    .X(net90));
 sky130_fd_sc_hd__buf_4 input91 (.A(la_data_out_mprj[63]),
    .X(net91));
 sky130_fd_sc_hd__buf_4 input92 (.A(la_data_out_mprj[64]),
    .X(net92));
 sky130_fd_sc_hd__buf_6 input93 (.A(la_data_out_mprj[65]),
    .X(net93));
 sky130_fd_sc_hd__buf_6 input94 (.A(la_data_out_mprj[66]),
    .X(net94));
 sky130_fd_sc_hd__buf_6 input95 (.A(la_data_out_mprj[67]),
    .X(net95));
 sky130_fd_sc_hd__buf_6 input96 (.A(la_data_out_mprj[68]),
    .X(net96));
 sky130_fd_sc_hd__buf_6 input97 (.A(la_data_out_mprj[69]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_4 input98 (.A(la_data_out_mprj[6]),
    .X(net98));
 sky130_fd_sc_hd__buf_6 input99 (.A(la_data_out_mprj[70]),
    .X(net99));
 sky130_fd_sc_hd__buf_6 input100 (.A(la_data_out_mprj[71]),
    .X(net100));
 sky130_fd_sc_hd__buf_4 input101 (.A(la_data_out_mprj[72]),
    .X(net101));
 sky130_fd_sc_hd__buf_4 input102 (.A(la_data_out_mprj[73]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_4 input103 (.A(la_data_out_mprj[74]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_4 input104 (.A(la_data_out_mprj[75]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_4 input105 (.A(la_data_out_mprj[76]),
    .X(net105));
 sky130_fd_sc_hd__buf_4 input106 (.A(la_data_out_mprj[77]),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_4 input107 (.A(la_data_out_mprj[78]),
    .X(net107));
 sky130_fd_sc_hd__buf_4 input108 (.A(la_data_out_mprj[79]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_4 input109 (.A(la_data_out_mprj[7]),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_8 input110 (.A(la_data_out_mprj[80]),
    .X(net110));
 sky130_fd_sc_hd__buf_6 input111 (.A(la_data_out_mprj[81]),
    .X(net111));
 sky130_fd_sc_hd__buf_6 input112 (.A(la_data_out_mprj[82]),
    .X(net112));
 sky130_fd_sc_hd__buf_6 input113 (.A(la_data_out_mprj[83]),
    .X(net113));
 sky130_fd_sc_hd__buf_8 input114 (.A(la_data_out_mprj[84]),
    .X(net114));
 sky130_fd_sc_hd__buf_8 input115 (.A(la_data_out_mprj[85]),
    .X(net115));
 sky130_fd_sc_hd__buf_8 input116 (.A(la_data_out_mprj[86]),
    .X(net116));
 sky130_fd_sc_hd__buf_8 input117 (.A(la_data_out_mprj[87]),
    .X(net117));
 sky130_fd_sc_hd__buf_8 input118 (.A(la_data_out_mprj[88]),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_4 input119 (.A(la_data_out_mprj[89]),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_4 input120 (.A(la_data_out_mprj[8]),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_4 input121 (.A(la_data_out_mprj[90]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_4 input122 (.A(la_data_out_mprj[91]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_4 input123 (.A(la_data_out_mprj[92]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_4 input124 (.A(la_data_out_mprj[93]),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_4 input125 (.A(la_data_out_mprj[94]),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_4 input126 (.A(la_data_out_mprj[95]),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_4 input127 (.A(la_data_out_mprj[96]),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_4 input128 (.A(la_data_out_mprj[97]),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_4 input129 (.A(la_data_out_mprj[98]),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_4 input130 (.A(la_data_out_mprj[99]),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_4 input131 (.A(la_data_out_mprj[9]),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_4 input132 (.A(la_iena_mprj[0]),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_4 input133 (.A(la_iena_mprj[100]),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_4 input134 (.A(la_iena_mprj[101]),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_4 input135 (.A(la_iena_mprj[102]),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_4 input136 (.A(la_iena_mprj[103]),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_4 input137 (.A(la_iena_mprj[104]),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_4 input138 (.A(la_iena_mprj[105]),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_4 input139 (.A(la_iena_mprj[106]),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_4 input140 (.A(la_iena_mprj[107]),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_4 input141 (.A(la_iena_mprj[108]),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_4 input142 (.A(la_iena_mprj[109]),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_4 input143 (.A(la_iena_mprj[10]),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_4 input144 (.A(la_iena_mprj[110]),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_4 input145 (.A(la_iena_mprj[111]),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_4 input146 (.A(la_iena_mprj[112]),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_4 input147 (.A(la_iena_mprj[113]),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_4 input148 (.A(la_iena_mprj[114]),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_4 input149 (.A(la_iena_mprj[115]),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_4 input150 (.A(la_iena_mprj[116]),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_4 input151 (.A(la_iena_mprj[117]),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_4 input152 (.A(la_iena_mprj[118]),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_4 input153 (.A(la_iena_mprj[119]),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_4 input154 (.A(la_iena_mprj[11]),
    .X(net154));
 sky130_fd_sc_hd__buf_4 input155 (.A(la_iena_mprj[120]),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_4 input156 (.A(la_iena_mprj[121]),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_4 input157 (.A(la_iena_mprj[122]),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_4 input158 (.A(la_iena_mprj[123]),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_4 input159 (.A(la_iena_mprj[124]),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_4 input160 (.A(la_iena_mprj[125]),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_4 input161 (.A(la_iena_mprj[126]),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_4 input162 (.A(la_iena_mprj[127]),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_4 input163 (.A(la_iena_mprj[12]),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_4 input164 (.A(la_iena_mprj[13]),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_4 input165 (.A(la_iena_mprj[14]),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_4 input166 (.A(la_iena_mprj[15]),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_4 input167 (.A(la_iena_mprj[16]),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_4 input168 (.A(la_iena_mprj[17]),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_4 input169 (.A(la_iena_mprj[18]),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_4 input170 (.A(la_iena_mprj[19]),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_4 input171 (.A(la_iena_mprj[1]),
    .X(net171));
 sky130_fd_sc_hd__buf_4 input172 (.A(la_iena_mprj[20]),
    .X(net172));
 sky130_fd_sc_hd__buf_4 input173 (.A(la_iena_mprj[21]),
    .X(net173));
 sky130_fd_sc_hd__buf_4 input174 (.A(la_iena_mprj[22]),
    .X(net174));
 sky130_fd_sc_hd__buf_4 input175 (.A(la_iena_mprj[23]),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_4 input176 (.A(la_iena_mprj[24]),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_4 input177 (.A(la_iena_mprj[25]),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_4 input178 (.A(la_iena_mprj[26]),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_4 input179 (.A(la_iena_mprj[27]),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_4 input180 (.A(la_iena_mprj[28]),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_4 input181 (.A(la_iena_mprj[29]),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_4 input182 (.A(la_iena_mprj[2]),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_4 input183 (.A(la_iena_mprj[30]),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_4 input184 (.A(la_iena_mprj[31]),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_4 input185 (.A(la_iena_mprj[32]),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_4 input186 (.A(la_iena_mprj[33]),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_4 input187 (.A(la_iena_mprj[34]),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_4 input188 (.A(la_iena_mprj[35]),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_4 input189 (.A(la_iena_mprj[36]),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_4 input190 (.A(la_iena_mprj[37]),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_4 input191 (.A(la_iena_mprj[38]),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_4 input192 (.A(la_iena_mprj[39]),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_4 input193 (.A(la_iena_mprj[3]),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_4 input194 (.A(la_iena_mprj[40]),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_4 input195 (.A(la_iena_mprj[41]),
    .X(net195));
 sky130_fd_sc_hd__buf_4 input196 (.A(la_iena_mprj[42]),
    .X(net196));
 sky130_fd_sc_hd__buf_4 input197 (.A(la_iena_mprj[43]),
    .X(net197));
 sky130_fd_sc_hd__buf_4 input198 (.A(la_iena_mprj[44]),
    .X(net198));
 sky130_fd_sc_hd__buf_4 input199 (.A(la_iena_mprj[45]),
    .X(net199));
 sky130_fd_sc_hd__buf_4 input200 (.A(la_iena_mprj[46]),
    .X(net200));
 sky130_fd_sc_hd__buf_4 input201 (.A(la_iena_mprj[47]),
    .X(net201));
 sky130_fd_sc_hd__buf_4 input202 (.A(la_iena_mprj[48]),
    .X(net202));
 sky130_fd_sc_hd__buf_4 input203 (.A(la_iena_mprj[49]),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_4 input204 (.A(la_iena_mprj[4]),
    .X(net204));
 sky130_fd_sc_hd__buf_4 input205 (.A(la_iena_mprj[50]),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_4 input206 (.A(la_iena_mprj[51]),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_4 input207 (.A(la_iena_mprj[52]),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_4 input208 (.A(la_iena_mprj[53]),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_4 input209 (.A(la_iena_mprj[54]),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_4 input210 (.A(la_iena_mprj[55]),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_4 input211 (.A(la_iena_mprj[56]),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_4 input212 (.A(la_iena_mprj[57]),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_4 input213 (.A(la_iena_mprj[58]),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_4 input214 (.A(la_iena_mprj[59]),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_4 input215 (.A(la_iena_mprj[5]),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_4 input216 (.A(la_iena_mprj[60]),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_4 input217 (.A(la_iena_mprj[61]),
    .X(net217));
 sky130_fd_sc_hd__buf_4 input218 (.A(la_iena_mprj[62]),
    .X(net218));
 sky130_fd_sc_hd__buf_4 input219 (.A(la_iena_mprj[63]),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_4 input220 (.A(la_iena_mprj[64]),
    .X(net220));
 sky130_fd_sc_hd__buf_4 input221 (.A(la_iena_mprj[65]),
    .X(net221));
 sky130_fd_sc_hd__buf_4 input222 (.A(la_iena_mprj[66]),
    .X(net222));
 sky130_fd_sc_hd__buf_4 input223 (.A(la_iena_mprj[67]),
    .X(net223));
 sky130_fd_sc_hd__buf_4 input224 (.A(la_iena_mprj[68]),
    .X(net224));
 sky130_fd_sc_hd__buf_4 input225 (.A(la_iena_mprj[69]),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_4 input226 (.A(la_iena_mprj[6]),
    .X(net226));
 sky130_fd_sc_hd__buf_4 input227 (.A(la_iena_mprj[70]),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_4 input228 (.A(la_iena_mprj[71]),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_4 input229 (.A(la_iena_mprj[72]),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_4 input230 (.A(la_iena_mprj[73]),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_4 input231 (.A(la_iena_mprj[74]),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_4 input232 (.A(la_iena_mprj[75]),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_4 input233 (.A(la_iena_mprj[76]),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_4 input234 (.A(la_iena_mprj[77]),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_4 input235 (.A(la_iena_mprj[78]),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_4 input236 (.A(la_iena_mprj[79]),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_4 input237 (.A(la_iena_mprj[7]),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_4 input238 (.A(la_iena_mprj[80]),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_4 input239 (.A(la_iena_mprj[81]),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_4 input240 (.A(la_iena_mprj[82]),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_4 input241 (.A(la_iena_mprj[83]),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_4 input242 (.A(la_iena_mprj[84]),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_4 input243 (.A(la_iena_mprj[85]),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_4 input244 (.A(la_iena_mprj[86]),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_4 input245 (.A(la_iena_mprj[87]),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_4 input246 (.A(la_iena_mprj[88]),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_4 input247 (.A(la_iena_mprj[89]),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_4 input248 (.A(la_iena_mprj[8]),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_4 input249 (.A(la_iena_mprj[90]),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_4 input250 (.A(la_iena_mprj[91]),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_4 input251 (.A(la_iena_mprj[92]),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_4 input252 (.A(la_iena_mprj[93]),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_4 input253 (.A(la_iena_mprj[94]),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_4 input254 (.A(la_iena_mprj[95]),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_4 input255 (.A(la_iena_mprj[96]),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_4 input256 (.A(la_iena_mprj[97]),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_4 input257 (.A(la_iena_mprj[98]),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_4 input258 (.A(la_iena_mprj[99]),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_4 input259 (.A(la_iena_mprj[9]),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_4 input260 (.A(la_oenb_mprj[0]),
    .X(net260));
 sky130_fd_sc_hd__buf_6 input261 (.A(la_oenb_mprj[100]),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_8 input262 (.A(la_oenb_mprj[101]),
    .X(net262));
 sky130_fd_sc_hd__buf_6 input263 (.A(la_oenb_mprj[102]),
    .X(net263));
 sky130_fd_sc_hd__buf_6 input264 (.A(la_oenb_mprj[103]),
    .X(net264));
 sky130_fd_sc_hd__buf_6 input265 (.A(la_oenb_mprj[104]),
    .X(net265));
 sky130_fd_sc_hd__buf_6 input266 (.A(la_oenb_mprj[105]),
    .X(net266));
 sky130_fd_sc_hd__buf_6 input267 (.A(la_oenb_mprj[106]),
    .X(net267));
 sky130_fd_sc_hd__buf_6 input268 (.A(la_oenb_mprj[107]),
    .X(net268));
 sky130_fd_sc_hd__buf_6 input269 (.A(la_oenb_mprj[108]),
    .X(net269));
 sky130_fd_sc_hd__buf_6 input270 (.A(la_oenb_mprj[109]),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_4 input271 (.A(la_oenb_mprj[10]),
    .X(net271));
 sky130_fd_sc_hd__buf_6 input272 (.A(la_oenb_mprj[110]),
    .X(net272));
 sky130_fd_sc_hd__buf_6 input273 (.A(la_oenb_mprj[111]),
    .X(net273));
 sky130_fd_sc_hd__buf_6 input274 (.A(la_oenb_mprj[112]),
    .X(net274));
 sky130_fd_sc_hd__buf_6 input275 (.A(la_oenb_mprj[113]),
    .X(net275));
 sky130_fd_sc_hd__buf_6 input276 (.A(la_oenb_mprj[114]),
    .X(net276));
 sky130_fd_sc_hd__buf_6 input277 (.A(la_oenb_mprj[115]),
    .X(net277));
 sky130_fd_sc_hd__buf_6 input278 (.A(la_oenb_mprj[116]),
    .X(net278));
 sky130_fd_sc_hd__buf_6 input279 (.A(la_oenb_mprj[117]),
    .X(net279));
 sky130_fd_sc_hd__buf_6 input280 (.A(la_oenb_mprj[118]),
    .X(net280));
 sky130_fd_sc_hd__buf_6 input281 (.A(la_oenb_mprj[119]),
    .X(net281));
 sky130_fd_sc_hd__clkbuf_4 input282 (.A(la_oenb_mprj[11]),
    .X(net282));
 sky130_fd_sc_hd__buf_6 input283 (.A(la_oenb_mprj[120]),
    .X(net283));
 sky130_fd_sc_hd__buf_6 input284 (.A(la_oenb_mprj[121]),
    .X(net284));
 sky130_fd_sc_hd__buf_6 input285 (.A(la_oenb_mprj[122]),
    .X(net285));
 sky130_fd_sc_hd__buf_6 input286 (.A(la_oenb_mprj[123]),
    .X(net286));
 sky130_fd_sc_hd__buf_6 input287 (.A(la_oenb_mprj[124]),
    .X(net287));
 sky130_fd_sc_hd__buf_6 input288 (.A(la_oenb_mprj[125]),
    .X(net288));
 sky130_fd_sc_hd__buf_6 input289 (.A(la_oenb_mprj[126]),
    .X(net289));
 sky130_fd_sc_hd__buf_6 input290 (.A(la_oenb_mprj[127]),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_4 input291 (.A(la_oenb_mprj[12]),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_4 input292 (.A(la_oenb_mprj[13]),
    .X(net292));
 sky130_fd_sc_hd__clkbuf_4 input293 (.A(la_oenb_mprj[14]),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_4 input294 (.A(la_oenb_mprj[15]),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_4 input295 (.A(la_oenb_mprj[16]),
    .X(net295));
 sky130_fd_sc_hd__clkbuf_4 input296 (.A(la_oenb_mprj[17]),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_4 input297 (.A(la_oenb_mprj[18]),
    .X(net297));
 sky130_fd_sc_hd__clkbuf_4 input298 (.A(la_oenb_mprj[19]),
    .X(net298));
 sky130_fd_sc_hd__clkbuf_4 input299 (.A(la_oenb_mprj[1]),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_4 input300 (.A(la_oenb_mprj[20]),
    .X(net300));
 sky130_fd_sc_hd__buf_6 input301 (.A(la_oenb_mprj[21]),
    .X(net301));
 sky130_fd_sc_hd__buf_4 input302 (.A(la_oenb_mprj[22]),
    .X(net302));
 sky130_fd_sc_hd__clkbuf_4 input303 (.A(la_oenb_mprj[23]),
    .X(net303));
 sky130_fd_sc_hd__buf_4 input304 (.A(la_oenb_mprj[24]),
    .X(net304));
 sky130_fd_sc_hd__buf_4 input305 (.A(la_oenb_mprj[25]),
    .X(net305));
 sky130_fd_sc_hd__buf_4 input306 (.A(la_oenb_mprj[26]),
    .X(net306));
 sky130_fd_sc_hd__buf_6 input307 (.A(la_oenb_mprj[27]),
    .X(net307));
 sky130_fd_sc_hd__clkbuf_8 input308 (.A(la_oenb_mprj[28]),
    .X(net308));
 sky130_fd_sc_hd__buf_6 input309 (.A(la_oenb_mprj[29]),
    .X(net309));
 sky130_fd_sc_hd__buf_4 input310 (.A(la_oenb_mprj[2]),
    .X(net310));
 sky130_fd_sc_hd__buf_6 input311 (.A(la_oenb_mprj[30]),
    .X(net311));
 sky130_fd_sc_hd__buf_8 input312 (.A(la_oenb_mprj[31]),
    .X(net312));
 sky130_fd_sc_hd__buf_6 input313 (.A(la_oenb_mprj[32]),
    .X(net313));
 sky130_fd_sc_hd__buf_4 input314 (.A(la_oenb_mprj[33]),
    .X(net314));
 sky130_fd_sc_hd__buf_4 input315 (.A(la_oenb_mprj[34]),
    .X(net315));
 sky130_fd_sc_hd__buf_6 input316 (.A(la_oenb_mprj[35]),
    .X(net316));
 sky130_fd_sc_hd__buf_8 input317 (.A(la_oenb_mprj[36]),
    .X(net317));
 sky130_fd_sc_hd__buf_8 input318 (.A(la_oenb_mprj[37]),
    .X(net318));
 sky130_fd_sc_hd__clkbuf_4 input319 (.A(la_oenb_mprj[38]),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_4 input320 (.A(la_oenb_mprj[39]),
    .X(net320));
 sky130_fd_sc_hd__clkbuf_4 input321 (.A(la_oenb_mprj[3]),
    .X(net321));
 sky130_fd_sc_hd__buf_8 input322 (.A(la_oenb_mprj[40]),
    .X(net322));
 sky130_fd_sc_hd__buf_4 input323 (.A(la_oenb_mprj[41]),
    .X(net323));
 sky130_fd_sc_hd__clkbuf_4 input324 (.A(la_oenb_mprj[42]),
    .X(net324));
 sky130_fd_sc_hd__buf_8 input325 (.A(la_oenb_mprj[43]),
    .X(net325));
 sky130_fd_sc_hd__buf_4 input326 (.A(la_oenb_mprj[44]),
    .X(net326));
 sky130_fd_sc_hd__buf_4 input327 (.A(la_oenb_mprj[45]),
    .X(net327));
 sky130_fd_sc_hd__buf_8 input328 (.A(la_oenb_mprj[46]),
    .X(net328));
 sky130_fd_sc_hd__buf_8 input329 (.A(la_oenb_mprj[47]),
    .X(net329));
 sky130_fd_sc_hd__buf_6 input330 (.A(la_oenb_mprj[48]),
    .X(net330));
 sky130_fd_sc_hd__buf_4 input331 (.A(la_oenb_mprj[49]),
    .X(net331));
 sky130_fd_sc_hd__clkbuf_4 input332 (.A(la_oenb_mprj[4]),
    .X(net332));
 sky130_fd_sc_hd__clkbuf_8 input333 (.A(la_oenb_mprj[50]),
    .X(net333));
 sky130_fd_sc_hd__buf_6 input334 (.A(la_oenb_mprj[51]),
    .X(net334));
 sky130_fd_sc_hd__buf_4 input335 (.A(la_oenb_mprj[52]),
    .X(net335));
 sky130_fd_sc_hd__buf_4 input336 (.A(la_oenb_mprj[53]),
    .X(net336));
 sky130_fd_sc_hd__buf_6 input337 (.A(la_oenb_mprj[54]),
    .X(net337));
 sky130_fd_sc_hd__clkbuf_4 input338 (.A(la_oenb_mprj[55]),
    .X(net338));
 sky130_fd_sc_hd__buf_4 input339 (.A(la_oenb_mprj[56]),
    .X(net339));
 sky130_fd_sc_hd__buf_4 input340 (.A(la_oenb_mprj[57]),
    .X(net340));
 sky130_fd_sc_hd__buf_6 input341 (.A(la_oenb_mprj[58]),
    .X(net341));
 sky130_fd_sc_hd__buf_4 input342 (.A(la_oenb_mprj[59]),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_4 input343 (.A(la_oenb_mprj[5]),
    .X(net343));
 sky130_fd_sc_hd__clkbuf_4 input344 (.A(la_oenb_mprj[60]),
    .X(net344));
 sky130_fd_sc_hd__clkbuf_4 input345 (.A(la_oenb_mprj[61]),
    .X(net345));
 sky130_fd_sc_hd__buf_6 input346 (.A(la_oenb_mprj[62]),
    .X(net346));
 sky130_fd_sc_hd__buf_6 input347 (.A(la_oenb_mprj[63]),
    .X(net347));
 sky130_fd_sc_hd__buf_6 input348 (.A(la_oenb_mprj[64]),
    .X(net348));
 sky130_fd_sc_hd__buf_6 input349 (.A(la_oenb_mprj[65]),
    .X(net349));
 sky130_fd_sc_hd__buf_6 input350 (.A(la_oenb_mprj[66]),
    .X(net350));
 sky130_fd_sc_hd__buf_6 input351 (.A(la_oenb_mprj[67]),
    .X(net351));
 sky130_fd_sc_hd__buf_8 input352 (.A(la_oenb_mprj[68]),
    .X(net352));
 sky130_fd_sc_hd__buf_8 input353 (.A(la_oenb_mprj[69]),
    .X(net353));
 sky130_fd_sc_hd__clkbuf_4 input354 (.A(la_oenb_mprj[6]),
    .X(net354));
 sky130_fd_sc_hd__buf_8 input355 (.A(la_oenb_mprj[70]),
    .X(net355));
 sky130_fd_sc_hd__buf_8 input356 (.A(la_oenb_mprj[71]),
    .X(net356));
 sky130_fd_sc_hd__buf_8 input357 (.A(la_oenb_mprj[72]),
    .X(net357));
 sky130_fd_sc_hd__buf_8 input358 (.A(la_oenb_mprj[73]),
    .X(net358));
 sky130_fd_sc_hd__buf_8 input359 (.A(la_oenb_mprj[74]),
    .X(net359));
 sky130_fd_sc_hd__buf_8 input360 (.A(la_oenb_mprj[75]),
    .X(net360));
 sky130_fd_sc_hd__buf_8 input361 (.A(la_oenb_mprj[76]),
    .X(net361));
 sky130_fd_sc_hd__buf_8 input362 (.A(la_oenb_mprj[77]),
    .X(net362));
 sky130_fd_sc_hd__buf_8 input363 (.A(la_oenb_mprj[78]),
    .X(net363));
 sky130_fd_sc_hd__buf_8 input364 (.A(la_oenb_mprj[79]),
    .X(net364));
 sky130_fd_sc_hd__clkbuf_4 input365 (.A(la_oenb_mprj[7]),
    .X(net365));
 sky130_fd_sc_hd__buf_8 input366 (.A(la_oenb_mprj[80]),
    .X(net366));
 sky130_fd_sc_hd__buf_8 input367 (.A(la_oenb_mprj[81]),
    .X(net367));
 sky130_fd_sc_hd__buf_8 input368 (.A(la_oenb_mprj[82]),
    .X(net368));
 sky130_fd_sc_hd__buf_8 input369 (.A(la_oenb_mprj[83]),
    .X(net369));
 sky130_fd_sc_hd__buf_8 input370 (.A(la_oenb_mprj[84]),
    .X(net370));
 sky130_fd_sc_hd__buf_8 input371 (.A(la_oenb_mprj[85]),
    .X(net371));
 sky130_fd_sc_hd__buf_8 input372 (.A(la_oenb_mprj[86]),
    .X(net372));
 sky130_fd_sc_hd__buf_8 input373 (.A(la_oenb_mprj[87]),
    .X(net373));
 sky130_fd_sc_hd__buf_8 input374 (.A(la_oenb_mprj[88]),
    .X(net374));
 sky130_fd_sc_hd__buf_4 input375 (.A(la_oenb_mprj[89]),
    .X(net375));
 sky130_fd_sc_hd__buf_4 input376 (.A(la_oenb_mprj[8]),
    .X(net376));
 sky130_fd_sc_hd__buf_4 input377 (.A(la_oenb_mprj[90]),
    .X(net377));
 sky130_fd_sc_hd__buf_6 input378 (.A(la_oenb_mprj[91]),
    .X(net378));
 sky130_fd_sc_hd__buf_6 input379 (.A(la_oenb_mprj[92]),
    .X(net379));
 sky130_fd_sc_hd__buf_8 input380 (.A(la_oenb_mprj[93]),
    .X(net380));
 sky130_fd_sc_hd__buf_8 input381 (.A(la_oenb_mprj[94]),
    .X(net381));
 sky130_fd_sc_hd__buf_8 input382 (.A(la_oenb_mprj[95]),
    .X(net382));
 sky130_fd_sc_hd__buf_6 input383 (.A(la_oenb_mprj[96]),
    .X(net383));
 sky130_fd_sc_hd__buf_6 input384 (.A(la_oenb_mprj[97]),
    .X(net384));
 sky130_fd_sc_hd__buf_6 input385 (.A(la_oenb_mprj[98]),
    .X(net385));
 sky130_fd_sc_hd__buf_6 input386 (.A(la_oenb_mprj[99]),
    .X(net386));
 sky130_fd_sc_hd__clkbuf_4 input387 (.A(la_oenb_mprj[9]),
    .X(net387));
 sky130_fd_sc_hd__buf_8 input388 (.A(mprj_adr_o_core[0]),
    .X(net388));
 sky130_fd_sc_hd__buf_8 input389 (.A(mprj_adr_o_core[10]),
    .X(net389));
 sky130_fd_sc_hd__buf_8 input390 (.A(mprj_adr_o_core[11]),
    .X(net390));
 sky130_fd_sc_hd__buf_8 input391 (.A(mprj_adr_o_core[12]),
    .X(net391));
 sky130_fd_sc_hd__buf_8 input392 (.A(mprj_adr_o_core[13]),
    .X(net392));
 sky130_fd_sc_hd__buf_8 input393 (.A(mprj_adr_o_core[14]),
    .X(net393));
 sky130_fd_sc_hd__buf_8 input394 (.A(mprj_adr_o_core[15]),
    .X(net394));
 sky130_fd_sc_hd__buf_8 input395 (.A(mprj_adr_o_core[16]),
    .X(net395));
 sky130_fd_sc_hd__buf_8 input396 (.A(mprj_adr_o_core[17]),
    .X(net396));
 sky130_fd_sc_hd__buf_8 input397 (.A(mprj_adr_o_core[18]),
    .X(net397));
 sky130_fd_sc_hd__buf_8 input398 (.A(mprj_adr_o_core[19]),
    .X(net398));
 sky130_fd_sc_hd__buf_8 input399 (.A(mprj_adr_o_core[1]),
    .X(net399));
 sky130_fd_sc_hd__buf_8 input400 (.A(mprj_adr_o_core[20]),
    .X(net400));
 sky130_fd_sc_hd__buf_8 input401 (.A(mprj_adr_o_core[21]),
    .X(net401));
 sky130_fd_sc_hd__buf_8 input402 (.A(mprj_adr_o_core[22]),
    .X(net402));
 sky130_fd_sc_hd__buf_8 input403 (.A(mprj_adr_o_core[23]),
    .X(net403));
 sky130_fd_sc_hd__buf_8 input404 (.A(mprj_adr_o_core[24]),
    .X(net404));
 sky130_fd_sc_hd__buf_8 input405 (.A(mprj_adr_o_core[25]),
    .X(net405));
 sky130_fd_sc_hd__buf_8 input406 (.A(mprj_adr_o_core[26]),
    .X(net406));
 sky130_fd_sc_hd__buf_8 input407 (.A(mprj_adr_o_core[27]),
    .X(net407));
 sky130_fd_sc_hd__buf_8 input408 (.A(mprj_adr_o_core[28]),
    .X(net408));
 sky130_fd_sc_hd__buf_8 input409 (.A(mprj_adr_o_core[29]),
    .X(net409));
 sky130_fd_sc_hd__buf_8 input410 (.A(mprj_adr_o_core[2]),
    .X(net410));
 sky130_fd_sc_hd__buf_8 input411 (.A(mprj_adr_o_core[30]),
    .X(net411));
 sky130_fd_sc_hd__buf_8 input412 (.A(mprj_adr_o_core[31]),
    .X(net412));
 sky130_fd_sc_hd__buf_8 input413 (.A(mprj_adr_o_core[3]),
    .X(net413));
 sky130_fd_sc_hd__buf_8 input414 (.A(mprj_adr_o_core[4]),
    .X(net414));
 sky130_fd_sc_hd__buf_8 input415 (.A(mprj_adr_o_core[5]),
    .X(net415));
 sky130_fd_sc_hd__buf_8 input416 (.A(mprj_adr_o_core[6]),
    .X(net416));
 sky130_fd_sc_hd__buf_8 input417 (.A(mprj_adr_o_core[7]),
    .X(net417));
 sky130_fd_sc_hd__buf_8 input418 (.A(mprj_adr_o_core[8]),
    .X(net418));
 sky130_fd_sc_hd__buf_8 input419 (.A(mprj_adr_o_core[9]),
    .X(net419));
 sky130_fd_sc_hd__buf_8 input420 (.A(mprj_cyc_o_core),
    .X(net420));
 sky130_fd_sc_hd__buf_8 input421 (.A(mprj_dat_o_core[0]),
    .X(net421));
 sky130_fd_sc_hd__buf_8 input422 (.A(mprj_dat_o_core[10]),
    .X(net422));
 sky130_fd_sc_hd__buf_8 input423 (.A(mprj_dat_o_core[11]),
    .X(net423));
 sky130_fd_sc_hd__buf_8 input424 (.A(mprj_dat_o_core[12]),
    .X(net424));
 sky130_fd_sc_hd__buf_8 input425 (.A(mprj_dat_o_core[13]),
    .X(net425));
 sky130_fd_sc_hd__buf_8 input426 (.A(mprj_dat_o_core[14]),
    .X(net426));
 sky130_fd_sc_hd__buf_8 input427 (.A(mprj_dat_o_core[15]),
    .X(net427));
 sky130_fd_sc_hd__buf_8 input428 (.A(mprj_dat_o_core[16]),
    .X(net428));
 sky130_fd_sc_hd__buf_8 input429 (.A(mprj_dat_o_core[17]),
    .X(net429));
 sky130_fd_sc_hd__buf_8 input430 (.A(mprj_dat_o_core[18]),
    .X(net430));
 sky130_fd_sc_hd__buf_8 input431 (.A(mprj_dat_o_core[19]),
    .X(net431));
 sky130_fd_sc_hd__buf_8 input432 (.A(mprj_dat_o_core[1]),
    .X(net432));
 sky130_fd_sc_hd__buf_8 input433 (.A(mprj_dat_o_core[20]),
    .X(net433));
 sky130_fd_sc_hd__buf_8 input434 (.A(mprj_dat_o_core[21]),
    .X(net434));
 sky130_fd_sc_hd__buf_8 input435 (.A(mprj_dat_o_core[22]),
    .X(net435));
 sky130_fd_sc_hd__buf_8 input436 (.A(mprj_dat_o_core[23]),
    .X(net436));
 sky130_fd_sc_hd__buf_8 input437 (.A(mprj_dat_o_core[24]),
    .X(net437));
 sky130_fd_sc_hd__buf_8 input438 (.A(mprj_dat_o_core[25]),
    .X(net438));
 sky130_fd_sc_hd__buf_8 input439 (.A(mprj_dat_o_core[26]),
    .X(net439));
 sky130_fd_sc_hd__buf_8 input440 (.A(mprj_dat_o_core[27]),
    .X(net440));
 sky130_fd_sc_hd__buf_6 input441 (.A(mprj_dat_o_core[28]),
    .X(net441));
 sky130_fd_sc_hd__buf_6 input442 (.A(mprj_dat_o_core[29]),
    .X(net442));
 sky130_fd_sc_hd__buf_8 input443 (.A(mprj_dat_o_core[2]),
    .X(net443));
 sky130_fd_sc_hd__buf_6 input444 (.A(mprj_dat_o_core[30]),
    .X(net444));
 sky130_fd_sc_hd__buf_6 input445 (.A(mprj_dat_o_core[31]),
    .X(net445));
 sky130_fd_sc_hd__buf_8 input446 (.A(mprj_dat_o_core[3]),
    .X(net446));
 sky130_fd_sc_hd__buf_8 input447 (.A(mprj_dat_o_core[4]),
    .X(net447));
 sky130_fd_sc_hd__buf_8 input448 (.A(mprj_dat_o_core[5]),
    .X(net448));
 sky130_fd_sc_hd__buf_8 input449 (.A(mprj_dat_o_core[6]),
    .X(net449));
 sky130_fd_sc_hd__buf_8 input450 (.A(mprj_dat_o_core[7]),
    .X(net450));
 sky130_fd_sc_hd__buf_8 input451 (.A(mprj_dat_o_core[8]),
    .X(net451));
 sky130_fd_sc_hd__buf_8 input452 (.A(mprj_dat_o_core[9]),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_4 input453 (.A(mprj_iena_wb),
    .X(net453));
 sky130_fd_sc_hd__buf_8 input454 (.A(mprj_sel_o_core[0]),
    .X(net454));
 sky130_fd_sc_hd__buf_8 input455 (.A(mprj_sel_o_core[1]),
    .X(net455));
 sky130_fd_sc_hd__buf_8 input456 (.A(mprj_sel_o_core[2]),
    .X(net456));
 sky130_fd_sc_hd__buf_8 input457 (.A(mprj_sel_o_core[3]),
    .X(net457));
 sky130_fd_sc_hd__buf_8 input458 (.A(mprj_stb_o_core),
    .X(net458));
 sky130_fd_sc_hd__buf_8 input459 (.A(mprj_we_o_core),
    .X(net459));
 sky130_fd_sc_hd__clkbuf_4 input460 (.A(user_irq_ena[0]),
    .X(net460));
 sky130_fd_sc_hd__clkbuf_4 input461 (.A(user_irq_ena[1]),
    .X(net461));
 sky130_fd_sc_hd__clkbuf_4 input462 (.A(user_irq_ena[2]),
    .X(net462));
 sky130_fd_sc_hd__buf_8 output463 (.A(net463),
    .X(la_data_in_core[0]));
 sky130_fd_sc_hd__buf_8 output464 (.A(net464),
    .X(la_data_in_core[100]));
 sky130_fd_sc_hd__buf_8 output465 (.A(net465),
    .X(la_data_in_core[101]));
 sky130_fd_sc_hd__buf_8 output466 (.A(net466),
    .X(la_data_in_core[102]));
 sky130_fd_sc_hd__buf_8 output467 (.A(net467),
    .X(la_data_in_core[103]));
 sky130_fd_sc_hd__buf_8 output468 (.A(net468),
    .X(la_data_in_core[104]));
 sky130_fd_sc_hd__buf_8 output469 (.A(net469),
    .X(la_data_in_core[105]));
 sky130_fd_sc_hd__buf_8 output470 (.A(net470),
    .X(la_data_in_core[106]));
 sky130_fd_sc_hd__buf_8 output471 (.A(net471),
    .X(la_data_in_core[107]));
 sky130_fd_sc_hd__buf_8 output472 (.A(net472),
    .X(la_data_in_core[108]));
 sky130_fd_sc_hd__buf_8 output473 (.A(net473),
    .X(la_data_in_core[109]));
 sky130_fd_sc_hd__buf_8 output474 (.A(net474),
    .X(la_data_in_core[10]));
 sky130_fd_sc_hd__buf_8 output475 (.A(net475),
    .X(la_data_in_core[110]));
 sky130_fd_sc_hd__buf_8 output476 (.A(net476),
    .X(la_data_in_core[111]));
 sky130_fd_sc_hd__buf_8 output477 (.A(net477),
    .X(la_data_in_core[112]));
 sky130_fd_sc_hd__buf_8 output478 (.A(net478),
    .X(la_data_in_core[113]));
 sky130_fd_sc_hd__buf_8 output479 (.A(net479),
    .X(la_data_in_core[114]));
 sky130_fd_sc_hd__buf_8 output480 (.A(net480),
    .X(la_data_in_core[115]));
 sky130_fd_sc_hd__buf_8 output481 (.A(net481),
    .X(la_data_in_core[116]));
 sky130_fd_sc_hd__buf_8 output482 (.A(net482),
    .X(la_data_in_core[117]));
 sky130_fd_sc_hd__buf_8 output483 (.A(net483),
    .X(la_data_in_core[118]));
 sky130_fd_sc_hd__buf_8 output484 (.A(net484),
    .X(la_data_in_core[119]));
 sky130_fd_sc_hd__buf_8 output485 (.A(net485),
    .X(la_data_in_core[11]));
 sky130_fd_sc_hd__buf_8 output486 (.A(net486),
    .X(la_data_in_core[120]));
 sky130_fd_sc_hd__buf_8 output487 (.A(net487),
    .X(la_data_in_core[121]));
 sky130_fd_sc_hd__buf_8 output488 (.A(net488),
    .X(la_data_in_core[122]));
 sky130_fd_sc_hd__buf_8 output489 (.A(net489),
    .X(la_data_in_core[123]));
 sky130_fd_sc_hd__buf_8 output490 (.A(net490),
    .X(la_data_in_core[124]));
 sky130_fd_sc_hd__buf_8 output491 (.A(net491),
    .X(la_data_in_core[125]));
 sky130_fd_sc_hd__buf_8 output492 (.A(net492),
    .X(la_data_in_core[126]));
 sky130_fd_sc_hd__buf_8 output493 (.A(net493),
    .X(la_data_in_core[127]));
 sky130_fd_sc_hd__buf_8 output494 (.A(net494),
    .X(la_data_in_core[12]));
 sky130_fd_sc_hd__buf_8 output495 (.A(net495),
    .X(la_data_in_core[13]));
 sky130_fd_sc_hd__buf_8 output496 (.A(net496),
    .X(la_data_in_core[14]));
 sky130_fd_sc_hd__buf_8 output497 (.A(net497),
    .X(la_data_in_core[15]));
 sky130_fd_sc_hd__buf_8 output498 (.A(net498),
    .X(la_data_in_core[16]));
 sky130_fd_sc_hd__buf_8 output499 (.A(net499),
    .X(la_data_in_core[17]));
 sky130_fd_sc_hd__buf_8 output500 (.A(net500),
    .X(la_data_in_core[18]));
 sky130_fd_sc_hd__buf_8 output501 (.A(net501),
    .X(la_data_in_core[19]));
 sky130_fd_sc_hd__buf_8 output502 (.A(net502),
    .X(la_data_in_core[1]));
 sky130_fd_sc_hd__buf_8 output503 (.A(net503),
    .X(la_data_in_core[20]));
 sky130_fd_sc_hd__buf_8 output504 (.A(net504),
    .X(la_data_in_core[21]));
 sky130_fd_sc_hd__buf_8 output505 (.A(net505),
    .X(la_data_in_core[22]));
 sky130_fd_sc_hd__buf_8 output506 (.A(net506),
    .X(la_data_in_core[23]));
 sky130_fd_sc_hd__buf_8 output507 (.A(net507),
    .X(la_data_in_core[24]));
 sky130_fd_sc_hd__buf_8 output508 (.A(net508),
    .X(la_data_in_core[25]));
 sky130_fd_sc_hd__buf_8 output509 (.A(net509),
    .X(la_data_in_core[26]));
 sky130_fd_sc_hd__buf_8 output510 (.A(net510),
    .X(la_data_in_core[27]));
 sky130_fd_sc_hd__buf_8 output511 (.A(net511),
    .X(la_data_in_core[28]));
 sky130_fd_sc_hd__buf_8 output512 (.A(net512),
    .X(la_data_in_core[29]));
 sky130_fd_sc_hd__buf_8 output513 (.A(net513),
    .X(la_data_in_core[2]));
 sky130_fd_sc_hd__buf_8 output514 (.A(net514),
    .X(la_data_in_core[30]));
 sky130_fd_sc_hd__buf_8 output515 (.A(net515),
    .X(la_data_in_core[31]));
 sky130_fd_sc_hd__buf_8 output516 (.A(net516),
    .X(la_data_in_core[32]));
 sky130_fd_sc_hd__buf_8 output517 (.A(net517),
    .X(la_data_in_core[33]));
 sky130_fd_sc_hd__buf_8 output518 (.A(net518),
    .X(la_data_in_core[34]));
 sky130_fd_sc_hd__buf_8 output519 (.A(net519),
    .X(la_data_in_core[35]));
 sky130_fd_sc_hd__buf_8 output520 (.A(net520),
    .X(la_data_in_core[36]));
 sky130_fd_sc_hd__buf_8 output521 (.A(net521),
    .X(la_data_in_core[37]));
 sky130_fd_sc_hd__buf_8 output522 (.A(net522),
    .X(la_data_in_core[38]));
 sky130_fd_sc_hd__buf_8 output523 (.A(net523),
    .X(la_data_in_core[39]));
 sky130_fd_sc_hd__buf_8 output524 (.A(net524),
    .X(la_data_in_core[3]));
 sky130_fd_sc_hd__buf_8 output525 (.A(net525),
    .X(la_data_in_core[40]));
 sky130_fd_sc_hd__buf_8 output526 (.A(net526),
    .X(la_data_in_core[41]));
 sky130_fd_sc_hd__buf_8 output527 (.A(net527),
    .X(la_data_in_core[42]));
 sky130_fd_sc_hd__buf_8 output528 (.A(net528),
    .X(la_data_in_core[43]));
 sky130_fd_sc_hd__buf_8 output529 (.A(net529),
    .X(la_data_in_core[44]));
 sky130_fd_sc_hd__buf_8 output530 (.A(net530),
    .X(la_data_in_core[45]));
 sky130_fd_sc_hd__buf_8 output531 (.A(net531),
    .X(la_data_in_core[46]));
 sky130_fd_sc_hd__buf_8 output532 (.A(net532),
    .X(la_data_in_core[47]));
 sky130_fd_sc_hd__buf_8 output533 (.A(net533),
    .X(la_data_in_core[48]));
 sky130_fd_sc_hd__buf_8 output534 (.A(net534),
    .X(la_data_in_core[49]));
 sky130_fd_sc_hd__buf_8 output535 (.A(net535),
    .X(la_data_in_core[4]));
 sky130_fd_sc_hd__buf_8 output536 (.A(net536),
    .X(la_data_in_core[50]));
 sky130_fd_sc_hd__buf_8 output537 (.A(net537),
    .X(la_data_in_core[51]));
 sky130_fd_sc_hd__buf_8 output538 (.A(net538),
    .X(la_data_in_core[52]));
 sky130_fd_sc_hd__buf_8 output539 (.A(net539),
    .X(la_data_in_core[53]));
 sky130_fd_sc_hd__buf_8 output540 (.A(net540),
    .X(la_data_in_core[54]));
 sky130_fd_sc_hd__buf_8 output541 (.A(net541),
    .X(la_data_in_core[55]));
 sky130_fd_sc_hd__buf_8 output542 (.A(net542),
    .X(la_data_in_core[56]));
 sky130_fd_sc_hd__buf_8 output543 (.A(net543),
    .X(la_data_in_core[57]));
 sky130_fd_sc_hd__buf_8 output544 (.A(net544),
    .X(la_data_in_core[58]));
 sky130_fd_sc_hd__buf_8 output545 (.A(net545),
    .X(la_data_in_core[59]));
 sky130_fd_sc_hd__buf_8 output546 (.A(net546),
    .X(la_data_in_core[5]));
 sky130_fd_sc_hd__buf_8 output547 (.A(net547),
    .X(la_data_in_core[60]));
 sky130_fd_sc_hd__buf_8 output548 (.A(net548),
    .X(la_data_in_core[61]));
 sky130_fd_sc_hd__buf_8 output549 (.A(net549),
    .X(la_data_in_core[62]));
 sky130_fd_sc_hd__buf_8 output550 (.A(net550),
    .X(la_data_in_core[63]));
 sky130_fd_sc_hd__buf_8 output551 (.A(net551),
    .X(la_data_in_core[64]));
 sky130_fd_sc_hd__buf_8 output552 (.A(net552),
    .X(la_data_in_core[65]));
 sky130_fd_sc_hd__buf_8 output553 (.A(net553),
    .X(la_data_in_core[66]));
 sky130_fd_sc_hd__buf_8 output554 (.A(net554),
    .X(la_data_in_core[67]));
 sky130_fd_sc_hd__buf_8 output555 (.A(net555),
    .X(la_data_in_core[68]));
 sky130_fd_sc_hd__buf_8 output556 (.A(net556),
    .X(la_data_in_core[69]));
 sky130_fd_sc_hd__buf_8 output557 (.A(net557),
    .X(la_data_in_core[6]));
 sky130_fd_sc_hd__buf_8 output558 (.A(net558),
    .X(la_data_in_core[70]));
 sky130_fd_sc_hd__buf_8 output559 (.A(net559),
    .X(la_data_in_core[71]));
 sky130_fd_sc_hd__buf_8 output560 (.A(net560),
    .X(la_data_in_core[72]));
 sky130_fd_sc_hd__buf_8 output561 (.A(net561),
    .X(la_data_in_core[73]));
 sky130_fd_sc_hd__buf_8 output562 (.A(net562),
    .X(la_data_in_core[74]));
 sky130_fd_sc_hd__buf_8 output563 (.A(net563),
    .X(la_data_in_core[75]));
 sky130_fd_sc_hd__buf_8 output564 (.A(net564),
    .X(la_data_in_core[76]));
 sky130_fd_sc_hd__buf_8 output565 (.A(net565),
    .X(la_data_in_core[77]));
 sky130_fd_sc_hd__buf_8 output566 (.A(net566),
    .X(la_data_in_core[78]));
 sky130_fd_sc_hd__buf_8 output567 (.A(net567),
    .X(la_data_in_core[79]));
 sky130_fd_sc_hd__buf_8 output568 (.A(net568),
    .X(la_data_in_core[7]));
 sky130_fd_sc_hd__buf_8 output569 (.A(net569),
    .X(la_data_in_core[80]));
 sky130_fd_sc_hd__buf_8 output570 (.A(net570),
    .X(la_data_in_core[81]));
 sky130_fd_sc_hd__buf_8 output571 (.A(net571),
    .X(la_data_in_core[82]));
 sky130_fd_sc_hd__buf_8 output572 (.A(net572),
    .X(la_data_in_core[83]));
 sky130_fd_sc_hd__buf_8 output573 (.A(net573),
    .X(la_data_in_core[84]));
 sky130_fd_sc_hd__buf_8 output574 (.A(net574),
    .X(la_data_in_core[85]));
 sky130_fd_sc_hd__buf_8 output575 (.A(net575),
    .X(la_data_in_core[86]));
 sky130_fd_sc_hd__buf_8 output576 (.A(net576),
    .X(la_data_in_core[87]));
 sky130_fd_sc_hd__buf_8 output577 (.A(net577),
    .X(la_data_in_core[88]));
 sky130_fd_sc_hd__buf_8 output578 (.A(net578),
    .X(la_data_in_core[89]));
 sky130_fd_sc_hd__buf_8 output579 (.A(net579),
    .X(la_data_in_core[8]));
 sky130_fd_sc_hd__buf_8 output580 (.A(net580),
    .X(la_data_in_core[90]));
 sky130_fd_sc_hd__buf_8 output581 (.A(net581),
    .X(la_data_in_core[91]));
 sky130_fd_sc_hd__buf_8 output582 (.A(net582),
    .X(la_data_in_core[92]));
 sky130_fd_sc_hd__buf_8 output583 (.A(net583),
    .X(la_data_in_core[93]));
 sky130_fd_sc_hd__buf_8 output584 (.A(net584),
    .X(la_data_in_core[94]));
 sky130_fd_sc_hd__buf_8 output585 (.A(net585),
    .X(la_data_in_core[95]));
 sky130_fd_sc_hd__buf_8 output586 (.A(net586),
    .X(la_data_in_core[96]));
 sky130_fd_sc_hd__buf_8 output587 (.A(net587),
    .X(la_data_in_core[97]));
 sky130_fd_sc_hd__buf_8 output588 (.A(net588),
    .X(la_data_in_core[98]));
 sky130_fd_sc_hd__buf_8 output589 (.A(net589),
    .X(la_data_in_core[99]));
 sky130_fd_sc_hd__buf_8 output590 (.A(net590),
    .X(la_data_in_core[9]));
 sky130_fd_sc_hd__buf_8 output591 (.A(net591),
    .X(la_data_in_mprj[0]));
 sky130_fd_sc_hd__buf_8 output592 (.A(net592),
    .X(la_data_in_mprj[100]));
 sky130_fd_sc_hd__buf_8 output593 (.A(net593),
    .X(la_data_in_mprj[101]));
 sky130_fd_sc_hd__buf_8 output594 (.A(net594),
    .X(la_data_in_mprj[102]));
 sky130_fd_sc_hd__buf_8 output595 (.A(net595),
    .X(la_data_in_mprj[103]));
 sky130_fd_sc_hd__buf_8 output596 (.A(net596),
    .X(la_data_in_mprj[104]));
 sky130_fd_sc_hd__buf_8 output597 (.A(net597),
    .X(la_data_in_mprj[105]));
 sky130_fd_sc_hd__buf_8 output598 (.A(net598),
    .X(la_data_in_mprj[106]));
 sky130_fd_sc_hd__buf_8 output599 (.A(net599),
    .X(la_data_in_mprj[107]));
 sky130_fd_sc_hd__buf_8 output600 (.A(net600),
    .X(la_data_in_mprj[108]));
 sky130_fd_sc_hd__buf_8 output601 (.A(net601),
    .X(la_data_in_mprj[109]));
 sky130_fd_sc_hd__buf_8 output602 (.A(net602),
    .X(la_data_in_mprj[10]));
 sky130_fd_sc_hd__buf_8 output603 (.A(net603),
    .X(la_data_in_mprj[110]));
 sky130_fd_sc_hd__buf_8 output604 (.A(net604),
    .X(la_data_in_mprj[111]));
 sky130_fd_sc_hd__buf_8 output605 (.A(net605),
    .X(la_data_in_mprj[112]));
 sky130_fd_sc_hd__buf_8 output606 (.A(net606),
    .X(la_data_in_mprj[113]));
 sky130_fd_sc_hd__buf_8 output607 (.A(net607),
    .X(la_data_in_mprj[114]));
 sky130_fd_sc_hd__buf_8 output608 (.A(net608),
    .X(la_data_in_mprj[115]));
 sky130_fd_sc_hd__buf_8 output609 (.A(net609),
    .X(la_data_in_mprj[116]));
 sky130_fd_sc_hd__buf_8 output610 (.A(net610),
    .X(la_data_in_mprj[117]));
 sky130_fd_sc_hd__buf_8 output611 (.A(net611),
    .X(la_data_in_mprj[118]));
 sky130_fd_sc_hd__buf_8 output612 (.A(net612),
    .X(la_data_in_mprj[119]));
 sky130_fd_sc_hd__buf_8 output613 (.A(net613),
    .X(la_data_in_mprj[11]));
 sky130_fd_sc_hd__buf_8 output614 (.A(net614),
    .X(la_data_in_mprj[120]));
 sky130_fd_sc_hd__buf_8 output615 (.A(net615),
    .X(la_data_in_mprj[121]));
 sky130_fd_sc_hd__buf_8 output616 (.A(net616),
    .X(la_data_in_mprj[122]));
 sky130_fd_sc_hd__buf_8 output617 (.A(net617),
    .X(la_data_in_mprj[123]));
 sky130_fd_sc_hd__buf_8 output618 (.A(net618),
    .X(la_data_in_mprj[124]));
 sky130_fd_sc_hd__buf_8 output619 (.A(net619),
    .X(la_data_in_mprj[125]));
 sky130_fd_sc_hd__buf_8 output620 (.A(net620),
    .X(la_data_in_mprj[126]));
 sky130_fd_sc_hd__buf_8 output621 (.A(net621),
    .X(la_data_in_mprj[127]));
 sky130_fd_sc_hd__buf_8 output622 (.A(net622),
    .X(la_data_in_mprj[12]));
 sky130_fd_sc_hd__buf_8 output623 (.A(net623),
    .X(la_data_in_mprj[13]));
 sky130_fd_sc_hd__buf_8 output624 (.A(net624),
    .X(la_data_in_mprj[14]));
 sky130_fd_sc_hd__buf_8 output625 (.A(net625),
    .X(la_data_in_mprj[15]));
 sky130_fd_sc_hd__buf_8 output626 (.A(net626),
    .X(la_data_in_mprj[16]));
 sky130_fd_sc_hd__buf_8 output627 (.A(net627),
    .X(la_data_in_mprj[17]));
 sky130_fd_sc_hd__buf_8 output628 (.A(net628),
    .X(la_data_in_mprj[18]));
 sky130_fd_sc_hd__buf_8 output629 (.A(net629),
    .X(la_data_in_mprj[19]));
 sky130_fd_sc_hd__buf_8 output630 (.A(net630),
    .X(la_data_in_mprj[1]));
 sky130_fd_sc_hd__buf_8 output631 (.A(net631),
    .X(la_data_in_mprj[20]));
 sky130_fd_sc_hd__buf_8 output632 (.A(net632),
    .X(la_data_in_mprj[21]));
 sky130_fd_sc_hd__buf_8 output633 (.A(net633),
    .X(la_data_in_mprj[22]));
 sky130_fd_sc_hd__buf_8 output634 (.A(net634),
    .X(la_data_in_mprj[23]));
 sky130_fd_sc_hd__buf_8 output635 (.A(net635),
    .X(la_data_in_mprj[24]));
 sky130_fd_sc_hd__buf_8 output636 (.A(net636),
    .X(la_data_in_mprj[25]));
 sky130_fd_sc_hd__buf_8 output637 (.A(net637),
    .X(la_data_in_mprj[26]));
 sky130_fd_sc_hd__buf_8 output638 (.A(net638),
    .X(la_data_in_mprj[27]));
 sky130_fd_sc_hd__buf_8 output639 (.A(net639),
    .X(la_data_in_mprj[28]));
 sky130_fd_sc_hd__buf_8 output640 (.A(net640),
    .X(la_data_in_mprj[29]));
 sky130_fd_sc_hd__buf_8 output641 (.A(net641),
    .X(la_data_in_mprj[2]));
 sky130_fd_sc_hd__buf_8 output642 (.A(net642),
    .X(la_data_in_mprj[30]));
 sky130_fd_sc_hd__buf_8 output643 (.A(net643),
    .X(la_data_in_mprj[31]));
 sky130_fd_sc_hd__buf_8 output644 (.A(net644),
    .X(la_data_in_mprj[32]));
 sky130_fd_sc_hd__buf_8 output645 (.A(net645),
    .X(la_data_in_mprj[33]));
 sky130_fd_sc_hd__buf_8 output646 (.A(net646),
    .X(la_data_in_mprj[34]));
 sky130_fd_sc_hd__buf_8 output647 (.A(net647),
    .X(la_data_in_mprj[35]));
 sky130_fd_sc_hd__buf_8 output648 (.A(net648),
    .X(la_data_in_mprj[36]));
 sky130_fd_sc_hd__buf_8 output649 (.A(net649),
    .X(la_data_in_mprj[37]));
 sky130_fd_sc_hd__buf_8 output650 (.A(net650),
    .X(la_data_in_mprj[38]));
 sky130_fd_sc_hd__buf_8 output651 (.A(net651),
    .X(la_data_in_mprj[39]));
 sky130_fd_sc_hd__buf_8 output652 (.A(net652),
    .X(la_data_in_mprj[3]));
 sky130_fd_sc_hd__buf_8 output653 (.A(net653),
    .X(la_data_in_mprj[40]));
 sky130_fd_sc_hd__buf_8 output654 (.A(net654),
    .X(la_data_in_mprj[41]));
 sky130_fd_sc_hd__buf_8 output655 (.A(net655),
    .X(la_data_in_mprj[42]));
 sky130_fd_sc_hd__buf_8 output656 (.A(net656),
    .X(la_data_in_mprj[43]));
 sky130_fd_sc_hd__buf_8 output657 (.A(net657),
    .X(la_data_in_mprj[44]));
 sky130_fd_sc_hd__buf_8 output658 (.A(net658),
    .X(la_data_in_mprj[45]));
 sky130_fd_sc_hd__buf_8 output659 (.A(net659),
    .X(la_data_in_mprj[46]));
 sky130_fd_sc_hd__buf_8 output660 (.A(net660),
    .X(la_data_in_mprj[47]));
 sky130_fd_sc_hd__buf_8 output661 (.A(net661),
    .X(la_data_in_mprj[48]));
 sky130_fd_sc_hd__buf_8 output662 (.A(net662),
    .X(la_data_in_mprj[49]));
 sky130_fd_sc_hd__buf_8 output663 (.A(net663),
    .X(la_data_in_mprj[4]));
 sky130_fd_sc_hd__buf_8 output664 (.A(net664),
    .X(la_data_in_mprj[50]));
 sky130_fd_sc_hd__buf_8 output665 (.A(net665),
    .X(la_data_in_mprj[51]));
 sky130_fd_sc_hd__buf_8 output666 (.A(net666),
    .X(la_data_in_mprj[52]));
 sky130_fd_sc_hd__buf_8 output667 (.A(net667),
    .X(la_data_in_mprj[53]));
 sky130_fd_sc_hd__buf_8 output668 (.A(net668),
    .X(la_data_in_mprj[54]));
 sky130_fd_sc_hd__buf_8 output669 (.A(net669),
    .X(la_data_in_mprj[55]));
 sky130_fd_sc_hd__buf_8 output670 (.A(net670),
    .X(la_data_in_mprj[56]));
 sky130_fd_sc_hd__buf_8 output671 (.A(net671),
    .X(la_data_in_mprj[57]));
 sky130_fd_sc_hd__buf_8 output672 (.A(net672),
    .X(la_data_in_mprj[58]));
 sky130_fd_sc_hd__buf_8 output673 (.A(net673),
    .X(la_data_in_mprj[59]));
 sky130_fd_sc_hd__buf_8 output674 (.A(net674),
    .X(la_data_in_mprj[5]));
 sky130_fd_sc_hd__buf_8 output675 (.A(net675),
    .X(la_data_in_mprj[60]));
 sky130_fd_sc_hd__buf_8 output676 (.A(net676),
    .X(la_data_in_mprj[61]));
 sky130_fd_sc_hd__buf_8 output677 (.A(net677),
    .X(la_data_in_mprj[62]));
 sky130_fd_sc_hd__buf_8 output678 (.A(net678),
    .X(la_data_in_mprj[63]));
 sky130_fd_sc_hd__buf_8 output679 (.A(net679),
    .X(la_data_in_mprj[64]));
 sky130_fd_sc_hd__buf_8 output680 (.A(net680),
    .X(la_data_in_mprj[65]));
 sky130_fd_sc_hd__buf_8 output681 (.A(net681),
    .X(la_data_in_mprj[66]));
 sky130_fd_sc_hd__buf_8 output682 (.A(net682),
    .X(la_data_in_mprj[67]));
 sky130_fd_sc_hd__buf_8 output683 (.A(net683),
    .X(la_data_in_mprj[68]));
 sky130_fd_sc_hd__buf_8 output684 (.A(net684),
    .X(la_data_in_mprj[69]));
 sky130_fd_sc_hd__buf_8 output685 (.A(net685),
    .X(la_data_in_mprj[6]));
 sky130_fd_sc_hd__buf_8 output686 (.A(net686),
    .X(la_data_in_mprj[70]));
 sky130_fd_sc_hd__buf_8 output687 (.A(net687),
    .X(la_data_in_mprj[71]));
 sky130_fd_sc_hd__buf_8 output688 (.A(net688),
    .X(la_data_in_mprj[72]));
 sky130_fd_sc_hd__buf_8 output689 (.A(net689),
    .X(la_data_in_mprj[73]));
 sky130_fd_sc_hd__buf_8 output690 (.A(net690),
    .X(la_data_in_mprj[74]));
 sky130_fd_sc_hd__buf_8 output691 (.A(net691),
    .X(la_data_in_mprj[75]));
 sky130_fd_sc_hd__buf_8 output692 (.A(net692),
    .X(la_data_in_mprj[76]));
 sky130_fd_sc_hd__buf_8 output693 (.A(net693),
    .X(la_data_in_mprj[77]));
 sky130_fd_sc_hd__buf_8 output694 (.A(net694),
    .X(la_data_in_mprj[78]));
 sky130_fd_sc_hd__buf_8 output695 (.A(net695),
    .X(la_data_in_mprj[79]));
 sky130_fd_sc_hd__buf_8 output696 (.A(net696),
    .X(la_data_in_mprj[7]));
 sky130_fd_sc_hd__buf_8 output697 (.A(net697),
    .X(la_data_in_mprj[80]));
 sky130_fd_sc_hd__buf_8 output698 (.A(net698),
    .X(la_data_in_mprj[81]));
 sky130_fd_sc_hd__buf_8 output699 (.A(net699),
    .X(la_data_in_mprj[82]));
 sky130_fd_sc_hd__buf_8 output700 (.A(net700),
    .X(la_data_in_mprj[83]));
 sky130_fd_sc_hd__buf_8 output701 (.A(net701),
    .X(la_data_in_mprj[84]));
 sky130_fd_sc_hd__buf_8 output702 (.A(net702),
    .X(la_data_in_mprj[85]));
 sky130_fd_sc_hd__buf_8 output703 (.A(net703),
    .X(la_data_in_mprj[86]));
 sky130_fd_sc_hd__buf_8 output704 (.A(net704),
    .X(la_data_in_mprj[87]));
 sky130_fd_sc_hd__buf_8 output705 (.A(net705),
    .X(la_data_in_mprj[88]));
 sky130_fd_sc_hd__buf_8 output706 (.A(net706),
    .X(la_data_in_mprj[89]));
 sky130_fd_sc_hd__buf_8 output707 (.A(net707),
    .X(la_data_in_mprj[8]));
 sky130_fd_sc_hd__buf_8 output708 (.A(net708),
    .X(la_data_in_mprj[90]));
 sky130_fd_sc_hd__buf_8 output709 (.A(net709),
    .X(la_data_in_mprj[91]));
 sky130_fd_sc_hd__buf_8 output710 (.A(net710),
    .X(la_data_in_mprj[92]));
 sky130_fd_sc_hd__buf_8 output711 (.A(net711),
    .X(la_data_in_mprj[93]));
 sky130_fd_sc_hd__buf_8 output712 (.A(net712),
    .X(la_data_in_mprj[94]));
 sky130_fd_sc_hd__buf_8 output713 (.A(net713),
    .X(la_data_in_mprj[95]));
 sky130_fd_sc_hd__buf_8 output714 (.A(net714),
    .X(la_data_in_mprj[96]));
 sky130_fd_sc_hd__buf_8 output715 (.A(net715),
    .X(la_data_in_mprj[97]));
 sky130_fd_sc_hd__buf_8 output716 (.A(net716),
    .X(la_data_in_mprj[98]));
 sky130_fd_sc_hd__buf_8 output717 (.A(net717),
    .X(la_data_in_mprj[99]));
 sky130_fd_sc_hd__buf_8 output718 (.A(net718),
    .X(la_data_in_mprj[9]));
 sky130_fd_sc_hd__buf_8 output719 (.A(net719),
    .X(la_oenb_core[0]));
 sky130_fd_sc_hd__buf_8 output720 (.A(net720),
    .X(la_oenb_core[100]));
 sky130_fd_sc_hd__buf_8 output721 (.A(net721),
    .X(la_oenb_core[101]));
 sky130_fd_sc_hd__buf_8 output722 (.A(net722),
    .X(la_oenb_core[102]));
 sky130_fd_sc_hd__buf_8 output723 (.A(net723),
    .X(la_oenb_core[103]));
 sky130_fd_sc_hd__buf_8 output724 (.A(net724),
    .X(la_oenb_core[104]));
 sky130_fd_sc_hd__buf_8 output725 (.A(net725),
    .X(la_oenb_core[105]));
 sky130_fd_sc_hd__buf_8 output726 (.A(net726),
    .X(la_oenb_core[106]));
 sky130_fd_sc_hd__buf_8 output727 (.A(net727),
    .X(la_oenb_core[107]));
 sky130_fd_sc_hd__buf_8 output728 (.A(net728),
    .X(la_oenb_core[108]));
 sky130_fd_sc_hd__buf_8 output729 (.A(net729),
    .X(la_oenb_core[109]));
 sky130_fd_sc_hd__buf_8 output730 (.A(net730),
    .X(la_oenb_core[10]));
 sky130_fd_sc_hd__buf_8 output731 (.A(net731),
    .X(la_oenb_core[110]));
 sky130_fd_sc_hd__buf_8 output732 (.A(net732),
    .X(la_oenb_core[111]));
 sky130_fd_sc_hd__buf_8 output733 (.A(net733),
    .X(la_oenb_core[112]));
 sky130_fd_sc_hd__buf_8 output734 (.A(net734),
    .X(la_oenb_core[113]));
 sky130_fd_sc_hd__buf_8 output735 (.A(net735),
    .X(la_oenb_core[114]));
 sky130_fd_sc_hd__buf_8 output736 (.A(net736),
    .X(la_oenb_core[115]));
 sky130_fd_sc_hd__buf_8 output737 (.A(net737),
    .X(la_oenb_core[116]));
 sky130_fd_sc_hd__buf_8 output738 (.A(net738),
    .X(la_oenb_core[117]));
 sky130_fd_sc_hd__buf_8 output739 (.A(net739),
    .X(la_oenb_core[118]));
 sky130_fd_sc_hd__buf_8 output740 (.A(net740),
    .X(la_oenb_core[119]));
 sky130_fd_sc_hd__buf_8 output741 (.A(net741),
    .X(la_oenb_core[11]));
 sky130_fd_sc_hd__buf_8 output742 (.A(net742),
    .X(la_oenb_core[120]));
 sky130_fd_sc_hd__buf_8 output743 (.A(net743),
    .X(la_oenb_core[121]));
 sky130_fd_sc_hd__buf_8 output744 (.A(net744),
    .X(la_oenb_core[122]));
 sky130_fd_sc_hd__buf_8 output745 (.A(net745),
    .X(la_oenb_core[123]));
 sky130_fd_sc_hd__buf_8 output746 (.A(net746),
    .X(la_oenb_core[124]));
 sky130_fd_sc_hd__buf_8 output747 (.A(net747),
    .X(la_oenb_core[125]));
 sky130_fd_sc_hd__buf_8 output748 (.A(net748),
    .X(la_oenb_core[126]));
 sky130_fd_sc_hd__buf_8 output749 (.A(net749),
    .X(la_oenb_core[127]));
 sky130_fd_sc_hd__buf_8 output750 (.A(net750),
    .X(la_oenb_core[12]));
 sky130_fd_sc_hd__buf_8 output751 (.A(net751),
    .X(la_oenb_core[13]));
 sky130_fd_sc_hd__buf_8 output752 (.A(net752),
    .X(la_oenb_core[14]));
 sky130_fd_sc_hd__buf_8 output753 (.A(net753),
    .X(la_oenb_core[15]));
 sky130_fd_sc_hd__buf_8 output754 (.A(net754),
    .X(la_oenb_core[16]));
 sky130_fd_sc_hd__buf_8 output755 (.A(net755),
    .X(la_oenb_core[17]));
 sky130_fd_sc_hd__buf_8 output756 (.A(net756),
    .X(la_oenb_core[18]));
 sky130_fd_sc_hd__buf_8 output757 (.A(net757),
    .X(la_oenb_core[19]));
 sky130_fd_sc_hd__buf_8 output758 (.A(net758),
    .X(la_oenb_core[1]));
 sky130_fd_sc_hd__buf_8 output759 (.A(net759),
    .X(la_oenb_core[20]));
 sky130_fd_sc_hd__buf_8 output760 (.A(net760),
    .X(la_oenb_core[21]));
 sky130_fd_sc_hd__buf_8 output761 (.A(net761),
    .X(la_oenb_core[22]));
 sky130_fd_sc_hd__buf_8 output762 (.A(net762),
    .X(la_oenb_core[23]));
 sky130_fd_sc_hd__buf_8 output763 (.A(net763),
    .X(la_oenb_core[24]));
 sky130_fd_sc_hd__buf_8 output764 (.A(net764),
    .X(la_oenb_core[25]));
 sky130_fd_sc_hd__buf_8 output765 (.A(net765),
    .X(la_oenb_core[26]));
 sky130_fd_sc_hd__buf_8 output766 (.A(net766),
    .X(la_oenb_core[27]));
 sky130_fd_sc_hd__buf_8 output767 (.A(net767),
    .X(la_oenb_core[28]));
 sky130_fd_sc_hd__buf_8 output768 (.A(net768),
    .X(la_oenb_core[29]));
 sky130_fd_sc_hd__buf_8 output769 (.A(net769),
    .X(la_oenb_core[2]));
 sky130_fd_sc_hd__buf_8 output770 (.A(net770),
    .X(la_oenb_core[30]));
 sky130_fd_sc_hd__buf_8 output771 (.A(net771),
    .X(la_oenb_core[31]));
 sky130_fd_sc_hd__buf_8 output772 (.A(net772),
    .X(la_oenb_core[32]));
 sky130_fd_sc_hd__buf_8 output773 (.A(net773),
    .X(la_oenb_core[33]));
 sky130_fd_sc_hd__buf_8 output774 (.A(net774),
    .X(la_oenb_core[34]));
 sky130_fd_sc_hd__buf_8 output775 (.A(net775),
    .X(la_oenb_core[35]));
 sky130_fd_sc_hd__buf_8 output776 (.A(net776),
    .X(la_oenb_core[36]));
 sky130_fd_sc_hd__buf_8 output777 (.A(net777),
    .X(la_oenb_core[37]));
 sky130_fd_sc_hd__buf_8 output778 (.A(net778),
    .X(la_oenb_core[38]));
 sky130_fd_sc_hd__buf_8 output779 (.A(net779),
    .X(la_oenb_core[39]));
 sky130_fd_sc_hd__buf_8 output780 (.A(net780),
    .X(la_oenb_core[3]));
 sky130_fd_sc_hd__buf_8 output781 (.A(net781),
    .X(la_oenb_core[40]));
 sky130_fd_sc_hd__buf_8 output782 (.A(net782),
    .X(la_oenb_core[41]));
 sky130_fd_sc_hd__buf_8 output783 (.A(net783),
    .X(la_oenb_core[42]));
 sky130_fd_sc_hd__buf_8 output784 (.A(net784),
    .X(la_oenb_core[43]));
 sky130_fd_sc_hd__buf_8 output785 (.A(net785),
    .X(la_oenb_core[44]));
 sky130_fd_sc_hd__buf_8 output786 (.A(net786),
    .X(la_oenb_core[45]));
 sky130_fd_sc_hd__buf_8 output787 (.A(net787),
    .X(la_oenb_core[46]));
 sky130_fd_sc_hd__buf_8 output788 (.A(net788),
    .X(la_oenb_core[47]));
 sky130_fd_sc_hd__buf_8 output789 (.A(net789),
    .X(la_oenb_core[48]));
 sky130_fd_sc_hd__buf_8 output790 (.A(net790),
    .X(la_oenb_core[49]));
 sky130_fd_sc_hd__buf_8 output791 (.A(net791),
    .X(la_oenb_core[4]));
 sky130_fd_sc_hd__buf_8 output792 (.A(net792),
    .X(la_oenb_core[50]));
 sky130_fd_sc_hd__buf_8 output793 (.A(net793),
    .X(la_oenb_core[51]));
 sky130_fd_sc_hd__buf_8 output794 (.A(net794),
    .X(la_oenb_core[52]));
 sky130_fd_sc_hd__buf_8 output795 (.A(net795),
    .X(la_oenb_core[53]));
 sky130_fd_sc_hd__buf_8 output796 (.A(net796),
    .X(la_oenb_core[54]));
 sky130_fd_sc_hd__buf_8 output797 (.A(net797),
    .X(la_oenb_core[55]));
 sky130_fd_sc_hd__buf_8 output798 (.A(net798),
    .X(la_oenb_core[56]));
 sky130_fd_sc_hd__buf_8 output799 (.A(net799),
    .X(la_oenb_core[57]));
 sky130_fd_sc_hd__buf_8 output800 (.A(net800),
    .X(la_oenb_core[58]));
 sky130_fd_sc_hd__buf_8 output801 (.A(net801),
    .X(la_oenb_core[59]));
 sky130_fd_sc_hd__buf_8 output802 (.A(net802),
    .X(la_oenb_core[5]));
 sky130_fd_sc_hd__buf_8 output803 (.A(net803),
    .X(la_oenb_core[60]));
 sky130_fd_sc_hd__buf_8 output804 (.A(net804),
    .X(la_oenb_core[61]));
 sky130_fd_sc_hd__buf_8 output805 (.A(net805),
    .X(la_oenb_core[62]));
 sky130_fd_sc_hd__buf_8 output806 (.A(net806),
    .X(la_oenb_core[63]));
 sky130_fd_sc_hd__buf_8 output807 (.A(net807),
    .X(la_oenb_core[64]));
 sky130_fd_sc_hd__buf_8 output808 (.A(net808),
    .X(la_oenb_core[65]));
 sky130_fd_sc_hd__buf_8 output809 (.A(net809),
    .X(la_oenb_core[66]));
 sky130_fd_sc_hd__buf_8 output810 (.A(net810),
    .X(la_oenb_core[67]));
 sky130_fd_sc_hd__buf_8 output811 (.A(net811),
    .X(la_oenb_core[68]));
 sky130_fd_sc_hd__buf_8 output812 (.A(net812),
    .X(la_oenb_core[69]));
 sky130_fd_sc_hd__buf_8 output813 (.A(net813),
    .X(la_oenb_core[6]));
 sky130_fd_sc_hd__buf_8 output814 (.A(net814),
    .X(la_oenb_core[70]));
 sky130_fd_sc_hd__buf_8 output815 (.A(net815),
    .X(la_oenb_core[71]));
 sky130_fd_sc_hd__buf_8 output816 (.A(net816),
    .X(la_oenb_core[72]));
 sky130_fd_sc_hd__buf_8 output817 (.A(net817),
    .X(la_oenb_core[73]));
 sky130_fd_sc_hd__buf_8 output818 (.A(net818),
    .X(la_oenb_core[74]));
 sky130_fd_sc_hd__buf_8 output819 (.A(net819),
    .X(la_oenb_core[75]));
 sky130_fd_sc_hd__buf_8 output820 (.A(net820),
    .X(la_oenb_core[76]));
 sky130_fd_sc_hd__buf_8 output821 (.A(net821),
    .X(la_oenb_core[77]));
 sky130_fd_sc_hd__buf_8 output822 (.A(net822),
    .X(la_oenb_core[78]));
 sky130_fd_sc_hd__buf_8 output823 (.A(net823),
    .X(la_oenb_core[79]));
 sky130_fd_sc_hd__buf_8 output824 (.A(net824),
    .X(la_oenb_core[7]));
 sky130_fd_sc_hd__buf_8 output825 (.A(net825),
    .X(la_oenb_core[80]));
 sky130_fd_sc_hd__buf_8 output826 (.A(net826),
    .X(la_oenb_core[81]));
 sky130_fd_sc_hd__buf_8 output827 (.A(net827),
    .X(la_oenb_core[82]));
 sky130_fd_sc_hd__buf_8 output828 (.A(net828),
    .X(la_oenb_core[83]));
 sky130_fd_sc_hd__buf_8 output829 (.A(net829),
    .X(la_oenb_core[84]));
 sky130_fd_sc_hd__buf_8 output830 (.A(net830),
    .X(la_oenb_core[85]));
 sky130_fd_sc_hd__buf_8 output831 (.A(net831),
    .X(la_oenb_core[86]));
 sky130_fd_sc_hd__buf_8 output832 (.A(net832),
    .X(la_oenb_core[87]));
 sky130_fd_sc_hd__buf_8 output833 (.A(net833),
    .X(la_oenb_core[88]));
 sky130_fd_sc_hd__buf_8 output834 (.A(net834),
    .X(la_oenb_core[89]));
 sky130_fd_sc_hd__buf_8 output835 (.A(net835),
    .X(la_oenb_core[8]));
 sky130_fd_sc_hd__buf_8 output836 (.A(net836),
    .X(la_oenb_core[90]));
 sky130_fd_sc_hd__buf_8 output837 (.A(net837),
    .X(la_oenb_core[91]));
 sky130_fd_sc_hd__buf_8 output838 (.A(net838),
    .X(la_oenb_core[92]));
 sky130_fd_sc_hd__buf_8 output839 (.A(net839),
    .X(la_oenb_core[93]));
 sky130_fd_sc_hd__buf_8 output840 (.A(net840),
    .X(la_oenb_core[94]));
 sky130_fd_sc_hd__buf_8 output841 (.A(net841),
    .X(la_oenb_core[95]));
 sky130_fd_sc_hd__buf_8 output842 (.A(net842),
    .X(la_oenb_core[96]));
 sky130_fd_sc_hd__buf_8 output843 (.A(net843),
    .X(la_oenb_core[97]));
 sky130_fd_sc_hd__buf_8 output844 (.A(net844),
    .X(la_oenb_core[98]));
 sky130_fd_sc_hd__buf_8 output845 (.A(net845),
    .X(la_oenb_core[99]));
 sky130_fd_sc_hd__buf_8 output846 (.A(net846),
    .X(la_oenb_core[9]));
 sky130_fd_sc_hd__buf_8 output847 (.A(net847),
    .X(mprj_ack_i_core));
 sky130_fd_sc_hd__buf_8 output848 (.A(net848),
    .X(mprj_adr_o_user[0]));
 sky130_fd_sc_hd__buf_8 output849 (.A(net849),
    .X(mprj_adr_o_user[10]));
 sky130_fd_sc_hd__buf_8 output850 (.A(net850),
    .X(mprj_adr_o_user[11]));
 sky130_fd_sc_hd__buf_8 output851 (.A(net851),
    .X(mprj_adr_o_user[12]));
 sky130_fd_sc_hd__buf_8 output852 (.A(net852),
    .X(mprj_adr_o_user[13]));
 sky130_fd_sc_hd__buf_8 output853 (.A(net853),
    .X(mprj_adr_o_user[14]));
 sky130_fd_sc_hd__buf_8 output854 (.A(net854),
    .X(mprj_adr_o_user[15]));
 sky130_fd_sc_hd__buf_8 output855 (.A(net855),
    .X(mprj_adr_o_user[16]));
 sky130_fd_sc_hd__buf_8 output856 (.A(net856),
    .X(mprj_adr_o_user[17]));
 sky130_fd_sc_hd__buf_8 output857 (.A(net857),
    .X(mprj_adr_o_user[18]));
 sky130_fd_sc_hd__buf_8 output858 (.A(net858),
    .X(mprj_adr_o_user[19]));
 sky130_fd_sc_hd__buf_8 output859 (.A(net859),
    .X(mprj_adr_o_user[1]));
 sky130_fd_sc_hd__buf_8 output860 (.A(net860),
    .X(mprj_adr_o_user[20]));
 sky130_fd_sc_hd__buf_8 output861 (.A(net861),
    .X(mprj_adr_o_user[21]));
 sky130_fd_sc_hd__buf_8 output862 (.A(net862),
    .X(mprj_adr_o_user[22]));
 sky130_fd_sc_hd__buf_8 output863 (.A(net863),
    .X(mprj_adr_o_user[23]));
 sky130_fd_sc_hd__buf_8 output864 (.A(net864),
    .X(mprj_adr_o_user[24]));
 sky130_fd_sc_hd__buf_8 output865 (.A(net865),
    .X(mprj_adr_o_user[25]));
 sky130_fd_sc_hd__buf_8 output866 (.A(net866),
    .X(mprj_adr_o_user[26]));
 sky130_fd_sc_hd__buf_8 output867 (.A(net867),
    .X(mprj_adr_o_user[27]));
 sky130_fd_sc_hd__buf_8 output868 (.A(net868),
    .X(mprj_adr_o_user[28]));
 sky130_fd_sc_hd__buf_8 output869 (.A(net869),
    .X(mprj_adr_o_user[29]));
 sky130_fd_sc_hd__buf_8 output870 (.A(net870),
    .X(mprj_adr_o_user[2]));
 sky130_fd_sc_hd__buf_8 output871 (.A(net871),
    .X(mprj_adr_o_user[30]));
 sky130_fd_sc_hd__buf_8 output872 (.A(net872),
    .X(mprj_adr_o_user[31]));
 sky130_fd_sc_hd__buf_8 output873 (.A(net873),
    .X(mprj_adr_o_user[3]));
 sky130_fd_sc_hd__buf_8 output874 (.A(net874),
    .X(mprj_adr_o_user[4]));
 sky130_fd_sc_hd__buf_8 output875 (.A(net875),
    .X(mprj_adr_o_user[5]));
 sky130_fd_sc_hd__buf_8 output876 (.A(net876),
    .X(mprj_adr_o_user[6]));
 sky130_fd_sc_hd__buf_8 output877 (.A(net877),
    .X(mprj_adr_o_user[7]));
 sky130_fd_sc_hd__buf_8 output878 (.A(net878),
    .X(mprj_adr_o_user[8]));
 sky130_fd_sc_hd__buf_8 output879 (.A(net879),
    .X(mprj_adr_o_user[9]));
 sky130_fd_sc_hd__buf_8 output880 (.A(net880),
    .X(mprj_cyc_o_user));
 sky130_fd_sc_hd__buf_8 output881 (.A(net881),
    .X(mprj_dat_i_core[0]));
 sky130_fd_sc_hd__buf_8 output882 (.A(net882),
    .X(mprj_dat_i_core[10]));
 sky130_fd_sc_hd__buf_8 output883 (.A(net883),
    .X(mprj_dat_i_core[11]));
 sky130_fd_sc_hd__buf_8 output884 (.A(net884),
    .X(mprj_dat_i_core[12]));
 sky130_fd_sc_hd__buf_8 output885 (.A(net885),
    .X(mprj_dat_i_core[13]));
 sky130_fd_sc_hd__buf_8 output886 (.A(net886),
    .X(mprj_dat_i_core[14]));
 sky130_fd_sc_hd__buf_8 output887 (.A(net887),
    .X(mprj_dat_i_core[15]));
 sky130_fd_sc_hd__buf_8 output888 (.A(net888),
    .X(mprj_dat_i_core[16]));
 sky130_fd_sc_hd__buf_8 output889 (.A(net889),
    .X(mprj_dat_i_core[17]));
 sky130_fd_sc_hd__buf_8 output890 (.A(net890),
    .X(mprj_dat_i_core[18]));
 sky130_fd_sc_hd__buf_8 output891 (.A(net891),
    .X(mprj_dat_i_core[19]));
 sky130_fd_sc_hd__buf_8 output892 (.A(net892),
    .X(mprj_dat_i_core[1]));
 sky130_fd_sc_hd__buf_8 output893 (.A(net893),
    .X(mprj_dat_i_core[20]));
 sky130_fd_sc_hd__buf_8 output894 (.A(net894),
    .X(mprj_dat_i_core[21]));
 sky130_fd_sc_hd__buf_8 output895 (.A(net895),
    .X(mprj_dat_i_core[22]));
 sky130_fd_sc_hd__buf_8 output896 (.A(net896),
    .X(mprj_dat_i_core[23]));
 sky130_fd_sc_hd__buf_8 output897 (.A(net897),
    .X(mprj_dat_i_core[24]));
 sky130_fd_sc_hd__buf_8 output898 (.A(net898),
    .X(mprj_dat_i_core[25]));
 sky130_fd_sc_hd__buf_8 output899 (.A(net899),
    .X(mprj_dat_i_core[26]));
 sky130_fd_sc_hd__buf_8 output900 (.A(net900),
    .X(mprj_dat_i_core[27]));
 sky130_fd_sc_hd__buf_8 output901 (.A(net901),
    .X(mprj_dat_i_core[28]));
 sky130_fd_sc_hd__buf_8 output902 (.A(net902),
    .X(mprj_dat_i_core[29]));
 sky130_fd_sc_hd__buf_8 output903 (.A(net903),
    .X(mprj_dat_i_core[2]));
 sky130_fd_sc_hd__buf_8 output904 (.A(net904),
    .X(mprj_dat_i_core[30]));
 sky130_fd_sc_hd__buf_8 output905 (.A(net905),
    .X(mprj_dat_i_core[31]));
 sky130_fd_sc_hd__buf_8 output906 (.A(net906),
    .X(mprj_dat_i_core[3]));
 sky130_fd_sc_hd__buf_8 output907 (.A(net907),
    .X(mprj_dat_i_core[4]));
 sky130_fd_sc_hd__buf_8 output908 (.A(net908),
    .X(mprj_dat_i_core[5]));
 sky130_fd_sc_hd__buf_8 output909 (.A(net909),
    .X(mprj_dat_i_core[6]));
 sky130_fd_sc_hd__buf_8 output910 (.A(net910),
    .X(mprj_dat_i_core[7]));
 sky130_fd_sc_hd__buf_8 output911 (.A(net911),
    .X(mprj_dat_i_core[8]));
 sky130_fd_sc_hd__buf_8 output912 (.A(net912),
    .X(mprj_dat_i_core[9]));
 sky130_fd_sc_hd__buf_8 output913 (.A(net913),
    .X(mprj_dat_o_user[0]));
 sky130_fd_sc_hd__buf_8 output914 (.A(net914),
    .X(mprj_dat_o_user[10]));
 sky130_fd_sc_hd__buf_8 output915 (.A(net915),
    .X(mprj_dat_o_user[11]));
 sky130_fd_sc_hd__buf_8 output916 (.A(net916),
    .X(mprj_dat_o_user[12]));
 sky130_fd_sc_hd__buf_8 output917 (.A(net917),
    .X(mprj_dat_o_user[13]));
 sky130_fd_sc_hd__buf_8 output918 (.A(net918),
    .X(mprj_dat_o_user[14]));
 sky130_fd_sc_hd__buf_8 output919 (.A(net919),
    .X(mprj_dat_o_user[15]));
 sky130_fd_sc_hd__buf_8 output920 (.A(net920),
    .X(mprj_dat_o_user[16]));
 sky130_fd_sc_hd__buf_8 output921 (.A(net921),
    .X(mprj_dat_o_user[17]));
 sky130_fd_sc_hd__buf_8 output922 (.A(net922),
    .X(mprj_dat_o_user[18]));
 sky130_fd_sc_hd__buf_8 output923 (.A(net923),
    .X(mprj_dat_o_user[19]));
 sky130_fd_sc_hd__buf_8 output924 (.A(net924),
    .X(mprj_dat_o_user[1]));
 sky130_fd_sc_hd__buf_8 output925 (.A(net925),
    .X(mprj_dat_o_user[20]));
 sky130_fd_sc_hd__buf_8 output926 (.A(net926),
    .X(mprj_dat_o_user[21]));
 sky130_fd_sc_hd__buf_8 output927 (.A(net927),
    .X(mprj_dat_o_user[22]));
 sky130_fd_sc_hd__buf_8 output928 (.A(net928),
    .X(mprj_dat_o_user[23]));
 sky130_fd_sc_hd__buf_8 output929 (.A(net929),
    .X(mprj_dat_o_user[24]));
 sky130_fd_sc_hd__buf_8 output930 (.A(net930),
    .X(mprj_dat_o_user[25]));
 sky130_fd_sc_hd__buf_8 output931 (.A(net931),
    .X(mprj_dat_o_user[26]));
 sky130_fd_sc_hd__buf_8 output932 (.A(net932),
    .X(mprj_dat_o_user[27]));
 sky130_fd_sc_hd__buf_8 output933 (.A(net933),
    .X(mprj_dat_o_user[28]));
 sky130_fd_sc_hd__buf_8 output934 (.A(net934),
    .X(mprj_dat_o_user[29]));
 sky130_fd_sc_hd__buf_8 output935 (.A(net935),
    .X(mprj_dat_o_user[2]));
 sky130_fd_sc_hd__buf_8 output936 (.A(net936),
    .X(mprj_dat_o_user[30]));
 sky130_fd_sc_hd__buf_8 output937 (.A(net937),
    .X(mprj_dat_o_user[31]));
 sky130_fd_sc_hd__buf_8 output938 (.A(net938),
    .X(mprj_dat_o_user[3]));
 sky130_fd_sc_hd__buf_8 output939 (.A(net939),
    .X(mprj_dat_o_user[4]));
 sky130_fd_sc_hd__buf_8 output940 (.A(net940),
    .X(mprj_dat_o_user[5]));
 sky130_fd_sc_hd__buf_8 output941 (.A(net941),
    .X(mprj_dat_o_user[6]));
 sky130_fd_sc_hd__buf_8 output942 (.A(net942),
    .X(mprj_dat_o_user[7]));
 sky130_fd_sc_hd__buf_8 output943 (.A(net943),
    .X(mprj_dat_o_user[8]));
 sky130_fd_sc_hd__buf_8 output944 (.A(net944),
    .X(mprj_dat_o_user[9]));
 sky130_fd_sc_hd__buf_8 output945 (.A(net945),
    .X(mprj_sel_o_user[0]));
 sky130_fd_sc_hd__buf_8 output946 (.A(net946),
    .X(mprj_sel_o_user[1]));
 sky130_fd_sc_hd__buf_8 output947 (.A(net947),
    .X(mprj_sel_o_user[2]));
 sky130_fd_sc_hd__buf_8 output948 (.A(net948),
    .X(mprj_sel_o_user[3]));
 sky130_fd_sc_hd__buf_8 output949 (.A(net949),
    .X(mprj_stb_o_user));
 sky130_fd_sc_hd__buf_8 output950 (.A(net950),
    .X(mprj_we_o_user));
 sky130_fd_sc_hd__buf_8 output951 (.A(net951),
    .X(user1_vcc_powergood));
 sky130_fd_sc_hd__buf_8 output952 (.A(net952),
    .X(user1_vdd_powergood));
 sky130_fd_sc_hd__buf_8 output953 (.A(net953),
    .X(user2_vcc_powergood));
 sky130_fd_sc_hd__buf_8 output954 (.A(net954),
    .X(user2_vdd_powergood));
 sky130_fd_sc_hd__buf_8 output955 (.A(net955),
    .X(user_clock));
 sky130_fd_sc_hd__buf_8 output956 (.A(net956),
    .X(user_clock2));
 sky130_fd_sc_hd__buf_8 output957 (.A(net957),
    .X(user_irq[0]));
 sky130_fd_sc_hd__buf_8 output958 (.A(net958),
    .X(user_irq[1]));
 sky130_fd_sc_hd__buf_8 output959 (.A(net959),
    .X(user_irq[2]));
 sky130_fd_sc_hd__buf_8 output960 (.A(net960),
    .X(user_reset));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(\la_data_in_mprj_bar[100] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(\la_data_in_mprj_bar[101] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(\la_data_in_mprj_bar[88] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(\la_data_in_mprj_bar[89] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(la_data_out_core[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(la_data_out_core[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(la_data_out_core[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(la_data_out_core[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(la_data_out_core[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(la_data_out_core[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(la_data_out_core[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(la_data_out_core[33]));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(la_data_out_core[33]));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(la_data_out_core[40]));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(la_data_out_core[41]));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(mprj_ack_i_user));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(mprj_ack_i_user));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(mprj_ack_i_user));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(mprj_ack_i_user));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(mprj_ack_i_user));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(mprj_ack_i_user));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(mprj_ack_i_user));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(mprj_ack_i_user));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(mprj_ack_i_user));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(mprj_ack_i_user));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(mprj_ack_i_user));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(mprj_dat_i_user[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(mprj_dat_i_user[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(mprj_dat_i_user[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(mprj_dat_i_user[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(mprj_dat_i_user[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(mprj_dat_i_user[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(mprj_dat_i_user[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(mprj_dat_i_user[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(mprj_dat_i_user[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(mprj_dat_i_user[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(mprj_dat_i_user[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(mprj_dat_i_user[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(mprj_dat_i_user[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(mprj_dat_i_user[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(mprj_dat_i_user[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(mprj_dat_i_user[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(mprj_dat_i_user[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(mprj_dat_i_user[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(mprj_dat_i_user[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(mprj_dat_i_user[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(mprj_dat_i_user[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(mprj_dat_i_user[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(mprj_dat_i_user[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(mprj_dat_i_user[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(mprj_dat_i_user[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(mprj_dat_i_user[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(mprj_dat_i_user[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(mprj_dat_i_user[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(mprj_dat_i_user[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(mprj_dat_i_user[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(mprj_dat_i_user[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(mprj_dat_i_user[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(mprj_dat_i_user[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(mprj_dat_i_user[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(mprj_dat_i_user[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(mprj_dat_i_user[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(mprj_dat_i_user[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(mprj_dat_i_user[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(mprj_dat_i_user[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(mprj_dat_i_user[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(mprj_dat_i_user[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(mprj_dat_i_user[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(mprj_dat_i_user[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(mprj_dat_i_user[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(mprj_dat_i_user[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(mprj_dat_i_user[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(mprj_dat_i_user[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(mprj_dat_i_user[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(mprj_dat_i_user[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(mprj_dat_i_user[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(mprj_dat_i_user[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(mprj_dat_i_user[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(mprj_dat_i_user[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(mprj_dat_i_user[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(mprj_dat_i_user[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(mprj_dat_i_user[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(mprj_dat_i_user[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(mprj_dat_i_user[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(mprj_dat_i_user[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(mprj_dat_i_user[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(mprj_dat_i_user[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(mprj_dat_i_user[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(mprj_dat_i_user[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(mprj_dat_i_user[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(mprj_dat_i_user[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(mprj_dat_i_user[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(mprj_dat_i_user[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(mprj_dat_i_user[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(mprj_dat_i_user[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(mprj_dat_i_user[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(mprj_dat_i_user[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(mprj_dat_i_user[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(mprj_dat_i_user[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(mprj_dat_i_user[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(mprj_dat_i_user[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(mprj_dat_i_user[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(mprj_dat_i_user[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(mprj_dat_i_user[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(mprj_dat_i_user[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(mprj_dat_i_user[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(mprj_dat_i_user[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(mprj_dat_i_user[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(mprj_dat_i_user[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(mprj_dat_i_user[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(mprj_dat_i_user[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(mprj_dat_i_user[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(mprj_dat_i_user[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(mprj_dat_i_user[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(mprj_dat_i_user[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(mprj_dat_i_user[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(mprj_dat_i_user[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(mprj_dat_i_user[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(mprj_dat_i_user[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(mprj_dat_i_user[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(mprj_dat_i_user[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(mprj_dat_i_user[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(mprj_dat_i_user[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(mprj_dat_i_user[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(mprj_dat_i_user[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(mprj_dat_i_user[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(mprj_dat_i_user[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(mprj_dat_i_user[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(mprj_dat_i_user[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(mprj_dat_i_user[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(mprj_dat_i_user[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(mprj_dat_i_user[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(mprj_dat_i_user[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(mprj_dat_i_user[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(mprj_dat_i_user[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(mprj_dat_i_user[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_137 (.DIODE(mprj_dat_i_user[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_138 (.DIODE(mprj_dat_i_user[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_139 (.DIODE(mprj_dat_i_user[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_140 (.DIODE(mprj_dat_i_user[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_141 (.DIODE(mprj_dat_i_user[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_142 (.DIODE(mprj_dat_i_user[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_143 (.DIODE(mprj_dat_i_user[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_144 (.DIODE(mprj_dat_i_user[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_145 (.DIODE(mprj_dat_i_user[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_146 (.DIODE(mprj_dat_i_user[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_147 (.DIODE(mprj_dat_i_user[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_148 (.DIODE(mprj_dat_i_user[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_149 (.DIODE(mprj_dat_i_user[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_150 (.DIODE(mprj_dat_i_user[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_151 (.DIODE(mprj_dat_i_user[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_152 (.DIODE(mprj_dat_i_user[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_153 (.DIODE(mprj_dat_i_user[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_154 (.DIODE(mprj_dat_i_user[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_155 (.DIODE(mprj_dat_i_user[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_156 (.DIODE(mprj_dat_i_user[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_157 (.DIODE(mprj_dat_i_user[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_158 (.DIODE(mprj_dat_i_user[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_159 (.DIODE(mprj_dat_i_user[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_160 (.DIODE(mprj_dat_i_user[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_161 (.DIODE(mprj_dat_i_user[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_162 (.DIODE(mprj_dat_i_user[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_163 (.DIODE(mprj_dat_i_user[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_164 (.DIODE(mprj_dat_i_user[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_165 (.DIODE(mprj_dat_i_user[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_166 (.DIODE(mprj_dat_i_user[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_167 (.DIODE(mprj_dat_i_user[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_168 (.DIODE(mprj_dat_i_user[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_169 (.DIODE(mprj_dat_i_user[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_170 (.DIODE(mprj_dat_i_user[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_171 (.DIODE(mprj_dat_i_user[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_172 (.DIODE(mprj_dat_i_user[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_173 (.DIODE(mprj_dat_i_user[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_174 (.DIODE(mprj_dat_i_user[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_175 (.DIODE(mprj_dat_i_user[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_176 (.DIODE(mprj_dat_i_user[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_177 (.DIODE(mprj_dat_i_user[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_178 (.DIODE(mprj_dat_i_user[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_179 (.DIODE(mprj_dat_i_user[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_180 (.DIODE(mprj_dat_i_user[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_181 (.DIODE(mprj_dat_i_user[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_182 (.DIODE(mprj_dat_i_user[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_183 (.DIODE(mprj_dat_i_user[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_184 (.DIODE(mprj_dat_i_user[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_185 (.DIODE(mprj_dat_i_user[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_186 (.DIODE(mprj_dat_i_user[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_187 (.DIODE(mprj_dat_i_user[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_188 (.DIODE(mprj_dat_i_user[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_189 (.DIODE(mprj_dat_i_user[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_190 (.DIODE(mprj_dat_i_user[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_191 (.DIODE(mprj_dat_i_user[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_192 (.DIODE(mprj_dat_i_user[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_193 (.DIODE(mprj_dat_i_user[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_194 (.DIODE(mprj_dat_i_user[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_195 (.DIODE(mprj_dat_i_user[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_196 (.DIODE(mprj_dat_i_user[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_197 (.DIODE(mprj_dat_i_user[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_198 (.DIODE(\mprj_logic1[101] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_199 (.DIODE(\mprj_logic1[103] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_200 (.DIODE(\mprj_logic1[103] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_201 (.DIODE(\mprj_logic1[117] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_202 (.DIODE(\mprj_logic1[128] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_203 (.DIODE(\mprj_logic1[128] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_204 (.DIODE(\mprj_logic1[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_205 (.DIODE(\mprj_logic1[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_206 (.DIODE(\mprj_logic1[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_207 (.DIODE(\mprj_logic1[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_208 (.DIODE(\mprj_logic1[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_209 (.DIODE(\mprj_logic1[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_210 (.DIODE(\mprj_logic1[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_211 (.DIODE(\mprj_logic1[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_212 (.DIODE(\mprj_logic1[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_213 (.DIODE(\mprj_logic1[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_214 (.DIODE(\mprj_logic1[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_215 (.DIODE(\mprj_logic1[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_216 (.DIODE(\mprj_logic1[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_217 (.DIODE(\mprj_logic1[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_218 (.DIODE(\mprj_logic1[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_219 (.DIODE(\mprj_logic1[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_220 (.DIODE(\mprj_logic1[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_221 (.DIODE(\mprj_logic1[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_222 (.DIODE(\mprj_logic1[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_223 (.DIODE(\mprj_logic1[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_224 (.DIODE(\mprj_logic1[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_225 (.DIODE(\mprj_logic1[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_226 (.DIODE(\mprj_logic1[130] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_227 (.DIODE(\mprj_logic1[130] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_228 (.DIODE(\mprj_logic1[134] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_229 (.DIODE(\mprj_logic1[135] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_230 (.DIODE(\mprj_logic1[139] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_231 (.DIODE(\mprj_logic1[139] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_232 (.DIODE(\mprj_logic1[139] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_233 (.DIODE(\mprj_logic1[139] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_234 (.DIODE(\mprj_logic1[139] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_235 (.DIODE(\mprj_logic1[139] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_236 (.DIODE(\mprj_logic1[140] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_237 (.DIODE(\mprj_logic1[140] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_238 (.DIODE(\mprj_logic1[140] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_239 (.DIODE(\mprj_logic1[140] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_240 (.DIODE(\mprj_logic1[140] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_241 (.DIODE(\mprj_logic1[140] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_242 (.DIODE(\mprj_logic1[145] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_243 (.DIODE(\mprj_logic1[145] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_244 (.DIODE(\mprj_logic1[145] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_245 (.DIODE(\mprj_logic1[145] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_246 (.DIODE(\mprj_logic1[145] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_247 (.DIODE(\mprj_logic1[145] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_248 (.DIODE(\mprj_logic1[145] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_249 (.DIODE(\mprj_logic1[145] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_250 (.DIODE(\mprj_logic1[145] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_251 (.DIODE(\mprj_logic1[145] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_252 (.DIODE(\mprj_logic1[146] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_253 (.DIODE(\mprj_logic1[146] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_254 (.DIODE(\mprj_logic1[146] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_255 (.DIODE(\mprj_logic1[146] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_256 (.DIODE(\mprj_logic1[146] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_257 (.DIODE(\mprj_logic1[146] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_258 (.DIODE(\mprj_logic1[148] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_259 (.DIODE(\mprj_logic1[150] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_260 (.DIODE(\mprj_logic1[150] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_261 (.DIODE(\mprj_logic1[150] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_262 (.DIODE(\mprj_logic1[150] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_263 (.DIODE(\mprj_logic1[150] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_264 (.DIODE(\mprj_logic1[152] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_265 (.DIODE(\mprj_logic1[152] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_266 (.DIODE(\mprj_logic1[152] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_267 (.DIODE(\mprj_logic1[152] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_268 (.DIODE(\mprj_logic1[152] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_269 (.DIODE(\mprj_logic1[152] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_270 (.DIODE(\mprj_logic1[153] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_271 (.DIODE(\mprj_logic1[153] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_272 (.DIODE(\mprj_logic1[153] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_273 (.DIODE(\mprj_logic1[153] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_274 (.DIODE(\mprj_logic1[153] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_275 (.DIODE(\mprj_logic1[153] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_276 (.DIODE(\mprj_logic1[153] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_277 (.DIODE(\mprj_logic1[153] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_278 (.DIODE(\mprj_logic1[154] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_279 (.DIODE(\mprj_logic1[154] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_280 (.DIODE(\mprj_logic1[154] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_281 (.DIODE(\mprj_logic1[154] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_282 (.DIODE(\mprj_logic1[154] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_283 (.DIODE(\mprj_logic1[156] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_284 (.DIODE(\mprj_logic1[156] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_285 (.DIODE(\mprj_logic1[156] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_286 (.DIODE(\mprj_logic1[156] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_287 (.DIODE(\mprj_logic1[156] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_288 (.DIODE(\mprj_logic1[156] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_289 (.DIODE(\mprj_logic1[156] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_290 (.DIODE(\mprj_logic1[156] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_291 (.DIODE(\mprj_logic1[156] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_292 (.DIODE(\mprj_logic1[156] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_293 (.DIODE(\mprj_logic1[156] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_294 (.DIODE(\mprj_logic1[156] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_295 (.DIODE(\mprj_logic1[156] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_296 (.DIODE(\mprj_logic1[156] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_297 (.DIODE(\mprj_logic1[156] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_298 (.DIODE(\mprj_logic1[156] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_299 (.DIODE(\mprj_logic1[156] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_300 (.DIODE(\mprj_logic1[156] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_301 (.DIODE(\mprj_logic1[157] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_302 (.DIODE(\mprj_logic1[157] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_303 (.DIODE(\mprj_logic1[157] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_304 (.DIODE(\mprj_logic1[157] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_305 (.DIODE(\mprj_logic1[157] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_306 (.DIODE(\mprj_logic1[157] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_307 (.DIODE(\mprj_logic1[157] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_308 (.DIODE(\mprj_logic1[157] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_309 (.DIODE(\mprj_logic1[157] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_310 (.DIODE(\mprj_logic1[157] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_311 (.DIODE(\mprj_logic1[157] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_312 (.DIODE(\mprj_logic1[157] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_313 (.DIODE(\mprj_logic1[157] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_314 (.DIODE(\mprj_logic1[157] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_315 (.DIODE(\mprj_logic1[157] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_316 (.DIODE(\mprj_logic1[157] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_317 (.DIODE(\mprj_logic1[157] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_318 (.DIODE(\mprj_logic1[157] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_319 (.DIODE(\mprj_logic1[158] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_320 (.DIODE(\mprj_logic1[158] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_321 (.DIODE(\mprj_logic1[158] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_322 (.DIODE(\mprj_logic1[158] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_323 (.DIODE(\mprj_logic1[158] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_324 (.DIODE(\mprj_logic1[158] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_325 (.DIODE(\mprj_logic1[158] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_326 (.DIODE(\mprj_logic1[158] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_327 (.DIODE(\mprj_logic1[158] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_328 (.DIODE(\mprj_logic1[158] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_329 (.DIODE(\mprj_logic1[158] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_330 (.DIODE(\mprj_logic1[159] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_331 (.DIODE(\mprj_logic1[159] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_332 (.DIODE(\mprj_logic1[159] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_333 (.DIODE(\mprj_logic1[159] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_334 (.DIODE(\mprj_logic1[159] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_335 (.DIODE(\mprj_logic1[159] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_336 (.DIODE(\mprj_logic1[159] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_337 (.DIODE(\mprj_logic1[159] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_338 (.DIODE(\mprj_logic1[159] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_339 (.DIODE(\mprj_logic1[159] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_340 (.DIODE(\mprj_logic1[159] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_341 (.DIODE(\mprj_logic1[159] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_342 (.DIODE(\mprj_logic1[159] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_343 (.DIODE(\mprj_logic1[159] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_344 (.DIODE(\mprj_logic1[159] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_345 (.DIODE(\mprj_logic1[159] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_346 (.DIODE(\mprj_logic1[159] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_347 (.DIODE(\mprj_logic1[159] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_348 (.DIODE(\mprj_logic1[159] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_349 (.DIODE(\mprj_logic1[159] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_350 (.DIODE(\mprj_logic1[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_351 (.DIODE(\mprj_logic1[161] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_352 (.DIODE(\mprj_logic1[161] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_353 (.DIODE(\mprj_logic1[161] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_354 (.DIODE(\mprj_logic1[161] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_355 (.DIODE(\mprj_logic1[161] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_356 (.DIODE(\mprj_logic1[161] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_357 (.DIODE(\mprj_logic1[161] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_358 (.DIODE(\mprj_logic1[161] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_359 (.DIODE(\mprj_logic1[161] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_360 (.DIODE(\mprj_logic1[161] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_361 (.DIODE(\mprj_logic1[161] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_362 (.DIODE(\mprj_logic1[161] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_363 (.DIODE(\mprj_logic1[161] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_364 (.DIODE(\mprj_logic1[161] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_365 (.DIODE(\mprj_logic1[161] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_366 (.DIODE(\mprj_logic1[161] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_367 (.DIODE(\mprj_logic1[161] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_368 (.DIODE(\mprj_logic1[161] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_369 (.DIODE(\mprj_logic1[161] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_370 (.DIODE(\mprj_logic1[161] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_371 (.DIODE(\mprj_logic1[161] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_372 (.DIODE(\mprj_logic1[161] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_373 (.DIODE(\mprj_logic1[162] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_374 (.DIODE(\mprj_logic1[162] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_375 (.DIODE(\mprj_logic1[162] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_376 (.DIODE(\mprj_logic1[170] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_377 (.DIODE(\mprj_logic1[171] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_378 (.DIODE(\mprj_logic1[171] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_379 (.DIODE(\mprj_logic1[173] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_380 (.DIODE(\mprj_logic1[174] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_381 (.DIODE(\mprj_logic1[175] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_382 (.DIODE(\mprj_logic1[177] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_383 (.DIODE(\mprj_logic1[177] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_384 (.DIODE(\mprj_logic1[177] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_385 (.DIODE(\mprj_logic1[177] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_386 (.DIODE(\mprj_logic1[177] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_387 (.DIODE(\mprj_logic1[177] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_388 (.DIODE(\mprj_logic1[177] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_389 (.DIODE(\mprj_logic1[177] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_390 (.DIODE(\mprj_logic1[177] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_391 (.DIODE(\mprj_logic1[177] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_392 (.DIODE(\mprj_logic1[177] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_393 (.DIODE(\mprj_logic1[177] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_394 (.DIODE(\mprj_logic1[177] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_395 (.DIODE(\mprj_logic1[177] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_396 (.DIODE(\mprj_logic1[178] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_397 (.DIODE(\mprj_logic1[178] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_398 (.DIODE(\mprj_logic1[178] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_399 (.DIODE(\mprj_logic1[178] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_400 (.DIODE(\mprj_logic1[178] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_401 (.DIODE(\mprj_logic1[178] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_402 (.DIODE(\mprj_logic1[178] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_403 (.DIODE(\mprj_logic1[178] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_404 (.DIODE(\mprj_logic1[178] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_405 (.DIODE(\mprj_logic1[178] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_406 (.DIODE(\mprj_logic1[180] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_407 (.DIODE(\mprj_logic1[182] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_408 (.DIODE(\mprj_logic1[182] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_409 (.DIODE(\mprj_logic1[182] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_410 (.DIODE(\mprj_logic1[182] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_411 (.DIODE(\mprj_logic1[182] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_412 (.DIODE(\mprj_logic1[182] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_413 (.DIODE(\mprj_logic1[182] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_414 (.DIODE(\mprj_logic1[182] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_415 (.DIODE(\mprj_logic1[182] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_416 (.DIODE(\mprj_logic1[182] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_417 (.DIODE(\mprj_logic1[182] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_418 (.DIODE(\mprj_logic1[182] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_419 (.DIODE(\mprj_logic1[182] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_420 (.DIODE(\mprj_logic1[182] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_421 (.DIODE(\mprj_logic1[182] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_422 (.DIODE(\mprj_logic1[182] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_423 (.DIODE(\mprj_logic1[182] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_424 (.DIODE(\mprj_logic1[182] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_425 (.DIODE(\mprj_logic1[182] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_426 (.DIODE(\mprj_logic1[182] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_427 (.DIODE(\mprj_logic1[184] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_428 (.DIODE(\mprj_logic1[184] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_429 (.DIODE(\mprj_logic1[184] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_430 (.DIODE(\mprj_logic1[185] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_431 (.DIODE(\mprj_logic1[187] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_432 (.DIODE(\mprj_logic1[187] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_433 (.DIODE(\mprj_logic1[187] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_434 (.DIODE(\mprj_logic1[188] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_435 (.DIODE(\mprj_logic1[188] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_436 (.DIODE(\mprj_logic1[188] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_437 (.DIODE(\mprj_logic1[188] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_438 (.DIODE(\mprj_logic1[188] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_439 (.DIODE(\mprj_logic1[188] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_440 (.DIODE(\mprj_logic1[188] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_441 (.DIODE(\mprj_logic1[188] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_442 (.DIODE(\mprj_logic1[188] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_443 (.DIODE(\mprj_logic1[188] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_444 (.DIODE(\mprj_logic1[188] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_445 (.DIODE(\mprj_logic1[188] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_446 (.DIODE(\mprj_logic1[188] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_447 (.DIODE(\mprj_logic1[188] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_448 (.DIODE(\mprj_logic1[188] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_449 (.DIODE(\mprj_logic1[188] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_450 (.DIODE(\mprj_logic1[188] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_451 (.DIODE(\mprj_logic1[188] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_452 (.DIODE(\mprj_logic1[188] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_453 (.DIODE(\mprj_logic1[188] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_454 (.DIODE(\mprj_logic1[188] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_455 (.DIODE(\mprj_logic1[188] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_456 (.DIODE(\mprj_logic1[189] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_457 (.DIODE(\mprj_logic1[189] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_458 (.DIODE(\mprj_logic1[189] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_459 (.DIODE(\mprj_logic1[189] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_460 (.DIODE(\mprj_logic1[189] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_461 (.DIODE(\mprj_logic1[189] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_462 (.DIODE(\mprj_logic1[189] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_463 (.DIODE(\mprj_logic1[189] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_464 (.DIODE(\mprj_logic1[189] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_465 (.DIODE(\mprj_logic1[189] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_466 (.DIODE(\mprj_logic1[189] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_467 (.DIODE(\mprj_logic1[189] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_468 (.DIODE(\mprj_logic1[189] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_469 (.DIODE(\mprj_logic1[189] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_470 (.DIODE(\mprj_logic1[189] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_471 (.DIODE(\mprj_logic1[189] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_472 (.DIODE(\mprj_logic1[189] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_473 (.DIODE(\mprj_logic1[189] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_474 (.DIODE(\mprj_logic1[189] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_475 (.DIODE(\mprj_logic1[189] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_476 (.DIODE(\mprj_logic1[191] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_477 (.DIODE(\mprj_logic1[191] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_478 (.DIODE(\mprj_logic1[191] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_479 (.DIODE(\mprj_logic1[192] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_480 (.DIODE(\mprj_logic1[192] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_481 (.DIODE(\mprj_logic1[192] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_482 (.DIODE(\mprj_logic1[192] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_483 (.DIODE(\mprj_logic1[192] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_484 (.DIODE(\mprj_logic1[192] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_485 (.DIODE(\mprj_logic1[192] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_486 (.DIODE(\mprj_logic1[192] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_487 (.DIODE(\mprj_logic1[192] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_488 (.DIODE(\mprj_logic1[192] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_489 (.DIODE(\mprj_logic1[192] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_490 (.DIODE(\mprj_logic1[193] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_491 (.DIODE(\mprj_logic1[193] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_492 (.DIODE(\mprj_logic1[193] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_493 (.DIODE(\mprj_logic1[193] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_494 (.DIODE(\mprj_logic1[193] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_495 (.DIODE(\mprj_logic1[193] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_496 (.DIODE(\mprj_logic1[193] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_497 (.DIODE(\mprj_logic1[193] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_498 (.DIODE(\mprj_logic1[193] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_499 (.DIODE(\mprj_logic1[193] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_500 (.DIODE(\mprj_logic1[193] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_501 (.DIODE(\mprj_logic1[195] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_502 (.DIODE(\mprj_logic1[195] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_503 (.DIODE(\mprj_logic1[195] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_504 (.DIODE(\mprj_logic1[195] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_505 (.DIODE(\mprj_logic1[195] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_506 (.DIODE(\mprj_logic1[195] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_507 (.DIODE(\mprj_logic1[195] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_508 (.DIODE(\mprj_logic1[195] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_509 (.DIODE(\mprj_logic1[195] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_510 (.DIODE(\mprj_logic1[195] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_511 (.DIODE(\mprj_logic1[195] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_512 (.DIODE(\mprj_logic1[196] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_513 (.DIODE(\mprj_logic1[196] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_514 (.DIODE(\mprj_logic1[196] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_515 (.DIODE(\mprj_logic1[196] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_516 (.DIODE(\mprj_logic1[196] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_517 (.DIODE(\mprj_logic1[196] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_518 (.DIODE(\mprj_logic1[196] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_519 (.DIODE(\mprj_logic1[196] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_520 (.DIODE(\mprj_logic1[196] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_521 (.DIODE(\mprj_logic1[196] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_522 (.DIODE(\mprj_logic1[197] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_523 (.DIODE(\mprj_logic1[198] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_524 (.DIODE(\mprj_logic1[198] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_525 (.DIODE(\mprj_logic1[199] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_526 (.DIODE(\mprj_logic1[200] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_527 (.DIODE(\mprj_logic1[200] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_528 (.DIODE(\mprj_logic1[200] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_529 (.DIODE(\mprj_logic1[200] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_530 (.DIODE(\mprj_logic1[200] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_531 (.DIODE(\mprj_logic1[200] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_532 (.DIODE(\mprj_logic1[200] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_533 (.DIODE(\mprj_logic1[200] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_534 (.DIODE(\mprj_logic1[201] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_535 (.DIODE(\mprj_logic1[201] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_536 (.DIODE(\mprj_logic1[201] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_537 (.DIODE(\mprj_logic1[201] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_538 (.DIODE(\mprj_logic1[201] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_539 (.DIODE(\mprj_logic1[201] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_540 (.DIODE(\mprj_logic1[201] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_541 (.DIODE(\mprj_logic1[201] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_542 (.DIODE(\mprj_logic1[202] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_543 (.DIODE(\mprj_logic1[203] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_544 (.DIODE(\mprj_logic1[203] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_545 (.DIODE(\mprj_logic1[203] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_546 (.DIODE(\mprj_logic1[203] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_547 (.DIODE(\mprj_logic1[203] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_548 (.DIODE(\mprj_logic1[203] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_549 (.DIODE(\mprj_logic1[203] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_550 (.DIODE(\mprj_logic1[203] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_551 (.DIODE(\mprj_logic1[203] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_552 (.DIODE(\mprj_logic1[203] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_553 (.DIODE(\mprj_logic1[203] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_554 (.DIODE(\mprj_logic1[203] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_555 (.DIODE(\mprj_logic1[203] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_556 (.DIODE(\mprj_logic1[203] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_557 (.DIODE(\mprj_logic1[203] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_558 (.DIODE(\mprj_logic1[203] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_559 (.DIODE(\mprj_logic1[203] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_560 (.DIODE(\mprj_logic1[203] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_561 (.DIODE(\mprj_logic1[204] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_562 (.DIODE(\mprj_logic1[204] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_563 (.DIODE(\mprj_logic1[204] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_564 (.DIODE(\mprj_logic1[204] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_565 (.DIODE(\mprj_logic1[204] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_566 (.DIODE(\mprj_logic1[204] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_567 (.DIODE(\mprj_logic1[204] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_568 (.DIODE(\mprj_logic1[205] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_569 (.DIODE(\mprj_logic1[206] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_570 (.DIODE(\mprj_logic1[207] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_571 (.DIODE(\mprj_logic1[207] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_572 (.DIODE(\mprj_logic1[207] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_573 (.DIODE(\mprj_logic1[207] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_574 (.DIODE(\mprj_logic1[207] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_575 (.DIODE(\mprj_logic1[207] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_576 (.DIODE(\mprj_logic1[207] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_577 (.DIODE(\mprj_logic1[207] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_578 (.DIODE(\mprj_logic1[207] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_579 (.DIODE(\mprj_logic1[207] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_580 (.DIODE(\mprj_logic1[207] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_581 (.DIODE(\mprj_logic1[207] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_582 (.DIODE(\mprj_logic1[207] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_583 (.DIODE(\mprj_logic1[207] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_584 (.DIODE(\mprj_logic1[207] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_585 (.DIODE(\mprj_logic1[207] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_586 (.DIODE(\mprj_logic1[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_587 (.DIODE(\mprj_logic1[211] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_588 (.DIODE(\mprj_logic1[211] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_589 (.DIODE(\mprj_logic1[211] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_590 (.DIODE(\mprj_logic1[211] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_591 (.DIODE(\mprj_logic1[211] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_592 (.DIODE(\mprj_logic1[212] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_593 (.DIODE(\mprj_logic1[215] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_594 (.DIODE(\mprj_logic1[215] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_595 (.DIODE(\mprj_logic1[215] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_596 (.DIODE(\mprj_logic1[215] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_597 (.DIODE(\mprj_logic1[215] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_598 (.DIODE(\mprj_logic1[215] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_599 (.DIODE(\mprj_logic1[215] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_600 (.DIODE(\mprj_logic1[215] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_601 (.DIODE(\mprj_logic1[215] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_602 (.DIODE(\mprj_logic1[215] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_603 (.DIODE(\mprj_logic1[216] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_604 (.DIODE(\mprj_logic1[216] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_605 (.DIODE(\mprj_logic1[216] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_606 (.DIODE(\mprj_logic1[216] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_607 (.DIODE(\mprj_logic1[216] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_608 (.DIODE(\mprj_logic1[216] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_609 (.DIODE(\mprj_logic1[216] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_610 (.DIODE(\mprj_logic1[216] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_611 (.DIODE(\mprj_logic1[216] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_612 (.DIODE(\mprj_logic1[216] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_613 (.DIODE(\mprj_logic1[216] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_614 (.DIODE(\mprj_logic1[216] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_615 (.DIODE(\mprj_logic1[218] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_616 (.DIODE(\mprj_logic1[219] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_617 (.DIODE(\mprj_logic1[221] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_618 (.DIODE(\mprj_logic1[221] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_619 (.DIODE(\mprj_logic1[222] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_620 (.DIODE(\mprj_logic1[222] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_621 (.DIODE(\mprj_logic1[223] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_622 (.DIODE(\mprj_logic1[224] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_623 (.DIODE(\mprj_logic1[224] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_624 (.DIODE(\mprj_logic1[225] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_625 (.DIODE(\mprj_logic1[226] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_626 (.DIODE(\mprj_logic1[226] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_627 (.DIODE(\mprj_logic1[229] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_628 (.DIODE(\mprj_logic1[240] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_629 (.DIODE(\mprj_logic1[246] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_630 (.DIODE(\mprj_logic1[254] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_631 (.DIODE(\mprj_logic1[257] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_632 (.DIODE(\mprj_logic1[257] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_633 (.DIODE(\mprj_logic1[262] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_634 (.DIODE(\mprj_logic1[263] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_635 (.DIODE(\mprj_logic1[264] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_636 (.DIODE(\mprj_logic1[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_637 (.DIODE(\mprj_logic1[270] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_638 (.DIODE(\mprj_logic1[270] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_639 (.DIODE(\mprj_logic1[270] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_640 (.DIODE(\mprj_logic1[271] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_641 (.DIODE(\mprj_logic1[271] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_642 (.DIODE(\mprj_logic1[271] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_643 (.DIODE(\mprj_logic1[272] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_644 (.DIODE(\mprj_logic1[272] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_645 (.DIODE(\mprj_logic1[272] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_646 (.DIODE(\mprj_logic1[273] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_647 (.DIODE(\mprj_logic1[273] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_648 (.DIODE(\mprj_logic1[273] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_649 (.DIODE(\mprj_logic1[273] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_650 (.DIODE(\mprj_logic1[273] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_651 (.DIODE(\mprj_logic1[273] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_652 (.DIODE(\mprj_logic1[273] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_653 (.DIODE(\mprj_logic1[273] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_654 (.DIODE(\mprj_logic1[273] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_655 (.DIODE(\mprj_logic1[273] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_656 (.DIODE(\mprj_logic1[273] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_657 (.DIODE(\mprj_logic1[274] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_658 (.DIODE(\mprj_logic1[274] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_659 (.DIODE(\mprj_logic1[274] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_660 (.DIODE(\mprj_logic1[274] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_661 (.DIODE(\mprj_logic1[274] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_662 (.DIODE(\mprj_logic1[274] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_663 (.DIODE(\mprj_logic1[275] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_664 (.DIODE(\mprj_logic1[276] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_665 (.DIODE(\mprj_logic1[279] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_666 (.DIODE(\mprj_logic1[279] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_667 (.DIODE(\mprj_logic1[279] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_668 (.DIODE(\mprj_logic1[279] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_669 (.DIODE(\mprj_logic1[279] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_670 (.DIODE(\mprj_logic1[279] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_671 (.DIODE(\mprj_logic1[279] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_672 (.DIODE(\mprj_logic1[279] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_673 (.DIODE(\mprj_logic1[279] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_674 (.DIODE(\mprj_logic1[279] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_675 (.DIODE(\mprj_logic1[281] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_676 (.DIODE(\mprj_logic1[281] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_677 (.DIODE(\mprj_logic1[281] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_678 (.DIODE(\mprj_logic1[281] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_679 (.DIODE(\mprj_logic1[281] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_680 (.DIODE(\mprj_logic1[281] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_681 (.DIODE(\mprj_logic1[281] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_682 (.DIODE(\mprj_logic1[281] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_683 (.DIODE(\mprj_logic1[281] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_684 (.DIODE(\mprj_logic1[282] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_685 (.DIODE(\mprj_logic1[283] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_686 (.DIODE(\mprj_logic1[284] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_687 (.DIODE(\mprj_logic1[284] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_688 (.DIODE(\mprj_logic1[284] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_689 (.DIODE(\mprj_logic1[285] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_690 (.DIODE(\mprj_logic1[286] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_691 (.DIODE(\mprj_logic1[287] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_692 (.DIODE(\mprj_logic1[287] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_693 (.DIODE(\mprj_logic1[287] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_694 (.DIODE(\mprj_logic1[287] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_695 (.DIODE(\mprj_logic1[287] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_696 (.DIODE(\mprj_logic1[287] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_697 (.DIODE(\mprj_logic1[287] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_698 (.DIODE(\mprj_logic1[288] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_699 (.DIODE(\mprj_logic1[288] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_700 (.DIODE(\mprj_logic1[288] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_701 (.DIODE(\mprj_logic1[288] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_702 (.DIODE(\mprj_logic1[288] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_703 (.DIODE(\mprj_logic1[288] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_704 (.DIODE(\mprj_logic1[288] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_705 (.DIODE(\mprj_logic1[288] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_706 (.DIODE(\mprj_logic1[288] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_707 (.DIODE(\mprj_logic1[289] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_708 (.DIODE(\mprj_logic1[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_709 (.DIODE(\mprj_logic1[290] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_710 (.DIODE(\mprj_logic1[293] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_711 (.DIODE(\mprj_logic1[296] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_712 (.DIODE(\mprj_logic1[298] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_713 (.DIODE(\mprj_logic1[299] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_714 (.DIODE(\mprj_logic1[299] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_715 (.DIODE(\mprj_logic1[299] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_716 (.DIODE(\mprj_logic1[299] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_717 (.DIODE(\mprj_logic1[299] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_718 (.DIODE(\mprj_logic1[299] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_719 (.DIODE(\mprj_logic1[299] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_720 (.DIODE(\mprj_logic1[299] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_721 (.DIODE(\mprj_logic1[299] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_722 (.DIODE(\mprj_logic1[299] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_723 (.DIODE(\mprj_logic1[299] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_724 (.DIODE(\mprj_logic1[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_725 (.DIODE(\mprj_logic1[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_726 (.DIODE(\mprj_logic1[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_727 (.DIODE(\mprj_logic1[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_728 (.DIODE(\mprj_logic1[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_729 (.DIODE(\mprj_logic1[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_730 (.DIODE(\mprj_logic1[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_731 (.DIODE(\mprj_logic1[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_732 (.DIODE(\mprj_logic1[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_733 (.DIODE(\mprj_logic1[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_734 (.DIODE(\mprj_logic1[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_735 (.DIODE(\mprj_logic1[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_736 (.DIODE(\mprj_logic1[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_737 (.DIODE(\mprj_logic1[300] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_738 (.DIODE(\mprj_logic1[300] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_739 (.DIODE(\mprj_logic1[300] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_740 (.DIODE(\mprj_logic1[300] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_741 (.DIODE(\mprj_logic1[300] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_742 (.DIODE(\mprj_logic1[300] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_743 (.DIODE(\mprj_logic1[300] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_744 (.DIODE(\mprj_logic1[300] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_745 (.DIODE(\mprj_logic1[300] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_746 (.DIODE(\mprj_logic1[300] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_747 (.DIODE(\mprj_logic1[300] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_748 (.DIODE(\mprj_logic1[301] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_749 (.DIODE(\mprj_logic1[302] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_750 (.DIODE(\mprj_logic1[302] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_751 (.DIODE(\mprj_logic1[302] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_752 (.DIODE(\mprj_logic1[302] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_753 (.DIODE(\mprj_logic1[302] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_754 (.DIODE(\mprj_logic1[302] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_755 (.DIODE(\mprj_logic1[302] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_756 (.DIODE(\mprj_logic1[302] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_757 (.DIODE(\mprj_logic1[302] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_758 (.DIODE(\mprj_logic1[302] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_759 (.DIODE(\mprj_logic1[302] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_760 (.DIODE(\mprj_logic1[302] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_761 (.DIODE(\mprj_logic1[303] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_762 (.DIODE(\mprj_logic1[303] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_763 (.DIODE(\mprj_logic1[303] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_764 (.DIODE(\mprj_logic1[303] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_765 (.DIODE(\mprj_logic1[303] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_766 (.DIODE(\mprj_logic1[303] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_767 (.DIODE(\mprj_logic1[303] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_768 (.DIODE(\mprj_logic1[303] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_769 (.DIODE(\mprj_logic1[303] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_770 (.DIODE(\mprj_logic1[304] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_771 (.DIODE(\mprj_logic1[305] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_772 (.DIODE(\mprj_logic1[306] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_773 (.DIODE(\mprj_logic1[308] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_774 (.DIODE(\mprj_logic1[308] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_775 (.DIODE(\mprj_logic1[308] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_776 (.DIODE(\mprj_logic1[308] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_777 (.DIODE(\mprj_logic1[308] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_778 (.DIODE(\mprj_logic1[308] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_779 (.DIODE(\mprj_logic1[308] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_780 (.DIODE(\mprj_logic1[308] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_781 (.DIODE(\mprj_logic1[309] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_782 (.DIODE(\mprj_logic1[309] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_783 (.DIODE(\mprj_logic1[309] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_784 (.DIODE(\mprj_logic1[309] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_785 (.DIODE(\mprj_logic1[309] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_786 (.DIODE(\mprj_logic1[309] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_787 (.DIODE(\mprj_logic1[309] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_788 (.DIODE(\mprj_logic1[309] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_789 (.DIODE(\mprj_logic1[309] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_790 (.DIODE(\mprj_logic1[309] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_791 (.DIODE(\mprj_logic1[309] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_792 (.DIODE(\mprj_logic1[309] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_793 (.DIODE(\mprj_logic1[309] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_794 (.DIODE(\mprj_logic1[310] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_795 (.DIODE(\mprj_logic1[310] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_796 (.DIODE(\mprj_logic1[310] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_797 (.DIODE(\mprj_logic1[310] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_798 (.DIODE(\mprj_logic1[310] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_799 (.DIODE(\mprj_logic1[310] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_800 (.DIODE(\mprj_logic1[310] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_801 (.DIODE(\mprj_logic1[310] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_802 (.DIODE(\mprj_logic1[310] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_803 (.DIODE(\mprj_logic1[310] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_804 (.DIODE(\mprj_logic1[310] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_805 (.DIODE(\mprj_logic1[310] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_806 (.DIODE(\mprj_logic1[310] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_807 (.DIODE(\mprj_logic1[311] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_808 (.DIODE(\mprj_logic1[312] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_809 (.DIODE(\mprj_logic1[313] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_810 (.DIODE(\mprj_logic1[313] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_811 (.DIODE(\mprj_logic1[314] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_812 (.DIODE(\mprj_logic1[314] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_813 (.DIODE(\mprj_logic1[316] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_814 (.DIODE(\mprj_logic1[316] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_815 (.DIODE(\mprj_logic1[316] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_816 (.DIODE(\mprj_logic1[316] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_817 (.DIODE(\mprj_logic1[316] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_818 (.DIODE(\mprj_logic1[316] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_819 (.DIODE(\mprj_logic1[316] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_820 (.DIODE(\mprj_logic1[316] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_821 (.DIODE(\mprj_logic1[316] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_822 (.DIODE(\mprj_logic1[316] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_823 (.DIODE(\mprj_logic1[316] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_824 (.DIODE(\mprj_logic1[316] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_825 (.DIODE(\mprj_logic1[316] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_826 (.DIODE(\mprj_logic1[317] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_827 (.DIODE(\mprj_logic1[317] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_828 (.DIODE(\mprj_logic1[317] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_829 (.DIODE(\mprj_logic1[317] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_830 (.DIODE(\mprj_logic1[317] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_831 (.DIODE(\mprj_logic1[317] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_832 (.DIODE(\mprj_logic1[317] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_833 (.DIODE(\mprj_logic1[317] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_834 (.DIODE(\mprj_logic1[317] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_835 (.DIODE(\mprj_logic1[317] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_836 (.DIODE(\mprj_logic1[317] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_837 (.DIODE(\mprj_logic1[317] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_838 (.DIODE(\mprj_logic1[317] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_839 (.DIODE(\mprj_logic1[317] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_840 (.DIODE(\mprj_logic1[317] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_841 (.DIODE(\mprj_logic1[317] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_842 (.DIODE(\mprj_logic1[317] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_843 (.DIODE(\mprj_logic1[317] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_844 (.DIODE(\mprj_logic1[317] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_845 (.DIODE(\mprj_logic1[317] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_846 (.DIODE(\mprj_logic1[317] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_847 (.DIODE(\mprj_logic1[317] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_848 (.DIODE(\mprj_logic1[318] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_849 (.DIODE(\mprj_logic1[318] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_850 (.DIODE(\mprj_logic1[318] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_851 (.DIODE(\mprj_logic1[319] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_852 (.DIODE(\mprj_logic1[319] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_853 (.DIODE(\mprj_logic1[319] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_854 (.DIODE(\mprj_logic1[319] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_855 (.DIODE(\mprj_logic1[319] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_856 (.DIODE(\mprj_logic1[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_857 (.DIODE(\mprj_logic1[320] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_858 (.DIODE(\mprj_logic1[322] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_859 (.DIODE(\mprj_logic1[322] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_860 (.DIODE(\mprj_logic1[322] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_861 (.DIODE(\mprj_logic1[322] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_862 (.DIODE(\mprj_logic1[322] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_863 (.DIODE(\mprj_logic1[322] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_864 (.DIODE(\mprj_logic1[322] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_865 (.DIODE(\mprj_logic1[322] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_866 (.DIODE(\mprj_logic1[322] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_867 (.DIODE(\mprj_logic1[322] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_868 (.DIODE(\mprj_logic1[322] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_869 (.DIODE(\mprj_logic1[322] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_870 (.DIODE(\mprj_logic1[322] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_871 (.DIODE(\mprj_logic1[322] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_872 (.DIODE(\mprj_logic1[322] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_873 (.DIODE(\mprj_logic1[322] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_874 (.DIODE(\mprj_logic1[322] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_875 (.DIODE(\mprj_logic1[322] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_876 (.DIODE(\mprj_logic1[322] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_877 (.DIODE(\mprj_logic1[322] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_878 (.DIODE(\mprj_logic1[322] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_879 (.DIODE(\mprj_logic1[322] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_880 (.DIODE(\mprj_logic1[323] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_881 (.DIODE(\mprj_logic1[323] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_882 (.DIODE(\mprj_logic1[323] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_883 (.DIODE(\mprj_logic1[323] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_884 (.DIODE(\mprj_logic1[323] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_885 (.DIODE(\mprj_logic1[323] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_886 (.DIODE(\mprj_logic1[323] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_887 (.DIODE(\mprj_logic1[323] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_888 (.DIODE(\mprj_logic1[323] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_889 (.DIODE(\mprj_logic1[323] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_890 (.DIODE(\mprj_logic1[323] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_891 (.DIODE(\mprj_logic1[323] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_892 (.DIODE(\mprj_logic1[323] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_893 (.DIODE(\mprj_logic1[323] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_894 (.DIODE(\mprj_logic1[323] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_895 (.DIODE(\mprj_logic1[323] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_896 (.DIODE(\mprj_logic1[323] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_897 (.DIODE(\mprj_logic1[323] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_898 (.DIODE(\mprj_logic1[323] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_899 (.DIODE(\mprj_logic1[323] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_900 (.DIODE(\mprj_logic1[323] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_901 (.DIODE(\mprj_logic1[323] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_902 (.DIODE(\mprj_logic1[324] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_903 (.DIODE(\mprj_logic1[324] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_904 (.DIODE(\mprj_logic1[324] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_905 (.DIODE(\mprj_logic1[324] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_906 (.DIODE(\mprj_logic1[324] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_907 (.DIODE(\mprj_logic1[324] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_908 (.DIODE(\mprj_logic1[324] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_909 (.DIODE(\mprj_logic1[324] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_910 (.DIODE(\mprj_logic1[324] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_911 (.DIODE(\mprj_logic1[324] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_912 (.DIODE(\mprj_logic1[324] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_913 (.DIODE(\mprj_logic1[324] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_914 (.DIODE(\mprj_logic1[324] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_915 (.DIODE(\mprj_logic1[324] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_916 (.DIODE(\mprj_logic1[324] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_917 (.DIODE(\mprj_logic1[324] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_918 (.DIODE(\mprj_logic1[324] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_919 (.DIODE(\mprj_logic1[324] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_920 (.DIODE(\mprj_logic1[324] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_921 (.DIODE(\mprj_logic1[324] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_922 (.DIODE(\mprj_logic1[325] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_923 (.DIODE(\mprj_logic1[325] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_924 (.DIODE(\mprj_logic1[325] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_925 (.DIODE(\mprj_logic1[325] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_926 (.DIODE(\mprj_logic1[325] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_927 (.DIODE(\mprj_logic1[325] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_928 (.DIODE(\mprj_logic1[325] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_929 (.DIODE(\mprj_logic1[325] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_930 (.DIODE(\mprj_logic1[325] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_931 (.DIODE(\mprj_logic1[325] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_932 (.DIODE(\mprj_logic1[325] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_933 (.DIODE(\mprj_logic1[325] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_934 (.DIODE(\mprj_logic1[325] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_935 (.DIODE(\mprj_logic1[326] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_936 (.DIODE(\mprj_logic1[326] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_937 (.DIODE(\mprj_logic1[326] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_938 (.DIODE(\mprj_logic1[326] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_939 (.DIODE(\mprj_logic1[326] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_940 (.DIODE(\mprj_logic1[326] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_941 (.DIODE(\mprj_logic1[326] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_942 (.DIODE(\mprj_logic1[326] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_943 (.DIODE(\mprj_logic1[326] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_944 (.DIODE(\mprj_logic1[326] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_945 (.DIODE(\mprj_logic1[326] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_946 (.DIODE(\mprj_logic1[327] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_947 (.DIODE(\mprj_logic1[327] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_948 (.DIODE(\mprj_logic1[327] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_949 (.DIODE(\mprj_logic1[327] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_950 (.DIODE(\mprj_logic1[327] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_951 (.DIODE(\mprj_logic1[327] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_952 (.DIODE(\mprj_logic1[327] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_953 (.DIODE(\mprj_logic1[327] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_954 (.DIODE(\mprj_logic1[327] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_955 (.DIODE(\mprj_logic1[327] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_956 (.DIODE(\mprj_logic1[327] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_957 (.DIODE(\mprj_logic1[327] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_958 (.DIODE(\mprj_logic1[327] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_959 (.DIODE(\mprj_logic1[327] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_960 (.DIODE(\mprj_logic1[327] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_961 (.DIODE(\mprj_logic1[327] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_962 (.DIODE(\mprj_logic1[327] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_963 (.DIODE(\mprj_logic1[327] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_964 (.DIODE(\mprj_logic1[327] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_965 (.DIODE(\mprj_logic1[327] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_966 (.DIODE(\mprj_logic1[327] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_967 (.DIODE(\mprj_logic1[327] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_968 (.DIODE(\mprj_logic1[328] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_969 (.DIODE(\mprj_logic1[328] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_970 (.DIODE(\mprj_logic1[328] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_971 (.DIODE(\mprj_logic1[328] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_972 (.DIODE(\mprj_logic1[328] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_973 (.DIODE(\mprj_logic1[328] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_974 (.DIODE(\mprj_logic1[328] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_975 (.DIODE(\mprj_logic1[328] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_976 (.DIODE(\mprj_logic1[328] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_977 (.DIODE(\mprj_logic1[328] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_978 (.DIODE(\mprj_logic1[328] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_979 (.DIODE(\mprj_logic1[328] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_980 (.DIODE(\mprj_logic1[328] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_981 (.DIODE(\mprj_logic1[329] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_982 (.DIODE(\mprj_logic1[329] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_983 (.DIODE(\mprj_logic1[329] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_984 (.DIODE(\mprj_logic1[329] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_985 (.DIODE(\mprj_logic1[329] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_986 (.DIODE(\mprj_logic1[329] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_987 (.DIODE(\mprj_logic1[329] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_988 (.DIODE(\mprj_logic1[329] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_989 (.DIODE(\mprj_logic1[329] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_990 (.DIODE(\mprj_logic1[329] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_991 (.DIODE(\mprj_logic1[329] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_992 (.DIODE(\mprj_logic1[329] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_993 (.DIODE(\mprj_logic1[329] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_994 (.DIODE(\mprj_logic1[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_995 (.DIODE(\mprj_logic1[330] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_996 (.DIODE(\mprj_logic1[330] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_997 (.DIODE(\mprj_logic1[330] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_998 (.DIODE(\mprj_logic1[330] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_999 (.DIODE(\mprj_logic1[330] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1000 (.DIODE(\mprj_logic1[330] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1001 (.DIODE(\mprj_logic1[330] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1002 (.DIODE(\mprj_logic1[330] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1003 (.DIODE(\mprj_logic1[330] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1004 (.DIODE(\mprj_logic1[330] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1005 (.DIODE(\mprj_logic1[330] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1006 (.DIODE(\mprj_logic1[330] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1007 (.DIODE(\mprj_logic1[330] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1008 (.DIODE(\mprj_logic1[330] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1009 (.DIODE(\mprj_logic1[330] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1010 (.DIODE(\mprj_logic1[330] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1011 (.DIODE(\mprj_logic1[330] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1012 (.DIODE(\mprj_logic1[330] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1013 (.DIODE(\mprj_logic1[330] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1014 (.DIODE(\mprj_logic1[330] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1015 (.DIODE(\mprj_logic1[330] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1016 (.DIODE(\mprj_logic1[330] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1017 (.DIODE(\mprj_logic1[331] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1018 (.DIODE(\mprj_logic1[331] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1019 (.DIODE(\mprj_logic1[331] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1020 (.DIODE(\mprj_logic1[331] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1021 (.DIODE(\mprj_logic1[331] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1022 (.DIODE(\mprj_logic1[331] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1023 (.DIODE(\mprj_logic1[331] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1024 (.DIODE(\mprj_logic1[331] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1025 (.DIODE(\mprj_logic1[331] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1026 (.DIODE(\mprj_logic1[331] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1027 (.DIODE(\mprj_logic1[331] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1028 (.DIODE(\mprj_logic1[331] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1029 (.DIODE(\mprj_logic1[331] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1030 (.DIODE(\mprj_logic1[331] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1031 (.DIODE(\mprj_logic1[331] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1032 (.DIODE(\mprj_logic1[331] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1033 (.DIODE(\mprj_logic1[331] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1034 (.DIODE(\mprj_logic1[331] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1035 (.DIODE(\mprj_logic1[331] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1036 (.DIODE(\mprj_logic1[331] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1037 (.DIODE(\mprj_logic1[331] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1038 (.DIODE(\mprj_logic1[331] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1039 (.DIODE(\mprj_logic1[332] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1040 (.DIODE(\mprj_logic1[332] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1041 (.DIODE(\mprj_logic1[332] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1042 (.DIODE(\mprj_logic1[333] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1043 (.DIODE(\mprj_logic1[333] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1044 (.DIODE(\mprj_logic1[333] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1045 (.DIODE(\mprj_logic1[333] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1046 (.DIODE(\mprj_logic1[334] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1047 (.DIODE(\mprj_logic1[334] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1048 (.DIODE(\mprj_logic1[334] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1049 (.DIODE(\mprj_logic1[334] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1050 (.DIODE(\mprj_logic1[334] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1051 (.DIODE(\mprj_logic1[335] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1052 (.DIODE(\mprj_logic1[336] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1053 (.DIODE(\mprj_logic1[337] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1054 (.DIODE(\mprj_logic1[339] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1055 (.DIODE(\mprj_logic1[340] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1056 (.DIODE(\mprj_logic1[341] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1057 (.DIODE(\mprj_logic1[342] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1058 (.DIODE(\mprj_logic1[343] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1059 (.DIODE(\mprj_logic1[343] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1060 (.DIODE(\mprj_logic1[343] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1061 (.DIODE(\mprj_logic1[343] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1062 (.DIODE(\mprj_logic1[343] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1063 (.DIODE(\mprj_logic1[344] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1064 (.DIODE(\mprj_logic1[345] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1065 (.DIODE(\mprj_logic1[346] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1066 (.DIODE(\mprj_logic1[347] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1067 (.DIODE(\mprj_logic1[348] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1068 (.DIODE(\mprj_logic1[349] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1069 (.DIODE(\mprj_logic1[349] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1070 (.DIODE(\mprj_logic1[349] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1071 (.DIODE(\mprj_logic1[349] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1072 (.DIODE(\mprj_logic1[349] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1073 (.DIODE(\mprj_logic1[349] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1074 (.DIODE(\mprj_logic1[349] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1075 (.DIODE(\mprj_logic1[349] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1076 (.DIODE(\mprj_logic1[349] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1077 (.DIODE(\mprj_logic1[349] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1078 (.DIODE(\mprj_logic1[349] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1079 (.DIODE(\mprj_logic1[34] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1080 (.DIODE(\mprj_logic1[350] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1081 (.DIODE(\mprj_logic1[350] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1082 (.DIODE(\mprj_logic1[350] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1083 (.DIODE(\mprj_logic1[350] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1084 (.DIODE(\mprj_logic1[350] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1085 (.DIODE(\mprj_logic1[350] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1086 (.DIODE(\mprj_logic1[350] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1087 (.DIODE(\mprj_logic1[350] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1088 (.DIODE(\mprj_logic1[350] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1089 (.DIODE(\mprj_logic1[350] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1090 (.DIODE(\mprj_logic1[350] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1091 (.DIODE(\mprj_logic1[350] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1092 (.DIODE(\mprj_logic1[350] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1093 (.DIODE(\mprj_logic1[350] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1094 (.DIODE(\mprj_logic1[350] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1095 (.DIODE(\mprj_logic1[350] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1096 (.DIODE(\mprj_logic1[350] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1097 (.DIODE(\mprj_logic1[350] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1098 (.DIODE(\mprj_logic1[350] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1099 (.DIODE(\mprj_logic1[350] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1100 (.DIODE(\mprj_logic1[350] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1101 (.DIODE(\mprj_logic1[350] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1102 (.DIODE(\mprj_logic1[351] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1103 (.DIODE(\mprj_logic1[351] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1104 (.DIODE(\mprj_logic1[351] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1105 (.DIODE(\mprj_logic1[351] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1106 (.DIODE(\mprj_logic1[351] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1107 (.DIODE(\mprj_logic1[351] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1108 (.DIODE(\mprj_logic1[351] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1109 (.DIODE(\mprj_logic1[351] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1110 (.DIODE(\mprj_logic1[351] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1111 (.DIODE(\mprj_logic1[351] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1112 (.DIODE(\mprj_logic1[351] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1113 (.DIODE(\mprj_logic1[351] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1114 (.DIODE(\mprj_logic1[351] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1115 (.DIODE(\mprj_logic1[351] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1116 (.DIODE(\mprj_logic1[351] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1117 (.DIODE(\mprj_logic1[351] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1118 (.DIODE(\mprj_logic1[351] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1119 (.DIODE(\mprj_logic1[351] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1120 (.DIODE(\mprj_logic1[351] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1121 (.DIODE(\mprj_logic1[351] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1122 (.DIODE(\mprj_logic1[351] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1123 (.DIODE(\mprj_logic1[351] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1124 (.DIODE(\mprj_logic1[352] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1125 (.DIODE(\mprj_logic1[352] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1126 (.DIODE(\mprj_logic1[352] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1127 (.DIODE(\mprj_logic1[352] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1128 (.DIODE(\mprj_logic1[353] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1129 (.DIODE(\mprj_logic1[353] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1130 (.DIODE(\mprj_logic1[353] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1131 (.DIODE(\mprj_logic1[355] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1132 (.DIODE(\mprj_logic1[356] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1133 (.DIODE(\mprj_logic1[357] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1134 (.DIODE(\mprj_logic1[357] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1135 (.DIODE(\mprj_logic1[358] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1136 (.DIODE(\mprj_logic1[358] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1137 (.DIODE(\mprj_logic1[359] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1138 (.DIODE(\mprj_logic1[361] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1139 (.DIODE(\mprj_logic1[361] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1140 (.DIODE(\mprj_logic1[362] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1141 (.DIODE(\mprj_logic1[362] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1142 (.DIODE(\mprj_logic1[362] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1143 (.DIODE(\mprj_logic1[362] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1144 (.DIODE(\mprj_logic1[363] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1145 (.DIODE(\mprj_logic1[363] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1146 (.DIODE(\mprj_logic1[363] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1147 (.DIODE(\mprj_logic1[363] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1148 (.DIODE(\mprj_logic1[363] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1149 (.DIODE(\mprj_logic1[363] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1150 (.DIODE(\mprj_logic1[364] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1151 (.DIODE(\mprj_logic1[364] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1152 (.DIODE(\mprj_logic1[364] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1153 (.DIODE(\mprj_logic1[364] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1154 (.DIODE(\mprj_logic1[365] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1155 (.DIODE(\mprj_logic1[365] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1156 (.DIODE(\mprj_logic1[365] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1157 (.DIODE(\mprj_logic1[365] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1158 (.DIODE(\mprj_logic1[366] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1159 (.DIODE(\mprj_logic1[366] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1160 (.DIODE(\mprj_logic1[366] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1161 (.DIODE(\mprj_logic1[367] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1162 (.DIODE(\mprj_logic1[368] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1163 (.DIODE(\mprj_logic1[368] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1164 (.DIODE(\mprj_logic1[36] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1165 (.DIODE(\mprj_logic1[372] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1166 (.DIODE(\mprj_logic1[373] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1167 (.DIODE(\mprj_logic1[374] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1168 (.DIODE(\mprj_logic1[376] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1169 (.DIODE(\mprj_logic1[377] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1170 (.DIODE(\mprj_logic1[378] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1171 (.DIODE(\mprj_logic1[379] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1172 (.DIODE(\mprj_logic1[37] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1173 (.DIODE(\mprj_logic1[380] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1174 (.DIODE(\mprj_logic1[381] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1175 (.DIODE(\mprj_logic1[381] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1176 (.DIODE(\mprj_logic1[381] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1177 (.DIODE(\mprj_logic1[382] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1178 (.DIODE(\mprj_logic1[382] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1179 (.DIODE(\mprj_logic1[382] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1180 (.DIODE(\mprj_logic1[383] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1181 (.DIODE(\mprj_logic1[384] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1182 (.DIODE(\mprj_logic1[384] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1183 (.DIODE(\mprj_logic1[386] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1184 (.DIODE(\mprj_logic1[386] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1185 (.DIODE(\mprj_logic1[387] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1186 (.DIODE(\mprj_logic1[387] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1187 (.DIODE(\mprj_logic1[388] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1188 (.DIODE(\mprj_logic1[388] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1189 (.DIODE(\mprj_logic1[38] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1190 (.DIODE(\mprj_logic1[390] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1191 (.DIODE(\mprj_logic1[393] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1192 (.DIODE(\mprj_logic1[393] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1193 (.DIODE(\mprj_logic1[394] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1194 (.DIODE(\mprj_logic1[394] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1195 (.DIODE(\mprj_logic1[395] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1196 (.DIODE(\mprj_logic1[395] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1197 (.DIODE(\mprj_logic1[396] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1198 (.DIODE(\mprj_logic1[396] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1199 (.DIODE(\mprj_logic1[398] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1200 (.DIODE(\mprj_logic1[400] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1201 (.DIODE(\mprj_logic1[400] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1202 (.DIODE(\mprj_logic1[401] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1203 (.DIODE(\mprj_logic1[403] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1204 (.DIODE(\mprj_logic1[406] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1205 (.DIODE(\mprj_logic1[407] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1206 (.DIODE(\mprj_logic1[409] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1207 (.DIODE(\mprj_logic1[411] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1208 (.DIODE(\mprj_logic1[411] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1209 (.DIODE(\mprj_logic1[412] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1210 (.DIODE(\mprj_logic1[413] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1211 (.DIODE(\mprj_logic1[414] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1212 (.DIODE(\mprj_logic1[415] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1213 (.DIODE(\mprj_logic1[416] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1214 (.DIODE(\mprj_logic1[417] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1215 (.DIODE(\mprj_logic1[418] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1216 (.DIODE(\mprj_logic1[419] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1217 (.DIODE(\mprj_logic1[41] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1218 (.DIODE(\mprj_logic1[420] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1219 (.DIODE(\mprj_logic1[421] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1220 (.DIODE(\mprj_logic1[423] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1221 (.DIODE(\mprj_logic1[426] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1222 (.DIODE(\mprj_logic1[427] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1223 (.DIODE(\mprj_logic1[428] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1224 (.DIODE(\mprj_logic1[428] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1225 (.DIODE(\mprj_logic1[429] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1226 (.DIODE(\mprj_logic1[429] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1227 (.DIODE(\mprj_logic1[429] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1228 (.DIODE(\mprj_logic1[429] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1229 (.DIODE(\mprj_logic1[429] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1230 (.DIODE(\mprj_logic1[429] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1231 (.DIODE(\mprj_logic1[429] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1232 (.DIODE(\mprj_logic1[429] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1233 (.DIODE(\mprj_logic1[42] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1234 (.DIODE(\mprj_logic1[433] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1235 (.DIODE(\mprj_logic1[433] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1236 (.DIODE(\mprj_logic1[435] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1237 (.DIODE(\mprj_logic1[436] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1238 (.DIODE(\mprj_logic1[436] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1239 (.DIODE(\mprj_logic1[436] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1240 (.DIODE(\mprj_logic1[436] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1241 (.DIODE(\mprj_logic1[436] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1242 (.DIODE(\mprj_logic1[436] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1243 (.DIODE(\mprj_logic1[436] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1244 (.DIODE(\mprj_logic1[436] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1245 (.DIODE(\mprj_logic1[436] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1246 (.DIODE(\mprj_logic1[436] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1247 (.DIODE(\mprj_logic1[437] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1248 (.DIODE(\mprj_logic1[437] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1249 (.DIODE(\mprj_logic1[438] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1250 (.DIODE(\mprj_logic1[439] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1251 (.DIODE(\mprj_logic1[439] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1252 (.DIODE(\mprj_logic1[439] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1253 (.DIODE(\mprj_logic1[439] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1254 (.DIODE(\mprj_logic1[439] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1255 (.DIODE(\mprj_logic1[439] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1256 (.DIODE(\mprj_logic1[439] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1257 (.DIODE(\mprj_logic1[439] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1258 (.DIODE(\mprj_logic1[439] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1259 (.DIODE(\mprj_logic1[439] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1260 (.DIODE(\mprj_logic1[440] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1261 (.DIODE(\mprj_logic1[440] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1262 (.DIODE(\mprj_logic1[441] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1263 (.DIODE(\mprj_logic1[441] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1264 (.DIODE(\mprj_logic1[441] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1265 (.DIODE(\mprj_logic1[441] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1266 (.DIODE(\mprj_logic1[441] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1267 (.DIODE(\mprj_logic1[441] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1268 (.DIODE(\mprj_logic1[441] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1269 (.DIODE(\mprj_logic1[441] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1270 (.DIODE(\mprj_logic1[442] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1271 (.DIODE(\mprj_logic1[442] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1272 (.DIODE(\mprj_logic1[442] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1273 (.DIODE(\mprj_logic1[442] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1274 (.DIODE(\mprj_logic1[442] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1275 (.DIODE(\mprj_logic1[442] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1276 (.DIODE(\mprj_logic1[442] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1277 (.DIODE(\mprj_logic1[442] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1278 (.DIODE(\mprj_logic1[442] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1279 (.DIODE(\mprj_logic1[442] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1280 (.DIODE(\mprj_logic1[443] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1281 (.DIODE(\mprj_logic1[443] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1282 (.DIODE(\mprj_logic1[443] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1283 (.DIODE(\mprj_logic1[443] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1284 (.DIODE(\mprj_logic1[443] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1285 (.DIODE(\mprj_logic1[443] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1286 (.DIODE(\mprj_logic1[443] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1287 (.DIODE(\mprj_logic1[443] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1288 (.DIODE(\mprj_logic1[445] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1289 (.DIODE(\mprj_logic1[445] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1290 (.DIODE(\mprj_logic1[446] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1291 (.DIODE(\mprj_logic1[446] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1292 (.DIODE(\mprj_logic1[446] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1293 (.DIODE(\mprj_logic1[446] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1294 (.DIODE(\mprj_logic1[446] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1295 (.DIODE(\mprj_logic1[446] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1296 (.DIODE(\mprj_logic1[446] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1297 (.DIODE(\mprj_logic1[446] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1298 (.DIODE(\mprj_logic1[446] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1299 (.DIODE(\mprj_logic1[446] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1300 (.DIODE(\mprj_logic1[447] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1301 (.DIODE(\mprj_logic1[447] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1302 (.DIODE(\mprj_logic1[449] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1303 (.DIODE(\mprj_logic1[449] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1304 (.DIODE(\mprj_logic1[449] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1305 (.DIODE(\mprj_logic1[449] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1306 (.DIODE(\mprj_logic1[449] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1307 (.DIODE(\mprj_logic1[449] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1308 (.DIODE(\mprj_logic1[449] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1309 (.DIODE(\mprj_logic1[449] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1310 (.DIODE(\mprj_logic1[449] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1311 (.DIODE(\mprj_logic1[449] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1312 (.DIODE(\mprj_logic1[449] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1313 (.DIODE(\mprj_logic1[449] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1314 (.DIODE(\mprj_logic1[449] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1315 (.DIODE(\mprj_logic1[449] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1316 (.DIODE(\mprj_logic1[449] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1317 (.DIODE(\mprj_logic1[449] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1318 (.DIODE(\mprj_logic1[449] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1319 (.DIODE(\mprj_logic1[449] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1320 (.DIODE(\mprj_logic1[449] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1321 (.DIODE(\mprj_logic1[449] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1322 (.DIODE(\mprj_logic1[449] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1323 (.DIODE(\mprj_logic1[449] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1324 (.DIODE(\mprj_logic1[450] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1325 (.DIODE(\mprj_logic1[450] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1326 (.DIODE(\mprj_logic1[451] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1327 (.DIODE(\mprj_logic1[451] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1328 (.DIODE(\mprj_logic1[452] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1329 (.DIODE(\mprj_logic1[452] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1330 (.DIODE(\mprj_logic1[454] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1331 (.DIODE(\mprj_logic1[454] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1332 (.DIODE(\mprj_logic1[454] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1333 (.DIODE(\mprj_logic1[454] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1334 (.DIODE(\mprj_logic1[454] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1335 (.DIODE(\mprj_logic1[454] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1336 (.DIODE(\mprj_logic1[454] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1337 (.DIODE(\mprj_logic1[454] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1338 (.DIODE(\mprj_logic1[454] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1339 (.DIODE(\mprj_logic1[454] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1340 (.DIODE(\mprj_logic1[454] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1341 (.DIODE(\mprj_logic1[454] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1342 (.DIODE(\mprj_logic1[454] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1343 (.DIODE(\mprj_logic1[454] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1344 (.DIODE(\mprj_logic1[454] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1345 (.DIODE(\mprj_logic1[454] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1346 (.DIODE(\mprj_logic1[456] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1347 (.DIODE(\mprj_logic1[456] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1348 (.DIODE(\mprj_logic1[456] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1349 (.DIODE(\mprj_logic1[456] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1350 (.DIODE(\mprj_logic1[456] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1351 (.DIODE(\mprj_logic1[457] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1352 (.DIODE(\mprj_logic1[457] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1353 (.DIODE(\mprj_logic1[458] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1354 (.DIODE(\mprj_logic1[458] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1355 (.DIODE(\mprj_logic1[458] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1356 (.DIODE(\mprj_logic1[458] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1357 (.DIODE(\mprj_logic1[458] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1358 (.DIODE(\mprj_logic1[458] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1359 (.DIODE(\mprj_logic1[458] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1360 (.DIODE(\mprj_logic1[458] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1361 (.DIODE(\mprj_logic1[458] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1362 (.DIODE(\mprj_logic1[458] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1363 (.DIODE(\mprj_logic1[458] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1364 (.DIODE(\mprj_logic1[459] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1365 (.DIODE(\mprj_logic1[459] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1366 (.DIODE(\mprj_logic1[460] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1367 (.DIODE(\mprj_logic1[460] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1368 (.DIODE(\mprj_logic1[462] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1369 (.DIODE(\mprj_logic1[462] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1370 (.DIODE(\mprj_logic1[47] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1371 (.DIODE(\mprj_logic1[48] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1372 (.DIODE(\mprj_logic1[49] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1373 (.DIODE(\mprj_logic1[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1374 (.DIODE(\mprj_logic1[50] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1375 (.DIODE(\mprj_logic1[51] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1376 (.DIODE(\mprj_logic1[52] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1377 (.DIODE(\mprj_logic1[54] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1378 (.DIODE(\mprj_logic1[55] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1379 (.DIODE(\mprj_logic1[57] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1380 (.DIODE(\mprj_logic1[58] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1381 (.DIODE(\mprj_logic1[59] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1382 (.DIODE(\mprj_logic1[60] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1383 (.DIODE(\mprj_logic1[61] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1384 (.DIODE(\mprj_logic1[64] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1385 (.DIODE(\mprj_logic1[66] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1386 (.DIODE(\mprj_logic1[67] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1387 (.DIODE(\mprj_logic1[68] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1388 (.DIODE(\mprj_logic1[69] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1389 (.DIODE(\mprj_logic1[70] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1390 (.DIODE(\mprj_logic1[70] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1391 (.DIODE(\mprj_logic1[70] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1392 (.DIODE(\mprj_logic1[70] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1393 (.DIODE(\mprj_logic1[70] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1394 (.DIODE(\mprj_logic1[70] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1395 (.DIODE(\mprj_logic1[70] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1396 (.DIODE(\mprj_logic1[70] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1397 (.DIODE(\mprj_logic1[70] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1398 (.DIODE(\mprj_logic1[70] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1399 (.DIODE(\mprj_logic1[70] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1400 (.DIODE(\mprj_logic1[70] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1401 (.DIODE(\mprj_logic1[70] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1402 (.DIODE(\mprj_logic1[70] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1403 (.DIODE(\mprj_logic1[72] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1404 (.DIODE(\mprj_logic1[72] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1405 (.DIODE(\mprj_logic1[72] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1406 (.DIODE(\mprj_logic1[72] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1407 (.DIODE(\mprj_logic1[72] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1408 (.DIODE(\mprj_logic1[72] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1409 (.DIODE(\mprj_logic1[72] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1410 (.DIODE(\mprj_logic1[72] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1411 (.DIODE(\mprj_logic1[72] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1412 (.DIODE(\mprj_logic1[72] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1413 (.DIODE(\mprj_logic1[72] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1414 (.DIODE(\mprj_logic1[72] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1415 (.DIODE(\mprj_logic1[72] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1416 (.DIODE(\mprj_logic1[72] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1417 (.DIODE(\mprj_logic1[73] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1418 (.DIODE(\mprj_logic1[73] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1419 (.DIODE(\mprj_logic1[73] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1420 (.DIODE(\mprj_logic1[73] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1421 (.DIODE(\mprj_logic1[73] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1422 (.DIODE(\mprj_logic1[73] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1423 (.DIODE(\mprj_logic1[73] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1424 (.DIODE(\mprj_logic1[73] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1425 (.DIODE(\mprj_logic1[73] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1426 (.DIODE(\mprj_logic1[73] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1427 (.DIODE(\mprj_logic1[73] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1428 (.DIODE(\mprj_logic1[73] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1429 (.DIODE(\mprj_logic1[73] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1430 (.DIODE(\mprj_logic1[73] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1431 (.DIODE(\mprj_logic1[73] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1432 (.DIODE(\mprj_logic1[73] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1433 (.DIODE(\mprj_logic1[74] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1434 (.DIODE(\mprj_logic1[74] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1435 (.DIODE(\mprj_logic1[74] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1436 (.DIODE(\mprj_logic1[74] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1437 (.DIODE(\mprj_logic1[74] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1438 (.DIODE(\mprj_logic1[75] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1439 (.DIODE(\mprj_logic1[75] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1440 (.DIODE(\mprj_logic1[75] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1441 (.DIODE(\mprj_logic1[76] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1442 (.DIODE(\mprj_logic1[76] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1443 (.DIODE(\mprj_logic1[76] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1444 (.DIODE(\mprj_logic1[76] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1445 (.DIODE(\mprj_logic1[76] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1446 (.DIODE(\mprj_logic1[77] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1447 (.DIODE(\mprj_logic1[77] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1448 (.DIODE(\mprj_logic1[77] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1449 (.DIODE(\mprj_logic1[77] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1450 (.DIODE(\mprj_logic1[77] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1451 (.DIODE(\mprj_logic1[77] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1452 (.DIODE(\mprj_logic1[78] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1453 (.DIODE(\mprj_logic1[78] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1454 (.DIODE(\mprj_logic1[78] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1455 (.DIODE(\mprj_logic1[79] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1456 (.DIODE(\mprj_logic1[79] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1457 (.DIODE(\mprj_logic1[79] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1458 (.DIODE(\mprj_logic1[80] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1459 (.DIODE(\mprj_logic1[80] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1460 (.DIODE(\mprj_logic1[81] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1461 (.DIODE(\mprj_logic1[81] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1462 (.DIODE(\mprj_logic1[81] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1463 (.DIODE(\mprj_logic1[81] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1464 (.DIODE(\mprj_logic1[81] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1465 (.DIODE(\mprj_logic1[81] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1466 (.DIODE(\mprj_logic1[81] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1467 (.DIODE(\mprj_logic1[81] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1468 (.DIODE(\mprj_logic1[81] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1469 (.DIODE(\mprj_logic1[81] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1470 (.DIODE(\mprj_logic1[81] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1471 (.DIODE(\mprj_logic1[81] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1472 (.DIODE(\mprj_logic1[81] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1473 (.DIODE(\mprj_logic1[81] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1474 (.DIODE(\mprj_logic1[81] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1475 (.DIODE(\mprj_logic1[81] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1476 (.DIODE(\mprj_logic1[81] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1477 (.DIODE(\mprj_logic1[81] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1478 (.DIODE(\mprj_logic1[81] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1479 (.DIODE(\mprj_logic1[81] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1480 (.DIODE(\mprj_logic1[82] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1481 (.DIODE(\mprj_logic1[82] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1482 (.DIODE(\mprj_logic1[82] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1483 (.DIODE(\mprj_logic1[82] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1484 (.DIODE(\mprj_logic1[82] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1485 (.DIODE(\mprj_logic1[82] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1486 (.DIODE(\mprj_logic1[82] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1487 (.DIODE(\mprj_logic1[82] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1488 (.DIODE(\mprj_logic1[82] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1489 (.DIODE(\mprj_logic1[82] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1490 (.DIODE(\mprj_logic1[82] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1491 (.DIODE(\mprj_logic1[82] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1492 (.DIODE(\mprj_logic1[82] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1493 (.DIODE(\mprj_logic1[82] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1494 (.DIODE(\mprj_logic1[82] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1495 (.DIODE(\mprj_logic1[82] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1496 (.DIODE(\mprj_logic1[82] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1497 (.DIODE(\mprj_logic1[82] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1498 (.DIODE(\mprj_logic1[82] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1499 (.DIODE(\mprj_logic1[82] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1500 (.DIODE(\mprj_logic1[84] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1501 (.DIODE(\mprj_logic1[84] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1502 (.DIODE(\mprj_logic1[85] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1503 (.DIODE(\mprj_logic1[86] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1504 (.DIODE(\mprj_logic1[86] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1505 (.DIODE(\mprj_logic1[86] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1506 (.DIODE(\mprj_logic1[86] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1507 (.DIODE(\mprj_logic1[86] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1508 (.DIODE(\mprj_logic1[86] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1509 (.DIODE(\mprj_logic1[86] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1510 (.DIODE(\mprj_logic1[86] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1511 (.DIODE(\mprj_logic1[86] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1512 (.DIODE(\mprj_logic1[86] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1513 (.DIODE(\mprj_logic1[86] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1514 (.DIODE(\mprj_logic1[86] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1515 (.DIODE(\mprj_logic1[86] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1516 (.DIODE(\mprj_logic1[88] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1517 (.DIODE(\mprj_logic1[88] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1518 (.DIODE(\mprj_logic1[88] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1519 (.DIODE(\mprj_logic1[88] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1520 (.DIODE(\mprj_logic1[88] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1521 (.DIODE(\mprj_logic1[88] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1522 (.DIODE(\mprj_logic1[88] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1523 (.DIODE(\mprj_logic1[88] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1524 (.DIODE(\mprj_logic1[88] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1525 (.DIODE(\mprj_logic1[88] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1526 (.DIODE(\mprj_logic1[88] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1527 (.DIODE(\mprj_logic1[88] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1528 (.DIODE(\mprj_logic1[88] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1529 (.DIODE(\mprj_logic1[88] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1530 (.DIODE(\mprj_logic1[89] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1531 (.DIODE(\mprj_logic1[89] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1532 (.DIODE(\mprj_logic1[89] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1533 (.DIODE(\mprj_logic1[89] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1534 (.DIODE(\mprj_logic1[89] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1535 (.DIODE(\mprj_logic1[89] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1536 (.DIODE(\mprj_logic1[89] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1537 (.DIODE(\mprj_logic1[89] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1538 (.DIODE(\mprj_logic1[89] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1539 (.DIODE(\mprj_logic1[89] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1540 (.DIODE(\mprj_logic1[91] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1541 (.DIODE(\mprj_logic1[91] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1542 (.DIODE(\mprj_logic1[91] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1543 (.DIODE(\mprj_logic1[91] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1544 (.DIODE(\mprj_logic1[91] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1545 (.DIODE(\mprj_logic1[91] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1546 (.DIODE(\mprj_logic1[91] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1547 (.DIODE(\mprj_logic1[91] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1548 (.DIODE(\mprj_logic1[91] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1549 (.DIODE(\mprj_logic1[91] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1550 (.DIODE(\mprj_logic1[91] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1551 (.DIODE(\mprj_logic1[91] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1552 (.DIODE(\mprj_logic1[91] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1553 (.DIODE(\mprj_logic1[91] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1554 (.DIODE(\mprj_logic1[92] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1555 (.DIODE(\mprj_logic1[92] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1556 (.DIODE(\mprj_logic1[92] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1557 (.DIODE(\mprj_logic1[92] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1558 (.DIODE(\mprj_logic1[95] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1559 (.DIODE(\mprj_logic1[95] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1560 (.DIODE(\mprj_logic1[96] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1561 (.DIODE(\mprj_logic1[96] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1562 (.DIODE(\mprj_logic1[97] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1563 (.DIODE(\mprj_logic1[97] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1564 (.DIODE(\mprj_logic1[97] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1565 (.DIODE(\mprj_logic1[97] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1566 (.DIODE(\mprj_logic1[97] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1567 (.DIODE(\mprj_logic1[97] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1568 (.DIODE(\mprj_logic1[99] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1569 (.DIODE(\mprj_logic1[99] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1570 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_1571 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_1572 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_1573 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_1574 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_1575 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_1576 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_1577 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_1578 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_1579 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_1580 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_1581 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_1582 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_1583 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_1584 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_1585 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_1586 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_1587 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_1588 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_1589 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_1590 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_1591 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_1592 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_1593 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_1594 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_1595 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_1596 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_1597 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_1598 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_1599 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_1600 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_1601 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_1602 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_1603 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_1604 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_1605 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_1606 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_1607 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_1608 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_1609 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_1610 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA_1611 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA_1612 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_1613 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_1614 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_1615 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_1616 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_1617 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_1618 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_1619 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_1620 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_1621 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_1622 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_1623 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_1624 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_1625 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_1626 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_1627 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_1628 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_1629 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_1630 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_1631 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_1632 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_1633 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_1634 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_1635 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_1636 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA_1637 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA_1638 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_1639 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_1640 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_1641 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_1642 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_1643 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_1644 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_1645 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_1646 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA_1647 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA_1648 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_1649 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_1650 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_1651 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_1652 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_1653 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_1654 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_1655 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_1656 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_1657 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_1658 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_1659 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_1660 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_1661 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_1662 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_1663 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_1664 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_1665 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_1666 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_1667 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_1668 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_1669 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_1670 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_1671 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_1672 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_1673 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_1674 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_1675 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_1676 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_1677 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_1678 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_1679 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_1680 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_1681 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_1682 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_1683 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_1684 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_1685 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_1686 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_1687 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_1688 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_1689 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_1690 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_1691 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_1692 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_1693 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_1694 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_1695 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_1696 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_1697 (.DIODE(net391));
 sky130_fd_sc_hd__diode_2 ANTENNA_1698 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_1699 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_1700 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_1701 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_1702 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_1703 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_1704 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_1705 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_1706 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_1707 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_1708 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_1709 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_1710 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_1711 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_1712 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_1713 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_1714 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_1715 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_1716 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_1717 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_1718 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_1719 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_1720 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_1721 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_1722 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_1723 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_1724 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_1725 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_1726 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_1727 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_1728 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_1729 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_1730 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_1731 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_1732 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_1733 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_1734 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_1735 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_1736 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_1737 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_1738 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_1739 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_1740 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_1741 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_1742 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_1743 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_1744 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_1745 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_1746 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_1747 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_1748 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_1749 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_1750 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_1751 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_1752 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_1753 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_1754 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_1755 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_1756 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_1757 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_1758 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_1759 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_1760 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_1761 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_1762 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_1763 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_1764 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_1765 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_1766 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_1767 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_1768 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_1769 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_1770 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_1771 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_1772 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_1773 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_1774 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_1775 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_1776 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_1777 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_1778 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_1779 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_1780 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_1781 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_1782 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_1783 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_1784 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_1785 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_1786 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_1787 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_1788 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_1789 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_1790 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_1791 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_1792 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_1793 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_1794 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_1795 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_1796 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_1797 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_1798 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_1799 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_1800 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_1801 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_1802 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_1803 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_1804 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_1805 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_1806 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_1807 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_1808 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_1809 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_1810 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_1811 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_1812 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_1813 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_1814 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_1815 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_1816 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_1817 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_1818 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_1819 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_1820 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_1821 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_1822 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_1823 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_1824 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_1825 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_1826 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_1827 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_1828 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_1829 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_1830 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_1831 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_1832 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_1833 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_1834 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_1835 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_1836 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_1837 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_1838 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_1839 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_1840 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_1841 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_1842 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_1843 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_1844 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_1845 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_1846 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_1847 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_1848 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_1849 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_1850 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_1851 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_1852 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_1853 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_1854 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_1855 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_1856 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_1857 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_1858 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_1859 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_1860 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_1861 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_1862 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_1863 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_1864 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_1865 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_1866 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_1867 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_1868 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_1869 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_1870 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_1871 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_1872 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_1873 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_1874 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_1875 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_1876 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_1877 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_1878 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_1879 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_1880 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_1881 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_1882 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_1883 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_1884 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_1885 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_1886 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_1887 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_1888 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_1889 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_1890 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_1891 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_1892 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_1893 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_1894 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_1895 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_1896 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_1897 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_1898 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_1899 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_1900 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_1901 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_1902 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_1903 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_1904 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_1905 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_1906 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_1907 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_1908 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_1909 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_1910 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_1911 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_1912 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_1913 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_1914 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_1915 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_1916 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_1917 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_1918 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_1919 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_1920 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_1921 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_1922 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_1923 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_1924 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_1925 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_1926 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_1927 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_1928 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_1929 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_1930 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_1931 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_1932 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_1933 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_1934 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_1935 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_1936 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_1937 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_1938 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_1939 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_1940 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_1941 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_1942 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_1943 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_1944 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_1945 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_1946 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_1947 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_1948 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_1949 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_1950 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_1951 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_1952 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_1953 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_1954 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_1955 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_1956 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_1957 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_1958 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_1959 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_1960 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_1961 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_1962 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_1963 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_1964 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_1965 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_1966 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_1967 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_1968 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_1969 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_1970 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA_1971 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_1972 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_1973 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA_1974 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_1975 (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA_1976 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_1977 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_1978 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_1979 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_1980 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_1981 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_1982 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA_1983 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_1984 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_1985 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_1986 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_1987 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_1988 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_1989 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_1990 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_1991 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_1992 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_1993 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_1994 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_1995 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_1996 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_1997 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_1998 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_1999 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_2000 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_2001 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_2002 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_2003 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_2004 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_2005 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_2006 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_2007 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_2008 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_2009 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_2010 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_2011 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_2012 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_2013 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_2014 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_2015 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_2016 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_2017 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_2018 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_2019 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_2020 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_2021 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_2022 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_2023 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_2024 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_2025 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_2026 (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA_2027 (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_2028 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_2029 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_2030 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_2031 (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_2032 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_2033 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_2034 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_2035 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA_2036 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_2037 (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_2038 (.DIODE(net837));
 sky130_fd_sc_hd__diode_2 ANTENNA_2039 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_2040 (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_2041 (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA_2042 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_2043 (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_2044 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_2045 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_2046 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_2047 (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_2048 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_2049 (.DIODE(net917));
 sky130_fd_sc_hd__diode_2 ANTENNA_2050 (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_2051 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_2052 (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_2053 (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_2054 (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_2055 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_2056 (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_2057 (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_2058 (.DIODE(net950));
 sky130_fd_sc_hd__diode_2 ANTENNA_2059 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_2060 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_2061 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_2062 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_2063 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_2064 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_2065 (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_2066 (.DIODE(\la_data_in_mprj_bar[86] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2067 (.DIODE(\la_data_in_mprj_bar[87] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2068 (.DIODE(\la_data_in_mprj_bar[90] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2069 (.DIODE(\la_data_in_mprj_bar[91] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2070 (.DIODE(la_data_out_core[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2071 (.DIODE(la_data_out_core[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2072 (.DIODE(mprj_dat_i_user[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2073 (.DIODE(mprj_dat_i_user[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2074 (.DIODE(\mprj_logic1[124] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2075 (.DIODE(\mprj_logic1[177] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2076 (.DIODE(\mprj_logic1[177] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2077 (.DIODE(\mprj_logic1[177] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2078 (.DIODE(\mprj_logic1[177] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2079 (.DIODE(\mprj_logic1[177] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2080 (.DIODE(\mprj_logic1[177] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2081 (.DIODE(\mprj_logic1[177] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2082 (.DIODE(\mprj_logic1[177] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2083 (.DIODE(\mprj_logic1[178] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2084 (.DIODE(\mprj_logic1[178] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2085 (.DIODE(\mprj_logic1[178] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2086 (.DIODE(\mprj_logic1[178] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2087 (.DIODE(\mprj_logic1[178] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2088 (.DIODE(\mprj_logic1[178] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2089 (.DIODE(\mprj_logic1[182] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2090 (.DIODE(\mprj_logic1[182] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2091 (.DIODE(\mprj_logic1[182] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2092 (.DIODE(\mprj_logic1[182] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2093 (.DIODE(\mprj_logic1[182] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2094 (.DIODE(\mprj_logic1[182] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2095 (.DIODE(\mprj_logic1[182] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2096 (.DIODE(\mprj_logic1[182] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2097 (.DIODE(\mprj_logic1[182] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2098 (.DIODE(\mprj_logic1[182] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2099 (.DIODE(\mprj_logic1[182] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2100 (.DIODE(\mprj_logic1[192] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2101 (.DIODE(\mprj_logic1[192] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2102 (.DIODE(\mprj_logic1[192] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2103 (.DIODE(\mprj_logic1[192] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2104 (.DIODE(\mprj_logic1[192] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2105 (.DIODE(\mprj_logic1[192] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2106 (.DIODE(\mprj_logic1[192] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2107 (.DIODE(\mprj_logic1[243] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2108 (.DIODE(\mprj_logic1[244] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2109 (.DIODE(\mprj_logic1[251] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2110 (.DIODE(\mprj_logic1[332] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2111 (.DIODE(\mprj_logic1[332] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2112 (.DIODE(\mprj_logic1[332] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2113 (.DIODE(\mprj_logic1[332] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2114 (.DIODE(\mprj_logic1[333] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2115 (.DIODE(\mprj_logic1[333] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2116 (.DIODE(\mprj_logic1[333] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2117 (.DIODE(\mprj_logic1[333] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2118 (.DIODE(\mprj_logic1[333] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2119 (.DIODE(\mprj_logic1[334] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2120 (.DIODE(\mprj_logic1[334] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2121 (.DIODE(\mprj_logic1[334] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2122 (.DIODE(\mprj_logic1[334] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2123 (.DIODE(\mprj_logic1[334] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2124 (.DIODE(\mprj_logic1[334] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2125 (.DIODE(\mprj_logic1[338] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2126 (.DIODE(\mprj_logic1[354] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2127 (.DIODE(\mprj_logic1[360] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2128 (.DIODE(\mprj_logic1[360] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2129 (.DIODE(\mprj_logic1[362] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2130 (.DIODE(\mprj_logic1[362] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2131 (.DIODE(\mprj_logic1[362] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2132 (.DIODE(\mprj_logic1[362] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2133 (.DIODE(\mprj_logic1[371] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2134 (.DIODE(\mprj_logic1[385] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2135 (.DIODE(\mprj_logic1[385] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2136 (.DIODE(\mprj_logic1[427] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2137 (.DIODE(\mprj_logic1[427] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2138 (.DIODE(\mprj_logic1[427] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2139 (.DIODE(\mprj_logic1[427] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2140 (.DIODE(\mprj_logic1[427] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2141 (.DIODE(\mprj_logic1[427] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2142 (.DIODE(\mprj_logic1[441] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2143 (.DIODE(\mprj_logic1[441] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2144 (.DIODE(\mprj_logic1[441] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2145 (.DIODE(\mprj_logic1[441] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2146 (.DIODE(\mprj_logic1[441] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2147 (.DIODE(\mprj_logic1[441] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2148 (.DIODE(\mprj_logic1[441] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2149 (.DIODE(\mprj_logic1[441] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2150 (.DIODE(\mprj_logic1[441] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2151 (.DIODE(\mprj_logic1[441] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2152 (.DIODE(\mprj_logic1[445] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2153 (.DIODE(\mprj_logic1[445] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2154 (.DIODE(\mprj_logic1[445] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2155 (.DIODE(\mprj_logic1[445] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2156 (.DIODE(\mprj_logic1[445] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2157 (.DIODE(\mprj_logic1[445] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2158 (.DIODE(\mprj_logic1[445] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2159 (.DIODE(\mprj_logic1[445] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2160 (.DIODE(\mprj_logic1[447] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2161 (.DIODE(\mprj_logic1[447] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2162 (.DIODE(\mprj_logic1[447] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2163 (.DIODE(\mprj_logic1[447] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2164 (.DIODE(\mprj_logic1[447] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2165 (.DIODE(\mprj_logic1[447] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2166 (.DIODE(\mprj_logic1[447] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2167 (.DIODE(\mprj_logic1[447] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2168 (.DIODE(\mprj_logic1[447] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2169 (.DIODE(\mprj_logic1[447] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2170 (.DIODE(\mprj_logic1[449] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2171 (.DIODE(\mprj_logic1[449] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2172 (.DIODE(\mprj_logic1[449] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2173 (.DIODE(\mprj_logic1[449] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2174 (.DIODE(\mprj_logic1[449] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2175 (.DIODE(\mprj_logic1[449] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2176 (.DIODE(\mprj_logic1[449] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2177 (.DIODE(\mprj_logic1[449] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2178 (.DIODE(\mprj_logic1[449] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2179 (.DIODE(\mprj_logic1[449] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2180 (.DIODE(\mprj_logic1[449] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2181 (.DIODE(\mprj_logic1[449] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2182 (.DIODE(\mprj_logic1[452] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2183 (.DIODE(\mprj_logic1[452] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2184 (.DIODE(\mprj_logic1[452] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2185 (.DIODE(\mprj_logic1[452] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2186 (.DIODE(\mprj_logic1[452] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2187 (.DIODE(\mprj_logic1[452] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2188 (.DIODE(\mprj_logic1[452] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2189 (.DIODE(\mprj_logic1[452] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2190 (.DIODE(\mprj_logic1[452] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2191 (.DIODE(\mprj_logic1[452] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2192 (.DIODE(\mprj_logic1[452] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2193 (.DIODE(\mprj_logic1[452] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2194 (.DIODE(\mprj_logic1[452] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2195 (.DIODE(\mprj_logic1[452] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2196 (.DIODE(\mprj_logic1[456] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2197 (.DIODE(\mprj_logic1[456] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2198 (.DIODE(\mprj_logic1[456] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2199 (.DIODE(\mprj_logic1[456] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2200 (.DIODE(\mprj_logic1[456] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2201 (.DIODE(\mprj_logic1[456] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2202 (.DIODE(\mprj_logic1[456] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2203 (.DIODE(\mprj_logic1[456] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2204 (.DIODE(\mprj_logic1[456] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2205 (.DIODE(\mprj_logic1[456] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2206 (.DIODE(\mprj_logic1[456] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2207 (.DIODE(\mprj_logic1[456] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2208 (.DIODE(\mprj_logic1[458] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2209 (.DIODE(\mprj_logic1[458] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2210 (.DIODE(\mprj_logic1[458] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2211 (.DIODE(\mprj_logic1[458] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2212 (.DIODE(\mprj_logic1[458] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2213 (.DIODE(\mprj_logic1[458] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2214 (.DIODE(\mprj_logic1[458] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2215 (.DIODE(\mprj_logic1[458] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2216 (.DIODE(\mprj_logic1[458] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2217 (.DIODE(\mprj_logic1[458] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2218 (.DIODE(\mprj_logic1[458] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2219 (.DIODE(\mprj_logic1[458] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2220 (.DIODE(\mprj_logic1[460] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2221 (.DIODE(\mprj_logic1[460] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2222 (.DIODE(\mprj_logic1[460] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2223 (.DIODE(\mprj_logic1[460] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2224 (.DIODE(\mprj_logic1[460] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2225 (.DIODE(\mprj_logic1[460] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2226 (.DIODE(\mprj_logic1[460] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2227 (.DIODE(\mprj_logic1[460] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2228 (.DIODE(\mprj_logic1[460] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2229 (.DIODE(\mprj_logic1[460] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2230 (.DIODE(\mprj_logic1[460] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2231 (.DIODE(\mprj_logic1[460] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2232 (.DIODE(\mprj_logic1[460] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2233 (.DIODE(\mprj_logic1[460] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2234 (.DIODE(\mprj_logic1[460] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2235 (.DIODE(\mprj_logic1[460] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2236 (.DIODE(\mprj_logic1[460] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2237 (.DIODE(\mprj_logic1[460] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2238 (.DIODE(\mprj_logic1[460] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2239 (.DIODE(\mprj_logic1[460] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2240 (.DIODE(\mprj_logic1[460] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2241 (.DIODE(\mprj_logic1[460] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2242 (.DIODE(\mprj_logic1[87] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2243 (.DIODE(\mprj_logic1[93] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2244 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_2245 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_2246 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_2247 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_2248 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA_2249 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_2250 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_2251 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_2252 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_2253 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_2254 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_2255 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_2256 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_2257 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_2258 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_2259 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_2260 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_2261 (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_2262 (.DIODE(net926));
 sky130_fd_sc_hd__diode_2 ANTENNA_2263 (.DIODE(net927));
 sky130_fd_sc_hd__diode_2 ANTENNA_2264 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_2265 (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_2266 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_2267 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_2268 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_2269 (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_2270 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_2271 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_2272 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_2273 (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_2274 (.DIODE(la_data_out_core[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2275 (.DIODE(la_data_out_core[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2276 (.DIODE(mprj_dat_i_user[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2277 (.DIODE(mprj_dat_i_user[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2278 (.DIODE(mprj_dat_i_user[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2279 (.DIODE(mprj_dat_i_user[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2280 (.DIODE(mprj_dat_i_user[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2281 (.DIODE(mprj_dat_i_user[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2282 (.DIODE(mprj_dat_i_user[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2283 (.DIODE(mprj_dat_i_user[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2284 (.DIODE(mprj_dat_i_user[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2285 (.DIODE(mprj_dat_i_user[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2286 (.DIODE(mprj_dat_i_user[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2287 (.DIODE(mprj_dat_i_user[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2288 (.DIODE(mprj_dat_i_user[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2289 (.DIODE(mprj_dat_i_user[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2290 (.DIODE(mprj_dat_i_user[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2291 (.DIODE(mprj_dat_i_user[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2292 (.DIODE(mprj_dat_i_user[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2293 (.DIODE(mprj_dat_i_user[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2294 (.DIODE(mprj_dat_i_user[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2295 (.DIODE(mprj_dat_i_user[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2296 (.DIODE(mprj_dat_i_user[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2297 (.DIODE(mprj_dat_i_user[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2298 (.DIODE(mprj_dat_i_user[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2299 (.DIODE(mprj_dat_i_user[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2300 (.DIODE(mprj_dat_i_user[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2301 (.DIODE(mprj_dat_i_user[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2302 (.DIODE(mprj_dat_i_user[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2303 (.DIODE(mprj_dat_i_user[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2304 (.DIODE(mprj_dat_i_user[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2305 (.DIODE(mprj_dat_i_user[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2306 (.DIODE(mprj_dat_i_user[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2307 (.DIODE(mprj_dat_i_user[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2308 (.DIODE(mprj_dat_i_user[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2309 (.DIODE(mprj_dat_i_user[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2310 (.DIODE(mprj_dat_i_user[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2311 (.DIODE(mprj_dat_i_user[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2312 (.DIODE(mprj_dat_i_user[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2313 (.DIODE(mprj_dat_i_user[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2314 (.DIODE(mprj_dat_i_user[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2315 (.DIODE(mprj_dat_i_user[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2316 (.DIODE(mprj_dat_i_user[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2317 (.DIODE(mprj_dat_i_user[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2318 (.DIODE(mprj_dat_i_user[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2319 (.DIODE(mprj_dat_i_user[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2320 (.DIODE(mprj_dat_i_user[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2321 (.DIODE(mprj_dat_i_user[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2322 (.DIODE(mprj_dat_i_user[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2323 (.DIODE(mprj_dat_i_user[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2324 (.DIODE(mprj_dat_i_user[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2325 (.DIODE(mprj_dat_i_user[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2326 (.DIODE(mprj_dat_i_user[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2327 (.DIODE(mprj_dat_i_user[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2328 (.DIODE(mprj_dat_i_user[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2329 (.DIODE(mprj_dat_i_user[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2330 (.DIODE(mprj_dat_i_user[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2331 (.DIODE(mprj_dat_i_user[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2332 (.DIODE(mprj_dat_i_user[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2333 (.DIODE(mprj_dat_i_user[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2334 (.DIODE(mprj_dat_i_user[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2335 (.DIODE(mprj_dat_i_user[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2336 (.DIODE(mprj_dat_i_user[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2337 (.DIODE(mprj_dat_i_user[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2338 (.DIODE(mprj_dat_i_user[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2339 (.DIODE(mprj_dat_i_user[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2340 (.DIODE(mprj_dat_i_user[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2341 (.DIODE(mprj_dat_i_user[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2342 (.DIODE(mprj_dat_i_user[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2343 (.DIODE(mprj_dat_i_user[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2344 (.DIODE(mprj_dat_i_user[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2345 (.DIODE(mprj_dat_i_user[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2346 (.DIODE(mprj_dat_i_user[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2347 (.DIODE(mprj_dat_i_user[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2348 (.DIODE(mprj_dat_i_user[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2349 (.DIODE(mprj_dat_i_user[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2350 (.DIODE(mprj_dat_i_user[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2351 (.DIODE(mprj_dat_i_user[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2352 (.DIODE(mprj_dat_i_user[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2353 (.DIODE(mprj_dat_i_user[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2354 (.DIODE(mprj_dat_i_user[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2355 (.DIODE(mprj_dat_i_user[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2356 (.DIODE(mprj_dat_i_user[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2357 (.DIODE(mprj_dat_i_user[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2358 (.DIODE(mprj_dat_i_user[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2359 (.DIODE(mprj_dat_i_user[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2360 (.DIODE(mprj_dat_i_user[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2361 (.DIODE(\mprj_logic1[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2362 (.DIODE(\mprj_logic1[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2363 (.DIODE(\mprj_logic1[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2364 (.DIODE(\mprj_logic1[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2365 (.DIODE(\mprj_logic1[159] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2366 (.DIODE(\mprj_logic1[159] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2367 (.DIODE(\mprj_logic1[159] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2368 (.DIODE(\mprj_logic1[159] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2369 (.DIODE(\mprj_logic1[159] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2370 (.DIODE(\mprj_logic1[159] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2371 (.DIODE(\mprj_logic1[159] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2372 (.DIODE(\mprj_logic1[159] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2373 (.DIODE(\mprj_logic1[159] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2374 (.DIODE(\mprj_logic1[159] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2375 (.DIODE(\mprj_logic1[159] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2376 (.DIODE(\mprj_logic1[211] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2377 (.DIODE(\mprj_logic1[211] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2378 (.DIODE(\mprj_logic1[211] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2379 (.DIODE(\mprj_logic1[211] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2380 (.DIODE(\mprj_logic1[211] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2381 (.DIODE(\mprj_logic1[211] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2382 (.DIODE(\mprj_logic1[211] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2383 (.DIODE(\mprj_logic1[211] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2384 (.DIODE(\mprj_logic1[211] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2385 (.DIODE(\mprj_logic1[211] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2386 (.DIODE(\mprj_logic1[211] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2387 (.DIODE(\mprj_logic1[211] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2388 (.DIODE(\mprj_logic1[240] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2389 (.DIODE(\mprj_logic1[35] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2390 (.DIODE(\mprj_logic1[40] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2391 (.DIODE(\mprj_logic1[438] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2392 (.DIODE(\mprj_logic1[438] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2393 (.DIODE(\mprj_logic1[438] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2394 (.DIODE(\mprj_logic1[438] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2395 (.DIODE(\mprj_logic1[438] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2396 (.DIODE(\mprj_logic1[438] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2397 (.DIODE(\mprj_logic1[438] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2398 (.DIODE(\mprj_logic1[438] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2399 (.DIODE(\mprj_logic1[438] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2400 (.DIODE(\mprj_logic1[457] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2401 (.DIODE(\mprj_logic1[457] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2402 (.DIODE(\mprj_logic1[457] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2403 (.DIODE(\mprj_logic1[457] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2404 (.DIODE(\mprj_logic1[457] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2405 (.DIODE(\mprj_logic1[457] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2406 (.DIODE(\mprj_logic1[457] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2407 (.DIODE(\mprj_logic1[457] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2408 (.DIODE(\mprj_logic1[457] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2409 (.DIODE(\mprj_logic1[457] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2410 (.DIODE(\mprj_logic1[457] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2411 (.DIODE(\mprj_logic1[457] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2412 (.DIODE(\mprj_logic1[457] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2413 (.DIODE(\mprj_logic1[457] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2414 (.DIODE(\mprj_logic1[459] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2415 (.DIODE(\mprj_logic1[459] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2416 (.DIODE(\mprj_logic1[459] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2417 (.DIODE(\mprj_logic1[459] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2418 (.DIODE(\mprj_logic1[459] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2419 (.DIODE(\mprj_logic1[459] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2420 (.DIODE(\mprj_logic1[459] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2421 (.DIODE(\mprj_logic1[459] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2422 (.DIODE(\mprj_logic1[459] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2423 (.DIODE(\mprj_logic1[459] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2424 (.DIODE(\mprj_logic1[459] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2425 (.DIODE(\mprj_logic1[459] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2426 (.DIODE(\mprj_logic1[459] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2427 (.DIODE(\mprj_logic1[459] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2428 (.DIODE(\mprj_logic1[459] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2429 (.DIODE(\mprj_logic1[459] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2430 (.DIODE(\mprj_logic1[459] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2431 (.DIODE(\mprj_logic1[459] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2432 (.DIODE(\mprj_logic1[459] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2433 (.DIODE(\mprj_logic1[459] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2434 (.DIODE(\mprj_logic1[459] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2435 (.DIODE(\mprj_logic1[459] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2436 (.DIODE(\mprj_logic1[62] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2437 (.DIODE(\mprj_logic1[63] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2438 (.DIODE(\mprj_logic1[65] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2439 (.DIODE(\mprj_logic1[71] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2440 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_2441 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_2442 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_2443 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_2444 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_2445 (.DIODE(mprj_dat_i_user[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2446 (.DIODE(mprj_dat_i_user[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2447 (.DIODE(mprj_dat_i_user[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2448 (.DIODE(mprj_dat_i_user[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2449 (.DIODE(mprj_dat_i_user[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2450 (.DIODE(mprj_dat_i_user[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2451 (.DIODE(mprj_dat_i_user[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2452 (.DIODE(mprj_dat_i_user[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2453 (.DIODE(mprj_dat_i_user[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2454 (.DIODE(mprj_dat_i_user[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2455 (.DIODE(mprj_dat_i_user[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2456 (.DIODE(mprj_dat_i_user[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2457 (.DIODE(mprj_dat_i_user[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2458 (.DIODE(mprj_dat_i_user[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2459 (.DIODE(\mprj_logic1[156] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2460 (.DIODE(\mprj_logic1[156] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2461 (.DIODE(\mprj_logic1[156] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2462 (.DIODE(\mprj_logic1[156] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2463 (.DIODE(\mprj_logic1[156] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2464 (.DIODE(\mprj_logic1[156] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2465 (.DIODE(\mprj_logic1[156] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2466 (.DIODE(\mprj_logic1[156] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2467 (.DIODE(\mprj_logic1[156] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2468 (.DIODE(\mprj_logic1[156] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2469 (.DIODE(\mprj_logic1[158] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2470 (.DIODE(\mprj_logic1[158] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2471 (.DIODE(\mprj_logic1[158] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2472 (.DIODE(\mprj_logic1[158] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2473 (.DIODE(\mprj_logic1[158] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2474 (.DIODE(\mprj_logic1[158] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2475 (.DIODE(\mprj_logic1[158] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2476 (.DIODE(\mprj_logic1[158] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2477 (.DIODE(\mprj_logic1[158] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2478 (.DIODE(\mprj_logic1[158] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2479 (.DIODE(\mprj_logic1[158] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2480 (.DIODE(\mprj_logic1[158] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2481 (.DIODE(\mprj_logic1[362] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2482 (.DIODE(\mprj_logic1[362] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2483 (.DIODE(\mprj_logic1[362] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2484 (.DIODE(\mprj_logic1[362] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2485 (.DIODE(\mprj_logic1[362] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2486 (.DIODE(\mprj_logic1[362] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2487 (.DIODE(\mprj_logic1[362] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2488 (.DIODE(\mprj_logic1[362] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2489 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_2490 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_2491 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_2492 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_2493 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_2494 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_2495 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_2496 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_2497 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_2498 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_2499 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_2500 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_2501 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_2502 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_2503 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_2504 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_2505 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_2506 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_2507 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_2508 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_2509 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_2510 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_2511 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_2512 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_2513 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_2514 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_2515 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_2516 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2517 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2518 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2519 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2520 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2521 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2522 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2523 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2524 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2525 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2526 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2527 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2528 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2529 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2530 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2531 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2532 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2533 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2534 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2535 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2536 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2537 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2538 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2539 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2540 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2541 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2542 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2543 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2544 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2545 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2546 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_2547 (.DIODE(\mprj_logic1[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2548 (.DIODE(\mprj_logic1[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2549 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_2550 (.DIODE(net778));
 sky130_fd_sc_hd__diode_2 ANTENNA_2551 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2552 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2553 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2554 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2555 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2556 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2557 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2558 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2559 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2560 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2561 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2562 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2563 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2564 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2565 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2566 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2567 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2568 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2569 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2570 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2571 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2572 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2573 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2574 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2575 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2576 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2577 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2578 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2579 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2580 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2581 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2582 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2583 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_2584 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_2585 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_2586 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_2587 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_2588 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_2589 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_2590 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_2591 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_2592 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_2593 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_2594 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_2595 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_2596 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_2597 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_2598 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_2599 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_2600 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_2601 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_2602 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_2603 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_2604 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_2605 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_2606 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_2607 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_2608 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_2609 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_2610 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_2611 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_2612 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_2613 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_2614 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_2615 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_2616 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_2617 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_2618 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_2619 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_2620 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_2621 (.DIODE(la_data_out_core[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2622 (.DIODE(\mprj_logic1[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2623 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_2624 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_2625 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_2626 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_2627 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_2628 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_2629 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_2630 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_2631 (.DIODE(net438));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_883 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_911 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_939 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_967 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1023 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1079 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1555 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1583 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1611 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1639 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1667 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1695 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1723 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1751 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1779 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1807 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1835 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1863 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1891 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1919 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1947 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1975 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2003 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2017 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2031 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2045 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2059 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2069 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2073 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2098 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2535 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2563 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2591 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2619 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2647 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2675 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2703 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2731 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2759 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2773 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2801 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2815 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2829 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2843 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2857 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2871 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2885 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2899 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2927 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2941 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2955 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2969 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2983 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2997 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3011 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3025 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3039 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3053 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3067 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3081 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3095 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3543 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3655 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3683 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3771 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3911 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3929 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3967 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4003 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4013 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4047 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4051 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4059 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4075 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4087 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4577 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1303 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1315 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1323 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1345 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1353 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1361 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1381 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1399 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1401 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1417 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1435 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1445 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1453 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1471 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1479 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1493 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1503 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1511 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1513 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1522 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1539 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1557 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1565 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1569 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1578 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1597 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1607 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1622 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1625 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1633 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1641 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1659 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1669 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1677 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1681 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1690 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1707 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1725 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1737 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1745 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1753 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1771 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1781 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1789 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1793 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1802 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1819 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1837 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1845 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1849 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1857 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1865 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1883 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1893 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1901 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1905 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1914 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1931 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1935 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1942 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1948 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1958 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1961 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1970 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1987 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1991 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2001 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2014 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_2017 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2029 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2033 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2043 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2047 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2057 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2070 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2073 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2087 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2095 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2122 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2129 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2143 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2151 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2178 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2185 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2199 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2207 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2221 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2231 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2239 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2241 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2255 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2263 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2277 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2287 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2295 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2311 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2323 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2327 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2334 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2346 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2353 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2367 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2383 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_2405 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2409 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2423 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2439 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2452 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2465 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2479 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2495 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2508 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2521 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2535 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2551 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2567 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2575 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2577 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2591 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2607 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2623 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2631 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2633 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2647 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2663 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2673 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2677 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2684 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_2689 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2698 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2712 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2726 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2732 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2742 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_2745 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2754 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2771 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2775 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2782 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2794 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2801 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2815 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2831 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_2853 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2857 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2871 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2884 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2894 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2900 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2910 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_2913 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2922 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2939 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2943 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2950 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2956 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2966 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_2969 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2978 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2995 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2999 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3006 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3010 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3022 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_3025 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_3034 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3051 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3055 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3062 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3068 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3078 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_3081 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_3090 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3107 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3111 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3118 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3124 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3134 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_3137 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_3146 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3163 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3167 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3174 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3180 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3190 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_3193 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_3202 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3219 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3223 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3230 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3236 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3246 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_3249 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_3258 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3275 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3279 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3286 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3292 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3302 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_3305 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3317 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3321 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3331 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3335 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3342 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3348 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3358 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_3361 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3373 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3377 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3387 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3391 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3398 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3404 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3414 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_3417 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_3426 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3443 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3447 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3454 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3460 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3470 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_3473 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_3482 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3499 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3503 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3510 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3516 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3526 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_3529 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_3538 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3555 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3559 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3566 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3572 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3582 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_3585 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_3594 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3611 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3615 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3622 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3628 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3638 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_3641 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3655 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3668 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3683 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3695 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_3697 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3711 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3730 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3734 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3738 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3742 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3746 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3750 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_3753 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3768 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3784 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3800 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3804 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_3809 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3814 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3818 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3821 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3825 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3829 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3833 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3837 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3841 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3855 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3859 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3863 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3865 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3869 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3873 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3877 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3881 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3895 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3899 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3903 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3907 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3911 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_3915 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3921 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3925 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3929 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3933 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3937 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3951 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3967 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_3971 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3977 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3981 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3985 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3989 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_4033 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_4047 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_4063 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_4079 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4087 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_4089 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_4103 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_4119 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_4135 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4143 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_4145 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_4159 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_4175 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_4191 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4199 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_4201 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_4215 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_4231 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_4247 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4255 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_4257 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_4271 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_4287 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_4303 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4311 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_4313 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_4327 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_4343 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_4359 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4367 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_4369 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_4383 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_4399 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4412 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4425 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4437 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4461 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_4473 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4479 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4481 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4493 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4517 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_4529 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4535 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4537 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4549 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_4561 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_4579 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1235 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1291 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1298 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1347 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1354 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1385 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1397 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1403 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1410 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1422 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1441 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1453 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1459 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1466 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1478 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1539 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1550 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1562 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1574 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1586 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1594 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1609 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1621 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1627 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1634 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1646 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1707 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1718 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1730 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1738 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1746 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1819 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1830 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1842 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1850 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1858 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2057 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2069 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2075 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2113 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2125 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2131 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2169 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2181 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2187 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2194 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2206 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2225 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2237 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2243 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2250 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2262 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2281 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2293 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2299 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2306 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2318 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2349 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_2361 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_2369 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2393 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2405 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2411 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2423 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2461 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2467 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2505 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2517 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2523 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2561 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2573 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2579 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2592 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2617 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2629 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2635 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2648 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2797 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_2809 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_2817 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2853 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_2865 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_2873 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2997 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3009 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3021 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3033 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3045 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3051 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3065 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3089 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3101 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3107 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3121 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3145 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3157 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3163 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3177 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3201 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3213 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3219 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3233 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3245 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3257 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3269 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3275 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3289 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3301 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3313 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3325 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3331 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3345 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3357 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3369 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3381 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3387 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3401 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3425 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3437 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3443 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3457 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3481 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3493 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3499 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3513 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3537 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3549 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3555 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3569 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3593 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3605 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3611 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3625 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3649 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3661 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3667 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3669 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3681 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3685 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3695 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3707 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3719 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3723 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3725 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_3739 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3757 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_3769 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_3777 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_3781 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3796 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3812 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3818 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3822 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3826 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3830 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3834 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_3837 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3852 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3868 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3872 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3876 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3880 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3884 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3888 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3893 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3897 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_3901 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3906 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3910 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3914 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3918 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3922 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3926 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3940 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3944 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3949 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3953 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3957 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3961 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_3965 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3980 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3996 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_4000 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_4005 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_4020 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_4036 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_4052 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_4061 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_4076 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_4092 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_4108 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_4117 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_4132 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_4148 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_4164 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_4173 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_4188 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_4204 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_4220 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_4229 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_4244 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_4260 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_4276 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_4285 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_4300 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_4316 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_4332 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_4341 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_4356 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_4372 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_4388 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_4397 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_4409 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4422 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4434 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_4446 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4453 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4465 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4489 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_4501 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4507 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4509 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4521 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4545 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_4557 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4563 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4565 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_4577 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3005 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3017 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3023 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3025 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3037 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3049 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3061 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3073 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3079 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3093 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3117 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3129 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3135 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3137 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3149 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3153 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3157 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3169 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3173 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3177 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3229 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3241 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3247 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3249 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3261 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3267 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3271 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3283 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_3295 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3303 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3317 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3329 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3341 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3353 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3359 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3373 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3397 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3409 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3415 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3429 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3453 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3465 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3471 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3497 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3509 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3521 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3527 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3541 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3565 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3577 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3583 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3597 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3621 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3633 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3639 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3653 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3677 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3689 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3695 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3709 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3733 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3745 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3751 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3765 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_3777 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_3785 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3790 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3794 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3798 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3802 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3809 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_3813 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3840 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3844 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3848 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3860 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3865 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3871 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3945 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_3967 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3972 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3977 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3982 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3989 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3993 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3997 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_4001 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_4005 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_4013 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_4017 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_4021 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4025 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4031 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4038 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4050 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4054 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4066 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4070 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4082 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_4089 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_4094 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4110 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4125 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4137 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4143 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4145 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4157 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4181 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4193 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4199 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4201 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4213 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4237 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4249 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4255 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4257 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4269 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4293 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4305 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4311 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4313 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_4325 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_4330 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_4339 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4343 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4355 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4367 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4369 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4381 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4405 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4417 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4423 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4425 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4437 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4461 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4473 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4479 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4481 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4493 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4517 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4529 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4535 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4537 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4549 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4561 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_4573 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2997 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3009 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3021 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3033 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3045 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3051 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3065 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3089 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3101 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3107 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3121 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3145 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3157 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3163 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3177 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3201 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3213 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3219 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3233 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3245 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3257 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3269 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3275 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3289 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3301 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3313 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3325 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3331 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3345 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3357 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3369 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3381 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3387 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3401 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3425 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3437 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3443 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3457 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3481 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3493 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3499 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3513 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3537 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3549 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3555 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3569 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3593 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3605 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3611 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3625 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3649 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3661 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3667 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3681 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3705 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3717 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3723 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3737 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3749 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3761 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3773 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3779 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3781 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3793 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3799 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3802 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3806 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3810 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3814 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3818 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3822 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3826 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3830 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3834 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3841 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3853 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3865 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3879 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3891 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3893 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_3905 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3913 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3917 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3921 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3935 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_3939 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3947 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3961 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3973 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3981 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3985 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3989 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3993 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3997 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4003 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4017 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4041 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4053 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4059 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4061 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4073 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_4082 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4090 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_4093 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_4097 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_4101 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_4105 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4109 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4115 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_4117 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_4123 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4131 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4134 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4146 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4158 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_4170 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4173 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4185 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4209 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4221 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4227 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4229 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4241 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4265 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4277 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4283 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4285 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4297 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4321 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4333 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4339 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4341 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4353 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4377 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4389 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4395 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4397 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4409 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4433 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4445 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4451 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4453 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4465 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4489 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4501 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4507 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4509 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4521 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4545 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4557 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4563 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_4565 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_4579 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3005 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3017 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3023 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3025 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3037 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3049 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3061 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3073 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3079 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3093 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3117 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3129 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3135 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3149 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3166 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3178 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3190 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3229 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3241 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3247 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3261 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3273 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3285 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3297 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3303 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3317 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3329 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3341 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3353 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3359 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3373 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3397 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3409 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3415 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3429 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3453 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3465 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3471 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3497 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3509 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3521 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3527 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3541 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3565 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3577 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3583 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3597 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3621 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3633 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3639 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3653 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3677 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3689 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3695 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3709 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3733 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3745 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3751 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3765 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3777 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3789 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3801 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3807 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3809 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3813 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3817 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_3821 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3826 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3830 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3834 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3846 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3858 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3865 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3877 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3889 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3901 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3913 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3919 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_3921 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3929 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3933 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3945 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_3957 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3967 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3971 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3975 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3977 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3985 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3989 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4013 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4025 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4031 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_4033 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4041 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_4045 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_4051 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_4055 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_4059 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_4063 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_4067 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_4071 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_4078 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_4082 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_4086 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_4089 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_4095 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_4099 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_4104 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_4108 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_4112 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_4116 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_4120 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_4124 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_4128 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_4132 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_4136 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_4140 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4145 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4157 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4181 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4193 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4199 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4201 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4213 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4237 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4249 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4255 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4257 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4269 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4293 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4305 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4311 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4313 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4325 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4349 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4361 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4367 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4369 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4381 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4405 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4417 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4423 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4425 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4437 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4461 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4473 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4479 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4481 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4493 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4517 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4529 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4535 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4537 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4549 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4561 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_4573 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2771 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_2773 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_2779 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2783 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2795 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2807 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_2819 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2997 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3011 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3023 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3035 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3047 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3051 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3065 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3089 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3101 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3107 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_3109 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3117 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3120 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3126 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_3138 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3148 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_3154 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3162 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3177 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3189 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3201 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_3211 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3219 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3233 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3245 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3257 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3269 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3275 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3289 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3301 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3313 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3325 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3331 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3345 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3357 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3369 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3381 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3387 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3401 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3425 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3437 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3443 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3457 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3481 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3493 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3499 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3513 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3537 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3549 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3555 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3569 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3593 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3605 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3611 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3625 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3649 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3661 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3667 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3681 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3705 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3717 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3723 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3737 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3749 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_3761 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3769 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3775 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3779 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3781 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3793 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3805 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3817 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3821 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3825 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3829 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3835 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3849 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3861 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3873 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3885 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3891 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3893 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3905 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3911 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3914 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3918 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3922 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3926 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3930 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3934 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3938 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3942 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3946 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_3949 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3954 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3959 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3963 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3967 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3971 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3975 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3979 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3983 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3989 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3993 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3997 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_4001 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_4005 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_4009 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4013 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4025 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4037 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_4049 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4061 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_4073 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4081 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4084 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_4096 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_4101 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_4105 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_4113 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_4117 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_4124 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4134 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4146 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4158 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_4170 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4173 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4185 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4209 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4221 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4227 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4229 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4241 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4265 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4277 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4283 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4285 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4297 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4321 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4333 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4339 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4341 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4353 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4377 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4389 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4395 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4397 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4409 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4433 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4445 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4451 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4453 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4465 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4489 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4501 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4507 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4509 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4521 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4545 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4557 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4563 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_4565 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_4579 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_986 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1973 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2477 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2713 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2717 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2725 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2734 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2742 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2749 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_2761 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2773 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_2792 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2825 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_2829 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2837 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2843 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2969 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2981 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2985 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2994 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_2997 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3005 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3008 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3020 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3025 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3037 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3049 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3065 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3093 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3121 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3149 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3177 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3205 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3233 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3245 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3261 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3273 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3289 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3301 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3317 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3329 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3345 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3357 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3373 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3401 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3429 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3457 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3469 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3478 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_3490 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3498 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3513 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3541 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3569 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3597 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3625 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3653 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3681 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3709 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3737 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3749 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3753 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3765 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3771 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3775 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3779 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3781 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3793 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3805 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3821 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3849 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3861 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3865 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3877 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3882 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3886 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3890 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3893 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3899 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3903 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3907 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3912 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3916 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3921 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3925 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3929 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3933 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3937 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3941 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3946 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3949 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3953 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3957 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3961 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3965 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3969 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3973 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3977 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3981 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3985 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3997 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4003 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4017 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4045 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_4057 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_4061 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_4070 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_4077 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_4084 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_4089 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4094 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_4106 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_4114 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4117 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_4129 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4133 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_4136 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_4145 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_4153 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4158 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_4170 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4173 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4185 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_4197 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4201 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4213 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_4225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4229 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4241 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_4253 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_4257 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4263 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_4275 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4283 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4285 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4297 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_4309 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4313 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4325 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_4337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4341 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4353 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_4365 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4369 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4381 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_4393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4397 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4409 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_4421 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4425 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4437 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_4449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4453 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4465 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_4477 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4481 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4493 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_4505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4509 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4521 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_4533 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4537 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4549 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_4561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4565 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_4577 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1016 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1067 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1123 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1179 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1235 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1267 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1279 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1291 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1323 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1335 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1347 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1367 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1379 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1391 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1403 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1423 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1435 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1447 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1459 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1471 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1479 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1491 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1503 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1515 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1529 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1535 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1547 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1559 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1571 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1583 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1591 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1603 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1615 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1627 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1635 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1640 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1644 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1647 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1659 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1671 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1683 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1695 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1703 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1715 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1727 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1739 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1751 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1757 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1759 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1766 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1778 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1790 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1802 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1815 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1827 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1839 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1851 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1863 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1869 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1871 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1883 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1895 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1907 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1919 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1927 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1939 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1951 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1963 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1975 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1981 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1983 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1988 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1992 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1996 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2000 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_2003 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2007 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2019 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2031 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2037 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2039 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2051 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2063 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2075 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2087 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2093 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2095 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2107 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2119 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2131 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2143 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2149 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2151 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2163 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2175 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2187 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2199 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2207 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2219 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2231 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2243 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2255 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2261 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2263 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2275 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2287 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2299 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2311 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2317 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2319 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2331 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2343 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2355 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2367 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2373 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2375 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2387 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2399 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2411 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2423 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2429 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2431 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2443 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2455 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2467 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2479 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2485 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2487 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2499 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2511 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2523 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2535 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2541 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2543 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2555 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2567 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2579 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2591 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2597 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2599 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2611 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2623 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2635 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2647 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2653 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2655 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2667 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2679 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2691 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3082 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3094 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3106 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3108 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3120 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3132 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3144 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3156 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3162 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3164 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3176 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3188 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3200 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3212 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3218 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3220 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3232 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3244 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3256 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3268 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3274 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3276 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3288 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3300 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3312 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3324 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3330 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3332 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3337 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3349 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3373 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3388 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3400 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3412 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3424 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3436 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3442 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3444 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3456 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3468 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3480 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3492 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3498 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3500 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3512 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3524 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3536 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3548 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3554 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3556 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3568 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3580 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3592 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3604 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3610 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3612 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3624 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3636 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3648 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3660 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3666 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3668 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3680 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3692 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3704 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3716 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3722 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_3724 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_3732 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3739 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3751 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3763 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3775 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3780 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3792 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3804 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3816 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3828 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3834 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3836 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3848 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3860 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3872 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3884 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3890 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3892 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3898 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3902 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3906 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3910 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3914 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3918 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3922 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3926 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3930 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3934 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3938 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3943 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3948 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3952 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3956 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3960 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3964 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3968 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3972 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3976 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3980 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3984 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3996 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4002 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4004 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4016 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_4028 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_4036 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_4040 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4044 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_4056 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4060 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_4072 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_4080 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4085 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4097 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4103 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_4106 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_4113 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_4116 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_4122 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_4126 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_4130 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_4134 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_4138 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_4142 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_4146 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_4151 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_4155 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_4159 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_4163 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_4167 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_4172 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4176 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4188 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4200 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4212 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_4217 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_4225 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4228 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_4240 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4248 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_4253 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_4261 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4269 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_4281 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4284 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4296 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4308 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4320 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4332 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4338 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4340 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4352 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4364 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4376 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4388 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4394 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4396 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4408 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4420 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4432 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4444 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4450 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4452 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4464 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4476 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4488 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4500 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4506 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4508 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4520 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4532 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4544 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4556 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4562 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_4564 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_4579 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1039 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1059 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1095 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1151 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1207 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1263 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1283 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1295 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1307 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1319 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1339 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1351 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1375 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1387 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1395 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1407 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1419 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1431 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1443 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1449 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1451 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1493 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1507 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1519 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1527 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1531 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1535 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1549 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1553 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1557 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1563 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1575 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1587 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1599 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1611 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1617 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1619 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1627 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1631 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1635 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1639 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1643 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1647 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1659 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1671 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1675 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1687 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1699 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1711 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1723 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1729 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1731 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1743 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1755 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1759 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1762 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1766 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1770 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1774 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1778 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1787 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1799 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1811 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1817 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1820 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1828 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1832 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1843 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1855 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1859 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1862 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1874 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1886 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1899 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1911 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1923 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1935 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1947 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1953 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1955 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1967 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1975 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1978 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1982 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1986 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1990 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1994 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1998 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_2002 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_2006 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_2011 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2027 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2039 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2042 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2054 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2067 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_2072 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2076 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2088 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2100 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2106 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_2111 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2119 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2123 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2135 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2147 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2159 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2171 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2177 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2179 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2191 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2203 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2215 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2227 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2233 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2235 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2247 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2251 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2255 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2267 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_2279 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2287 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2291 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2303 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2315 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2327 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2339 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2345 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2347 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2359 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2371 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2383 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2395 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2401 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2403 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2422 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_2434 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_2444 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2459 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_2471 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2479 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_2484 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2490 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2502 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2515 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2527 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2539 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2551 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2563 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2569 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2571 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2583 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_2595 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_2599 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2604 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_2616 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_2624 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2627 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2639 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2651 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2663 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2675 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2681 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_2683 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_2688 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2692 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2704 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3082 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3094 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3106 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3118 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3130 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3134 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3136 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3148 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3160 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3172 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3184 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3190 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3192 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3204 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3208 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3211 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3215 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3227 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_3239 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3248 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3260 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3272 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3284 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3296 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3301 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3304 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3310 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3314 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3326 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3338 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_3350 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3358 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3360 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3367 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3379 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3403 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3416 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3428 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3440 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3445 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3451 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3455 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3467 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3472 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3484 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3496 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3508 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3520 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3526 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3528 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3540 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3552 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3564 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3576 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3582 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3584 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3596 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3608 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3620 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3632 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3638 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3640 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3652 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3664 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3676 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3688 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3694 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3696 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3708 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3720 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3732 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3744 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3750 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3752 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3764 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3776 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3788 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3800 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3806 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3808 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3820 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3832 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3844 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3856 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3862 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3864 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3876 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3888 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3900 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3912 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3918 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_3920 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3928 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3933 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3945 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_3957 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_3967 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3976 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3988 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3993 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3997 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4001 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4005 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4009 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4013 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4018 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4022 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4026 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_4032 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_4036 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4039 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4043 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4047 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4051 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4055 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4059 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4063 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4067 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4071 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4075 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4079 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4084 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4088 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4092 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4096 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4100 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4104 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4108 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4112 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4116 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4120 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4127 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4131 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4135 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4139 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4144 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4148 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4152 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4164 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4176 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_4188 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4196 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4200 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4212 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4224 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4236 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_4248 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_4254 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4256 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_4262 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4270 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4282 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4294 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_4306 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_4310 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4312 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4324 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4336 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4348 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_4360 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_4366 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4368 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4380 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4392 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4404 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_4416 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_4422 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4424 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4436 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4448 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4460 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_4472 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_4478 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4480 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4492 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4504 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4516 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_4528 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_4534 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4536 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4548 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4560 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4572 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4577 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1011 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1067 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1084 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1120 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1179 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1235 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1267 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1279 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1291 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1323 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1335 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1347 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1365 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1367 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1389 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1401 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1423 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1435 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1447 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1459 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1471 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1479 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1491 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1499 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1511 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1521 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1525 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1529 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1533 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1535 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1539 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1543 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1547 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1551 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1555 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1559 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1563 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1567 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1571 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1577 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1581 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1585 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1589 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1591 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1596 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1608 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1618 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1622 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1626 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1630 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1643 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1647 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1651 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1655 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1659 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1663 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1671 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1683 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1687 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1691 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1699 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1703 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1707 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1710 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1715 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1719 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1723 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1735 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1743 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1750 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1754 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1759 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1763 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1766 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1770 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1774 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1778 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1789 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1801 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1805 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1808 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1815 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1820 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1825 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1832 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1836 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1840 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1844 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1850 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1854 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1858 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1867 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1871 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1883 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1906 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1918 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1927 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1939 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1951 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1963 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1969 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1974 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1978 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1983 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1987 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1990 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1994 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1998 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_2002 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2006 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_2012 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2020 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_2034 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_2039 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_2043 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_2047 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_2051 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2059 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_2062 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_2070 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_2074 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_2078 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2082 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2095 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2107 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2119 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2131 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2143 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2149 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2151 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2163 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2175 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2187 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2199 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2207 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2219 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2231 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2243 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2255 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2261 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2263 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2275 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2287 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2299 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2311 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2317 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2319 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2331 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2343 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2355 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2367 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2373 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2375 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2387 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2399 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2411 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2423 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2429 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_2431 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_2439 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2457 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2469 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2481 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2485 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2487 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2499 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_2511 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2521 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_2533 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2541 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2543 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_2555 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2564 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2576 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_2587 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_2595 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2599 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2611 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2623 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2635 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2647 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2653 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2655 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2667 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2679 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2691 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3082 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3094 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3106 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3108 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3120 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3132 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3144 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_3156 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3161 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3164 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3176 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3180 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3192 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3204 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_3216 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3220 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3232 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3244 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3256 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3268 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3274 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3276 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3288 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3300 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3312 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3324 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3330 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3332 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3344 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3356 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3368 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3380 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3386 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3388 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_3400 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3408 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3412 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3424 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3436 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3442 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3444 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3456 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3468 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3472 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3482 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3494 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3498 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3500 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3512 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3524 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3536 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3548 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3554 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3556 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3568 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3580 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3592 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3597 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3609 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3612 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3623 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3635 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3647 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_3659 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3668 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3674 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3686 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3690 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3694 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3706 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3718 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3722 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3724 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3736 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3748 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3760 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3772 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3778 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3780 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3792 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3804 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3816 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3828 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3834 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3836 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3848 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3860 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3872 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3884 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3890 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3892 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3904 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3916 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3928 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3940 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3946 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3948 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3960 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3972 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3984 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3996 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_4002 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4004 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_4016 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4020 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_4032 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_4038 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_4041 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_4045 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_4049 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_4053 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_4057 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_4060 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_4066 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_4070 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_4074 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_4078 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_4082 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_4087 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_4091 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_4095 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_4099 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_4103 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_4107 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_4111 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_4116 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_4121 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_4125 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_4129 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_4133 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_4137 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_4141 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_4145 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_4149 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4153 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_4165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4172 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4184 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4196 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4208 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_4220 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_4226 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4228 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4240 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_4252 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4260 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_4272 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_4280 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4284 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4296 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4308 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4320 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_4332 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_4338 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4340 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4352 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4364 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4376 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_4388 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_4394 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4396 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4408 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4420 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4432 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_4444 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_4450 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4452 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4464 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4476 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4488 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_4500 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_4506 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4508 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4520 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_4532 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_4540 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_4545 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_4549 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_4553 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_4557 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_4561 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_4564 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_4579 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1022 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1127 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1155 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1183 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1211 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1239 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1251 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1283 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1295 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1307 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1323 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1339 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1351 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1367 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1379 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1395 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1407 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1419 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1423 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1435 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1447 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1451 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1463 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1475 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1479 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1487 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1499 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1505 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1507 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1511 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1514 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1518 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1522 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1526 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1530 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1535 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1539 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1543 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1547 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1551 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1555 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1559 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1563 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1572 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1576 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1580 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1584 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1588 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1591 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1603 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1606 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1610 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1614 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1619 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1623 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1627 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1631 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1635 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1639 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1643 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1647 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1651 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1655 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1658 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1664 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1672 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1675 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1683 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1688 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1703 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1708 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1716 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1721 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1725 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1729 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1731 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1740 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1744 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1750 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1754 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1759 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1764 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1772 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1778 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1784 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1787 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1791 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1795 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1803 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1806 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1810 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1815 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1824 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1828 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1832 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1836 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1843 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1849 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1853 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1864 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1868 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1871 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1880 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1892 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1899 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1907 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1916 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1922 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1927 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1939 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1951 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1955 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1961 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1972 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1978 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1983 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1987 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1990 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1994 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1998 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2002 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2006 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2011 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2015 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2019 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2023 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2027 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2030 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2034 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2039 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2043 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2047 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2051 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2055 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2058 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2062 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2067 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2071 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2075 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2079 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2083 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2092 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2095 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2099 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2103 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2107 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_2119 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2123 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2135 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_2147 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2151 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2163 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_2175 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2179 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2188 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2200 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2207 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2219 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_2231 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2235 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2247 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_2259 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2263 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2275 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_2287 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2291 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2303 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_2315 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2319 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2331 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_2343 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2347 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2359 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_2371 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2375 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2387 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_2399 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2403 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2409 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_2421 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2429 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2431 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2443 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_2455 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2459 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2471 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_2483 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2487 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2499 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_2511 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2515 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2527 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_2539 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2543 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2555 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_2567 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2571 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2583 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_2595 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2599 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2611 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_2623 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2627 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2639 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_2651 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2655 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2667 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_2679 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2683 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_2695 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3082 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3094 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3106 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3108 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3120 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3132 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_3136 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3144 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3149 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3164 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3176 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3188 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3192 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3211 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3215 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3220 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3224 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_3236 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3244 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3248 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3260 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3272 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3276 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3288 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_3292 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3300 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3304 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3316 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3328 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3332 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3344 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3356 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_3360 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3368 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3371 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_3383 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3388 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3400 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3412 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3416 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3428 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3440 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3444 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3456 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3468 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3472 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3484 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3496 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_3500 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3508 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_3518 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3526 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3528 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_3540 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3548 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3553 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3556 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3568 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3572 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_3576 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3582 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_3584 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3592 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3596 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3608 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3612 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3624 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3636 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3640 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3652 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3664 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3668 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3680 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3692 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3696 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3708 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3720 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3724 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3736 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3748 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3752 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3764 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3776 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3780 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3792 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3804 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3808 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3820 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3832 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3836 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3848 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3860 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3864 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3876 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3888 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3892 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3904 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3916 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3920 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3932 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3944 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3948 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3960 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3972 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3976 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3988 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_4000 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4004 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4016 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_4028 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4032 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4044 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_4056 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4060 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4072 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_4084 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4088 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4100 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_4112 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_4116 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4120 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_4132 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_4140 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4144 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4156 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_4168 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4172 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4184 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_4196 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4200 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4212 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_4224 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4228 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4240 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_4252 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_4256 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_4262 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4267 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_4279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4284 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4296 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_4308 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_4312 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4317 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_4329 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_4337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4340 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4352 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_4364 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4368 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4380 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_4392 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4396 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4408 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_4420 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4424 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4436 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_4448 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4452 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4464 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_4476 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4480 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4492 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_4504 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4508 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4520 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_4532 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4536 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4548 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_4560 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_4564 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_4572 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_4577 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_972 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1123 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1179 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1235 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1267 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1279 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1291 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1323 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1335 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1347 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1367 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1379 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1391 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1403 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1423 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1435 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2249 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2273 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2275 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2287 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2299 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2311 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2323 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2329 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2331 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2343 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2355 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2367 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2379 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2385 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_2387 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_2395 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2419 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_2431 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_2439 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2443 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2455 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2467 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2483 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_2495 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2499 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2511 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2523 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2535 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2547 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2553 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_2555 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_2563 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2572 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2584 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2596 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_2608 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2611 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2623 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2635 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2647 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2659 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2665 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2667 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2679 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2691 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3082 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3094 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3097 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3101 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3105 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3108 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3112 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3116 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3120 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3129 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3133 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3137 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3141 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3145 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3149 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3153 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3157 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3161 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3164 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3176 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3180 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3184 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3188 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3192 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3196 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3208 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3212 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_3216 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3220 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3224 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3228 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3232 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3236 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3240 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3244 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3248 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3260 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_3272 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3276 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3288 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3300 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3304 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3319 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3332 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3344 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3356 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3368 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3380 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3386 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3388 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3400 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3412 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3424 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3436 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3442 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3444 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3456 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3468 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3471 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3483 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3495 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3500 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_3512 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3517 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3521 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3525 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3529 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3533 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3537 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3541 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3545 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3549 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3553 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3556 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3568 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3572 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3576 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3580 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3584 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3588 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3592 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3596 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3600 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3604 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_3608 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3612 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3616 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_3628 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_3636 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3655 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3661 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_3664 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3668 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3680 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3692 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3704 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3716 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3722 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3724 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3736 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3748 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3760 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3772 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3778 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3780 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3792 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3804 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3816 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3828 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3834 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3836 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3848 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3860 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3872 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3889 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_3892 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3900 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3903 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3907 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3919 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3925 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3937 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3941 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3948 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3960 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3972 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3984 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3996 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_4002 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4004 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4022 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4034 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4046 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_4058 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4060 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4072 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4084 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4096 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_4108 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_4114 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4116 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4130 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4134 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4138 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4142 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4146 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4150 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4155 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4159 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4163 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_4167 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4172 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4176 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4180 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4192 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4204 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_4216 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_4222 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4225 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_4228 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_4232 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4235 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4239 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4243 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4247 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4254 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4258 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4262 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4266 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4270 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4274 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_4278 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_4282 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4284 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4291 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4295 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4299 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4303 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4307 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4311 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4315 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4319 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4323 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_4335 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4340 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4352 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4364 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4376 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_4388 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_4394 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4396 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4408 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4420 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4432 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_4444 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_4450 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4452 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4464 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4476 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4488 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_4500 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_4506 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4508 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4520 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4532 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4544 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_4556 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_4562 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4564 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_4576 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_4580 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1008 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1095 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1207 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1263 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1283 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1295 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1307 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1319 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1339 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1357 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1368 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1372 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1384 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1392 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1395 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1413 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1416 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1428 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1436 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2261 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2273 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2285 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2297 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2301 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2303 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2315 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2327 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2339 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_2351 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2357 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2359 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2371 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_2383 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_2391 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_2395 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_2407 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2413 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2415 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2427 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2432 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2444 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2456 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_2468 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2471 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2483 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2495 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2507 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_2519 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2525 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_2527 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2539 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2551 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2563 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_2575 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2581 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2583 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2595 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2607 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2619 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_2631 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2637 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2639 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2651 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2663 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2675 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_2687 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2693 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_2695 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3082 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3094 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3098 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3110 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3122 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3134 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3136 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3148 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3160 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3172 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_3184 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3190 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_3192 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3200 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3203 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3212 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3216 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3220 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3232 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3244 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3248 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3260 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_3272 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3278 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3290 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3302 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3304 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3316 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3328 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3340 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_3352 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3358 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3360 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3372 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3384 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3396 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_3408 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3414 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3416 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3428 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3440 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3452 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_3464 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3470 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3472 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3484 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3496 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3508 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_3520 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3526 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3528 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3537 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3541 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3565 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_3577 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3584 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3596 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3608 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_3620 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3626 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3640 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3652 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3656 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3660 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3664 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3668 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3677 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3681 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3685 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_3689 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3696 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3714 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3726 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3738 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3750 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3752 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3764 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3776 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3788 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_3800 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3806 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3808 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3820 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_3832 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3840 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3845 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3849 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3853 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3857 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3861 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3864 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3877 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3891 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3895 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3899 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3903 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3907 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3911 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3915 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3920 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3932 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3944 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3956 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_3968 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3974 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3976 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3988 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4000 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4012 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_4024 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_4030 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4032 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_4044 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_4050 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_4053 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_4057 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_4061 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_4065 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_4069 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_4073 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_4085 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_4088 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_4092 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_4096 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_4100 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_4104 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4117 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4129 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_4141 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4144 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4156 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4168 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4180 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_4192 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_4198 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4200 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4212 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4224 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4236 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_4248 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_4254 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_4256 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_4262 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4267 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4291 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_4303 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_4312 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_4317 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_4321 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_4325 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_4329 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_4333 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_4337 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_4349 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_4353 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_4357 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_4361 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_4365 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4368 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4380 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4392 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4404 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_4416 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_4422 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4424 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4436 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4448 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4460 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_4476 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4480 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4492 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4504 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4516 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_4528 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_4534 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4536 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4548 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_4560 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_4566 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_4579 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1011 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1031 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1051 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1127 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1179 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1235 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1253 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1263 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1274 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1298 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1323 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1335 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1347 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1365 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1367 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_1375 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1380 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1392 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1404 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1416 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1423 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_1435 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2249 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2273 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2275 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2287 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2299 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2311 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_2323 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2329 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2331 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2343 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2355 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2367 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_2379 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2385 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_2387 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2395 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_2398 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_2410 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_2424 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2428 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_2440 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2443 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2455 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2467 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2479 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_2491 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2497 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2499 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2511 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2523 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2535 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_2547 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2553 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_2555 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2564 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2576 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2588 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_2600 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_2608 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2611 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2623 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2635 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2647 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_2659 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2665 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2667 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_2679 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_2687 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_2691 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_2703 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3082 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3087 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_3099 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3108 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3120 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3132 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3144 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_3156 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_3162 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3164 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3176 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3188 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3200 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_3209 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3220 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3232 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3244 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3256 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_3268 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_3274 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3276 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3288 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3300 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3312 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_3323 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3332 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3344 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3356 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3368 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_3380 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_3386 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3388 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3400 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3412 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3424 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_3436 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_3442 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3444 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3456 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3468 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3480 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_3492 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_3498 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3500 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3512 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3524 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3536 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_3548 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_3554 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3556 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3562 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3566 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3570 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3579 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3583 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3587 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3591 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3597 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3601 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3605 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3609 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_3612 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3617 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3621 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3625 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3629 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3641 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3652 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3656 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3660 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_3664 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3668 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3672 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_3676 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3679 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3683 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3687 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3691 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3695 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3699 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3703 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3707 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3719 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3724 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3728 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3740 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3752 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3764 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_3776 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3780 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3792 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3796 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3800 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3804 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3816 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_3828 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_3834 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3836 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_3848 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_3856 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3861 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3873 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_3885 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_3892 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3911 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3923 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3935 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3948 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3960 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3972 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3984 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_3996 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_4002 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_4004 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_4016 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_4028 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_4036 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_4048 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_4056 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_4060 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_4072 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_4084 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_4096 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_4108 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_4114 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_4116 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_4128 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_4142 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_4146 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_4155 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_4159 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_4172 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_4184 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_4196 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_4208 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_4220 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_4226 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_4228 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_4240 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_4252 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_4264 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_4276 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_4282 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_4284 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_4296 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_4308 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_4316 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_4321 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_4325 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_4329 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_4333 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_4337 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_4340 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_4352 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_4356 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_4360 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_4364 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_4368 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_4372 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_4384 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_4392 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_4396 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_4408 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_4420 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_4432 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_4444 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_4450 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_4452 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_4464 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_4476 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_4488 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_4500 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_4506 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_4508 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_4520 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_4532 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_4544 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_4556 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_4562 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_4564 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_4572 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_4577 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1027 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1039 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1139 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1151 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1171 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1207 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1225 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1235 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1238 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1266 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1278 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1283 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1291 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1296 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1304 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1325 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1337 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1339 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1351 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1375 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1387 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1393 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1395 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1407 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1419 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1431 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1437 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2261 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2273 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2285 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2297 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2301 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2303 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2315 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2327 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2339 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_2351 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2357 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2359 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2371 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_2374 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_2383 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2392 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_2404 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_2412 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2415 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2427 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_2430 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2439 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2451 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_2463 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2469 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_2471 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_2480 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2487 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2499 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2511 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_2523 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_2527 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2536 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2563 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_2575 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2581 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2583 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2595 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2607 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2619 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_2631 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2637 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2639 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2651 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2663 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_2675 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_2687 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2693 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_2695 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_2703 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3082 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3094 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3098 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_3110 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_3118 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_3128 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_3134 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3136 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3148 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3160 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_3172 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_3180 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3185 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3189 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3192 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3201 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3205 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3216 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_3220 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3228 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_3240 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_3246 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3248 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3257 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3269 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3281 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_3293 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3301 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3304 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3319 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3331 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3343 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3355 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3360 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_3372 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_3378 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3382 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3394 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_3406 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_3414 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3416 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3428 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3440 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3452 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3464 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3472 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3484 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3496 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3508 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_3520 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_3526 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3528 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3540 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3552 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3564 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_3576 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_3582 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_3584 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3589 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3593 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3597 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3601 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3605 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3609 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3613 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3617 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3626 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3630 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3634 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_3638 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3640 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3644 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3648 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3652 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3656 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3660 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_3664 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_3667 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_3673 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3676 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_3680 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3691 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3696 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3700 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_3704 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3707 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3711 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3720 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3724 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_3733 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3741 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3745 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3749 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3752 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3756 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3760 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3764 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3776 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3780 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3784 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3788 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3792 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3798 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3808 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3820 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3832 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3844 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_3856 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_3862 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3864 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3876 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3888 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3900 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_3912 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_3918 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_3920 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_3928 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3933 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_3937 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3945 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3953 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_3965 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3973 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3976 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3994 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_4006 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_4018 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_4030 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_4032 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_4044 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_4056 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_4068 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_4080 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_4086 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_4088 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4096 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4100 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4104 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4108 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4112 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4116 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4120 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4129 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4133 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4137 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4141 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4144 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4148 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4152 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_4156 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_4168 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_4180 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_4192 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_4198 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_4200 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_4212 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_4224 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_4232 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4237 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4241 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4245 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4249 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4253 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4256 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4265 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4269 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4273 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4277 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4281 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4285 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4289 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_4293 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_4305 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4312 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4324 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_4328 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_4340 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_4352 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_4364 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_4368 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_4380 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_4392 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_4404 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_4416 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_4422 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_4424 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_4436 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_4448 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_4460 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_4472 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_4478 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_4480 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_4492 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_4504 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_4516 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_4528 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_4534 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_4536 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_4542 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4545 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4549 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4553 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4557 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4561 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4565 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4579 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1011 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1067 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1085 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1112 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1132 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1212 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1216 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1252 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1255 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1270 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1282 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1290 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1294 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1298 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1302 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1323 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1335 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1347 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1365 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1367 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1379 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1391 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1403 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1435 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2249 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_2269 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2272 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2275 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2284 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2288 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2300 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2312 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_2324 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2331 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2343 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2355 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2367 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_2379 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_2385 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2387 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_2396 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2408 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2420 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_2426 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_2430 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_2435 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_2441 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2443 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2456 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_2468 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2471 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_2480 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2491 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_2495 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2499 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2511 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2523 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2535 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_2547 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_2553 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2555 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2567 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2579 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2591 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_2603 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_2609 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2611 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2623 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2635 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_2647 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_2655 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2660 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2664 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_2667 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2681 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2685 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2689 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2693 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_2697 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3082 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3094 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_3106 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3108 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3120 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3132 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3144 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_3156 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_3162 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3164 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3176 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3188 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3200 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_3212 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_3218 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_3220 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_3228 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3236 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3248 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3260 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_3272 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_3276 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_3282 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3290 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3298 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3310 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_3322 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_3330 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3332 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_3344 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3353 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3360 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3372 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_3384 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_3388 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3398 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3410 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3422 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_3434 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_3442 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3444 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3448 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_3460 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3465 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3477 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_3489 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3497 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3500 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3512 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3524 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3536 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_3548 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_3554 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3556 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3568 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3580 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3592 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_3604 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_3610 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3612 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_3624 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_3632 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3635 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3647 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_3659 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3668 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_3680 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_3688 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3691 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3695 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3699 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3703 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3707 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3711 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_3720 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3724 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3735 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3739 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3743 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_3747 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3750 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3754 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3758 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3762 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3774 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_3778 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3780 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_3792 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3821 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3836 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3848 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3860 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3872 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_3884 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3889 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3892 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_3896 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3899 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3903 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3907 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3911 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3923 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3927 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_3931 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3941 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3945 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_3948 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3953 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3957 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_3969 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_3977 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_3980 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3988 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3992 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4001 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4004 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_4008 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4018 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_4022 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_4034 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_4046 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_4058 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_4060 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_4072 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_4084 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_4092 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4097 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4101 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4105 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4109 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4113 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_4116 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_4120 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4128 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4132 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4136 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4140 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4144 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4148 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4152 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_4156 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_4162 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4165 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4169 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4172 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4181 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4185 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4189 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_4193 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_4205 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_4217 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4225 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_4228 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4236 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4240 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4244 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4256 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_4260 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_4272 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_4280 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_4284 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_4296 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_4308 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_4320 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_4332 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_4338 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_4340 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_4352 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_4364 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_4376 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_4388 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_4394 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_4396 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_4408 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_4420 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_4432 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_4444 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_4450 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_4452 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_4460 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4465 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4469 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4473 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4477 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4486 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4490 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4494 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_4498 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_4506 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_4508 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_4520 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_4532 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_4544 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_4556 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_4562 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_4564 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_4572 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4577 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_984 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1039 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1095 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1127 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1207 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1225 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1235 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1238 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1266 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1278 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1283 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1291 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1296 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1320 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1332 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1339 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1351 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1375 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1387 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1393 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1395 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1407 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1419 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1431 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1437 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2249 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_2261 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2270 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2282 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_2294 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2303 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2315 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2327 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2339 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_2351 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_2357 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2359 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2371 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_2383 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_2389 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2393 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_2405 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_2413 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2415 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2427 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2439 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_2451 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_2459 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_2464 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_2471 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_2479 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_2485 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2498 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2510 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_2522 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2527 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2539 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2551 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2563 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_2575 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_2581 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2583 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2595 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2607 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2619 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_2631 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_2637 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2639 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2651 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2663 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_2675 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_2687 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_2693 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3082 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3094 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3106 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3118 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3130 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3134 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3136 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3148 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3160 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3172 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3184 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3190 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3192 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3204 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3208 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3216 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3228 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3240 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3246 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3248 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3260 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3272 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_3284 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3289 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3293 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3297 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3301 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3304 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3315 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3319 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3323 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3327 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3331 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3335 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3343 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3355 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3360 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3372 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3376 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3380 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3384 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3388 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3392 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3396 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3407 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3411 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3416 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3420 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3424 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3428 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3434 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_3441 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3448 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3452 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3456 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3460 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_3464 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3469 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3472 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3476 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3488 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3500 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3512 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_3524 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3528 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3540 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3552 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3564 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3576 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3582 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3584 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3596 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3608 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3620 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3626 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3629 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3633 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3637 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3640 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3644 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3648 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3657 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3661 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3665 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3669 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3673 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3677 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3681 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3718 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3730 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3742 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3746 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3750 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3752 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_3764 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_3772 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3777 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3781 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3785 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3789 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3793 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3802 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3806 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3808 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3812 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3816 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3820 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3824 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3836 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3842 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3845 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3849 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3853 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3857 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3861 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3864 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3873 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3877 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3881 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3885 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3889 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3893 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_3897 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3907 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3911 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3915 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3920 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3924 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3928 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3948 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3952 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3958 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3961 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3965 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3969 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3973 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3976 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3980 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3992 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_4003 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_4007 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_4011 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_4015 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_4019 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_4022 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_4026 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_4030 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_4032 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_4044 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_4056 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_4068 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_4080 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_4086 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_4088 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_4098 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_4102 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_4114 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_4118 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_4130 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_4142 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_4144 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_4156 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_4168 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_4180 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_4192 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_4198 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_4200 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_4212 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_4224 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_4236 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_4248 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_4254 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_4256 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_4266 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_4270 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_4274 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_4278 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_4282 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_4286 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_4295 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_4299 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_4303 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_4307 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_4312 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_4316 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_4320 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_4332 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_4344 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_4356 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_4364 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_4368 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_4380 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_4392 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_4404 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_4416 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_4422 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_4424 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_4436 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_4448 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_4460 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_4472 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_4478 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_4480 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_4492 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_4504 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_4516 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_4528 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_4534 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_4536 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_4548 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_4560 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_4566 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_4579 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_975 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1001 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1123 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1267 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1279 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1291 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1323 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1334 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1346 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1358 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1367 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1381 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1409 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1423 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1435 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2249 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_2273 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2275 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2287 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2299 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2311 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_2323 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_2329 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2331 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2343 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2355 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2367 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_2379 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_2385 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_2387 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_2395 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2417 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_2441 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2443 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2455 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2467 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_2473 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2482 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2494 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_2507 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2515 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2527 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2539 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_2551 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2555 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2567 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_2579 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_2589 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_2593 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2605 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_2609 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2611 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2623 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2635 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_2647 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_2650 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2662 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_2667 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_2679 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_2683 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_2687 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_2691 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3082 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3094 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_3106 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3108 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3120 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3132 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3144 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3156 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_3162 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3164 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3176 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3188 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3200 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3212 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_3218 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3220 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3232 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3244 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3256 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3268 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_3274 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3276 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3288 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3300 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3312 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3324 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_3330 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_3332 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3340 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3344 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3348 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3352 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3356 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3360 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_3372 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3377 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3381 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3385 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_3388 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3393 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3397 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3401 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3405 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3409 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3413 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3417 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3421 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3433 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3437 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3441 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3444 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3448 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3452 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_3456 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3466 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3470 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3474 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3478 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3482 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3488 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3492 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_3496 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3500 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3504 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3508 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3512 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3516 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3520 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3524 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3535 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_3547 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3556 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3568 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3580 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3592 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3604 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_3610 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3612 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_3624 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_3632 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3649 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3661 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3668 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_3680 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3690 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3694 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3698 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3702 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_3706 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3709 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3718 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_3722 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3724 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3728 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3732 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3736 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3740 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3744 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3748 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3752 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3764 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_3776 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3780 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3792 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3804 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3816 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3828 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_3834 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3836 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3848 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3860 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3872 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3884 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_3890 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3892 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_3896 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3899 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_3911 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_3919 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3924 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3928 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3937 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3941 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3948 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3960 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3972 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3984 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3996 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_4002 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_4004 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4018 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_4022 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_4030 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_4036 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_4043 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_4050 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_4058 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_4060 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_4072 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_4084 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_4092 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_4097 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_4109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_4116 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_4128 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_4140 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_4152 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_4164 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_4170 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_4172 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_4180 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4183 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4192 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_4196 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_4208 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_4218 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_4226 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_4228 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_4240 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_4252 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_4264 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_4276 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_4282 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_4284 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4292 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_4310 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_4318 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4321 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4325 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4329 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4333 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4337 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4340 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4349 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4353 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4357 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4361 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_4369 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_4381 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4393 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_4396 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_4408 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_4420 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_4432 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_4444 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_4450 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_4452 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4458 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4462 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4466 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4470 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4474 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4478 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4487 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4491 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4495 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4499 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_4503 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4508 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_4512 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_4524 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_4536 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_4548 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_4560 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_4564 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_4576 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_4580 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1425 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1437 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2249 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_2273 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2275 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2287 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_2299 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2303 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_2315 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_2318 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_2327 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_2331 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_2343 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_2347 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_2355 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2359 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2371 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_2383 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2387 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2399 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_2411 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_2415 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_2424 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2428 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_2440 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_2443 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_2452 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_2463 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_2469 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2471 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2483 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_2495 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2499 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2511 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_2523 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2527 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2539 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_2551 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2555 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2567 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_2579 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_2583 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_2591 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_2596 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_2608 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2611 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2623 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_2635 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2639 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2651 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_2663 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2667 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2679 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_2691 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_2695 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3082 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3094 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_3106 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3108 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3120 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3132 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3136 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_3148 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3156 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3161 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3164 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3173 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3177 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3192 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_3204 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3212 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3217 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3220 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3229 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3233 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3245 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_3248 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_3256 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3261 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3273 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3276 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3288 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3300 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3304 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3313 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_3325 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_3332 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3340 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3344 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3348 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3352 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3356 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3360 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3364 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3368 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3372 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_3376 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3384 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3388 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3392 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3404 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3412 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3416 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3421 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3425 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3429 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3433 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3437 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3441 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3444 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3448 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3452 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3456 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3465 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3469 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3472 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3476 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3490 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3494 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_3498 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3500 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3504 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_3518 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_3526 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_3528 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_3534 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3537 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3541 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3545 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3549 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3553 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3556 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3567 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3571 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3575 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3579 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3584 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3588 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_3600 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3608 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3612 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3624 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3636 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_3640 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_3648 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3665 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3668 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3673 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3677 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3681 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3685 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3689 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3693 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3696 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3705 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3709 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3713 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3717 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3721 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3724 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3728 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3732 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_3744 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_3750 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3752 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3764 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3776 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3780 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3792 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3804 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3808 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3820 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3832 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3836 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3848 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3860 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3864 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3876 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3888 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3892 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3904 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3916 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_3920 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3928 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3933 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3948 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3960 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3972 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3976 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_3996 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_4002 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_4004 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_4016 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_4028 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_4032 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_4040 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4045 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4049 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4053 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4057 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_4060 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4066 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4071 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4075 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4079 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_4083 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4088 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4092 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_4096 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4101 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4105 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4109 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4113 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4116 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4121 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4125 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4129 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4133 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4137 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4141 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4144 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4148 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_4152 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_4164 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_4170 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_4172 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_4184 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_4196 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_4200 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_4212 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_4224 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_4228 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_4240 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_4252 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_4256 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_4268 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_4280 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_4284 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_4296 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_4308 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_4312 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4324 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4333 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4337 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4340 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_4347 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4356 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_4360 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_4366 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_4368 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_4380 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_4383 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_4396 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_4408 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_4420 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_4424 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_4436 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_4448 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_4452 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_4458 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4461 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4465 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4469 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4473 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4477 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4480 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4489 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4493 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4497 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4501 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4505 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4508 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4512 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4516 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_4520 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_4532 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_4536 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_4548 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_4560 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_4564 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_4576 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_4580 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1179 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1248 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1397 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1409 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1414 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1426 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1435 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2249 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_2273 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2275 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2287 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2299 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2311 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_2323 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_2329 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2331 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2343 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2355 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2367 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_2379 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_2385 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2387 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2399 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2411 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2423 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_2435 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_2441 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_2443 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2476 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_2488 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_2496 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_2499 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_2508 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_2512 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_2522 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2531 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_2543 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_2551 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2555 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_2567 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_2571 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2579 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2591 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_2603 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_2609 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2611 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_2623 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_2631 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_2635 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2644 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_2656 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_2664 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2667 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2679 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2691 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3082 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3094 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_3106 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3108 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3120 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3132 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_3144 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_3150 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3153 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3157 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3161 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3164 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3173 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3177 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3181 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3185 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3197 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_3209 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3220 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3232 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3244 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3256 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_3268 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_3274 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3276 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_3288 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_3296 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3301 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3305 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3309 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3313 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3317 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3321 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3325 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3329 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3332 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3344 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3348 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_3352 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3355 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3359 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3363 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3367 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3376 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_3380 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_3386 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3388 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_3400 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3408 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_3417 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3432 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3436 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_3440 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3444 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3453 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3457 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3461 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3465 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3469 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3476 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_3488 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_3494 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3497 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_3500 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3505 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3509 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3513 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3517 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3526 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3530 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_3534 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3537 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3541 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3545 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3549 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3553 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3556 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3568 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3572 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3576 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3580 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3584 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3588 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3592 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_3604 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_3610 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3612 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3621 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3625 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3649 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_3661 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_3668 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_3676 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_3686 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3694 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3703 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3715 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3719 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3724 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3728 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3740 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3752 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3764 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_3776 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3780 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3792 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3804 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3816 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_3828 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_3834 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3836 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3848 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_3860 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3877 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3889 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3892 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3904 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3916 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3928 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_3940 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_3946 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3948 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_3960 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3979 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3999 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_4004 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_4016 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_4028 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_4040 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_4052 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_4058 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_4060 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_4072 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_4084 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_4096 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_4108 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_4114 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_4116 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_4124 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4129 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4133 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4137 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4141 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4145 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4149 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4154 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4158 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4162 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_4166 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_4170 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4172 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4176 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_4180 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_4192 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_4204 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_4216 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_4224 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_4228 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_4240 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_4252 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_4264 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_4276 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_4282 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_4284 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_4296 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_4308 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_4320 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_4332 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_4338 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_4340 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_4352 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_4358 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_4370 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_4374 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4377 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4381 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4385 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4389 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4393 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_4396 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4401 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4410 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4414 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4418 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4422 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4426 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4430 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4434 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_4438 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_4450 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_4452 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4457 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4461 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4465 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4469 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4473 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4477 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4486 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4490 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4494 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4498 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_4502 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_4506 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4508 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_4512 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_4524 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_4536 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_4548 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_4560 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_4564 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_4576 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_4580 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1425 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1436 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_2249 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2257 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2281 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_2293 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_2301 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2303 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2315 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2327 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2339 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_2351 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_2357 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_2359 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2368 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2380 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2392 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_2404 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_2412 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2415 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2427 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2441 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2453 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2465 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_2469 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_2471 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2484 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2496 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2508 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_2520 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2527 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2539 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_2551 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_2555 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2563 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_2573 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_2581 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2583 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2595 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2607 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2619 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_2631 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_2637 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2639 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2651 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2663 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_2675 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_2683 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_2692 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_2695 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_2703 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3082 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3094 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3106 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3118 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3130 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_3134 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3136 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3148 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3160 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3172 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_3184 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_3190 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3192 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3204 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3216 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3228 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_3240 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_3246 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3248 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3260 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3272 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3284 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_3296 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_3302 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_3304 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3314 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3318 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3322 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3326 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3335 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3339 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3343 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3347 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3353 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3357 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3360 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3364 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3368 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3372 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3376 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3387 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_3391 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3399 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3410 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_3414 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3416 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3420 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3424 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3428 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3432 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3444 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3456 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_3468 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3472 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3484 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3496 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_3508 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_3514 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_3517 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3528 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_3540 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3548 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3552 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3564 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_3576 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_3582 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3584 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3602 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3614 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3626 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_3630 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3633 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3637 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3640 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3652 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3656 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3660 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3672 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_3684 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_3692 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3696 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3708 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3720 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3732 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_3744 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_3750 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3752 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3764 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3776 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3788 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_3800 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_3806 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3808 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3820 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3832 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3844 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_3856 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_3862 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3864 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3876 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3888 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3900 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_3912 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_3918 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3920 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3932 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3944 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3956 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_3968 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_3974 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3976 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3994 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_4006 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_4018 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_4030 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_4032 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_4044 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_4056 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_4068 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_4081 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_4088 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_4100 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_4112 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_4124 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_4136 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_4142 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_4144 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_4156 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_4168 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_4180 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_4192 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_4198 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_4200 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_4212 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_4224 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_4231 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_4243 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_4256 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_4268 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_4280 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_4292 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_4304 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_4310 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_4312 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_4324 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_4330 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_4334 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_4338 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_4342 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_4346 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_4350 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_4357 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_4361 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_4365 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_4368 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_4373 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_4380 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_4384 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_4388 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_4392 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_4396 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_4400 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_4404 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_4408 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_4412 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_4420 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_4424 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_4436 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_4448 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_4460 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_4472 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_4478 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_4480 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_4492 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_4504 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_4516 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_4528 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_4534 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_4536 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_4548 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_4560 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_4572 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_4580 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1427 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1434 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_2249 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2253 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_2265 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_2273 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2275 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2287 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2299 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2311 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_2323 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_2329 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2331 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2343 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2355 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2367 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_2379 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_2385 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2387 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2399 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2411 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2423 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_2435 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_2441 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2443 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2455 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2467 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2479 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_2491 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_2497 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2499 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2518 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2530 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2542 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2555 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2567 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2579 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2591 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_2603 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_2609 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2611 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2623 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2635 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2647 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_2659 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_2665 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2667 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2679 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_2691 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_2703 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3082 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3091 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3095 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3108 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3120 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3132 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3144 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_3156 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_3162 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3164 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3176 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_3188 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3201 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_3213 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3220 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3232 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3244 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3256 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_3268 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_3274 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3276 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3288 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3300 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3312 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_3324 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_3330 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_3332 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_3340 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3345 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3349 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3353 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3357 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3361 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3365 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3374 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3378 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_3382 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_3386 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3388 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3392 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_3412 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3420 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3424 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3428 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3432 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3441 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3444 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3448 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3452 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3464 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3476 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_3488 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_3496 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3500 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3512 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3524 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_3536 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3556 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3568 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3580 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3592 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_3604 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_3610 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3612 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3624 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3636 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3648 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_3660 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_3666 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_3668 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_3672 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3675 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3679 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3683 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3687 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3696 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3700 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3704 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3708 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_3712 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_3720 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3724 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3736 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3748 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3760 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_3772 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_3778 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3780 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3792 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3804 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3816 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_3828 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_3834 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3836 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3854 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3866 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3878 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_3890 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3892 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3904 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_3916 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_3922 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_3939 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3948 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3960 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3972 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3984 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_3996 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_4002 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_4004 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_4016 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_4028 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_4040 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_4052 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_4058 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_4060 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_4066 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_4083 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_4095 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_4107 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_4116 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_4128 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_4140 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_4152 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_4164 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_4170 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_4172 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_4184 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_4196 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_4208 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_4220 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_4226 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_4228 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_4240 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_4252 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_4264 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_4276 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_4282 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_4284 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_4296 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_4320 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_4332 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_4338 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_4340 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_4352 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_4364 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_4372 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_4377 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_4381 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_4388 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_4392 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_4396 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_4408 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_4420 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_4432 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_4444 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_4450 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_4452 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_4464 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_4476 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_4488 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_4500 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_4506 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_4508 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_4520 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_4532 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_4544 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_4556 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_4562 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_4564 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_4576 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_4580 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1118 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1301 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1325 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1401 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1426 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1430 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1434 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_2249 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_2255 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2263 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2275 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2287 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_2299 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2303 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_2315 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2326 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2338 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_2350 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2359 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2371 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2383 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_2395 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_2401 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_2404 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_2412 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2415 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2427 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2439 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2451 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_2463 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_2469 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2471 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_2483 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_2497 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_2505 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_2508 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_2517 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_2525 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_2527 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_2572 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_2580 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2583 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_2595 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_2601 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_2604 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_2608 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_2620 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2624 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_2636 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2639 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2651 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2663 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2675 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_2687 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_2693 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_2695 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_2703 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_3082 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_3090 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3095 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3104 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3108 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3120 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_3132 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3136 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3148 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3154 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3166 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3172 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_3181 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3192 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3204 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3216 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3228 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_3240 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_3246 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3248 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3260 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3272 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3284 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_3296 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_3302 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3304 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3316 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_3328 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3357 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3360 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3372 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3384 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_3396 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3416 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3428 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3440 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3452 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_3464 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_3470 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3472 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3484 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3496 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3508 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_3520 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_3526 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3528 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3546 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3558 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3570 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_3582 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3584 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3596 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3608 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3620 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_3632 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_3638 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3640 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3652 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_3664 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_3672 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3682 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_3694 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3696 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3708 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3720 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3732 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_3744 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_3750 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3752 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3773 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3785 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_3797 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3805 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3808 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3820 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3832 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3844 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_3856 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_3862 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3864 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3876 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3888 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3900 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_3912 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_3918 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3920 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3932 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3944 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3956 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_3968 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_3974 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3976 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3988 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4000 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4012 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_4024 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_4030 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4032 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4044 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4056 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_4068 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_4085 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4088 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4100 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4112 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4124 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_4136 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_4142 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4144 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_4156 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4174 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4186 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_4198 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4200 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4212 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4224 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4236 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_4248 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_4254 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4256 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4268 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4280 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4292 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_4304 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_4310 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4312 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_4324 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_4332 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4339 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4351 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_4363 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4368 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_4380 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_4383 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_4389 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4396 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4408 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_4420 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4424 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4436 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4448 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4460 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_4472 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_4478 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4480 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4492 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4504 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4516 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_4528 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_4534 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4536 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4548 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4560 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_4572 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_4580 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1297 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1397 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1401 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1409 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1418 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1434 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2249 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2253 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2257 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_2273 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2275 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2287 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_2299 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2303 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2315 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_2327 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2331 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2343 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_2355 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2359 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2371 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_2383 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2387 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2399 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2403 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2412 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2415 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2427 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_2439 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2443 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2455 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_2467 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2471 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2483 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_2495 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2499 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2511 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_2523 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2527 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2536 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2540 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2552 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2555 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2567 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_2579 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2583 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2595 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_2607 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2611 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2620 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_2632 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2639 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2651 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_2663 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2667 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2671 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2683 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2687 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_2691 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_2695 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2700 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2704 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2708 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2720 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2723 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2735 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2746 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_2751 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2759 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_2770 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2779 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2791 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_2803 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2807 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2819 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2829 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_2833 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_2835 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_2841 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2844 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2848 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2852 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2856 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2860 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2863 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2875 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2885 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_2889 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2891 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2895 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_2907 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_2915 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2919 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2931 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_2943 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2947 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2959 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_2971 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2975 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2979 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2991 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_2995 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_3001 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3003 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3015 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3027 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3031 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3043 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3055 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3059 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3071 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3083 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3087 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3099 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3111 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3115 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3127 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3143 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3155 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3167 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3171 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3183 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3199 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3211 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3223 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3227 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3239 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3251 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3255 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3267 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3279 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_3283 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3291 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3296 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3300 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3304 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3308 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3311 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3320 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3331 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3335 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3339 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3343 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3348 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_3360 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3367 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3379 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3391 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3395 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3407 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3419 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3423 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3435 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3447 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3451 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_3469 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_3477 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3479 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3491 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3503 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3507 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3519 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3531 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3535 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3544 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_3556 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_3563 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_3571 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3588 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3591 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3603 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3615 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3619 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_3637 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_3645 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3647 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3659 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3671 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3675 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3687 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3699 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3703 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3715 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3727 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3731 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3742 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3754 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3759 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3771 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3783 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3787 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3799 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3811 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3815 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3827 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3839 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3843 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3855 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3867 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_3871 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_3879 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3896 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3899 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3911 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3923 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3927 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3939 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3943 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3952 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3955 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3967 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3979 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3983 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3995 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_4007 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_4011 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_4029 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_4037 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_4039 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_4051 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_4063 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_4067 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_4079 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_4091 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_4095 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_4113 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_4121 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_4123 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_4135 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_4147 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_4151 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_4163 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_4175 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_4179 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_4191 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_4203 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_4207 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_4219 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_4231 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_4235 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_4247 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_4259 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_4263 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_4275 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_4287 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_4291 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_4303 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_4315 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_4319 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_4331 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_4343 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_4347 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_4359 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_4371 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_4375 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_4387 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_4399 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_4403 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_4415 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_4427 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_4431 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_4443 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_4448 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_4452 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_4456 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_4459 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_4465 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_4469 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_4474 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_4478 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_4482 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_4487 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_4491 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_4495 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_4499 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_4503 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_4511 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_4515 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_4527 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_4539 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_4543 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_4555 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_4567 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_4571 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_928 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_942 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_946 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1112 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1413 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1425 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_1433 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2249 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2261 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2273 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2285 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2297 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_2301 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2303 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2315 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_2327 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_2335 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2340 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2344 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2348 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2352 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2356 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2359 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2368 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2372 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2376 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2380 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2384 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_2388 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2402 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2415 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_2427 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2444 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2456 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2468 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2471 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2483 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2495 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2507 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_2519 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_2525 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2527 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2535 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_2539 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2556 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2568 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2580 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_2583 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_2591 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2596 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2604 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2616 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_2628 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2636 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2639 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_2651 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2665 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2677 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2689 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_2693 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2707 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2719 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_2723 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2726 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2735 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_2747 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2751 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2760 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_2764 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2772 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2776 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2789 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2801 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_2805 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2807 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2819 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_2831 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2847 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_2859 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2863 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2875 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2887 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_2901 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2914 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2919 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2931 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2943 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2955 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_2967 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2972 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2975 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2988 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3000 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3012 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_3024 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3031 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3043 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_3055 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3070 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_3082 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3087 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3099 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3123 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_3135 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_3141 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3143 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_3155 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3179 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_3191 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_3197 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3199 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3211 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3235 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_3247 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_3251 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3255 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3259 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3268 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_3280 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3283 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3287 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3291 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3300 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3304 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3308 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3311 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3320 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3324 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3328 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_3332 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3340 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3352 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3364 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3367 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3379 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3391 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3403 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_3415 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_3421 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3423 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3435 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3447 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3459 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_3471 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_3477 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3479 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3491 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3503 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3515 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_3527 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_3533 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3535 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3547 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3559 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3571 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_3583 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_3589 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3591 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3603 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3615 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3627 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_3639 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_3645 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3647 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3659 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3671 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3683 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_3695 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_3701 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3703 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3715 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3727 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3739 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_3751 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_3757 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3759 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3771 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3783 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_3795 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_3801 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3804 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3808 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3812 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_3815 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3821 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3825 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3829 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3833 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3837 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3841 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3845 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3849 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3857 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3861 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3865 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_3869 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3871 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3875 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3879 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3883 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3887 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3891 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3895 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3899 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3903 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_3915 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_3923 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3927 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3939 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3951 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3963 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_3975 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_3981 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3983 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3995 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4007 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4019 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_4031 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_4037 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4039 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4051 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4063 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4075 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_4087 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_4093 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4095 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4107 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4119 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4131 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_4143 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_4149 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4151 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4163 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4175 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4187 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_4199 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_4205 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4207 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4219 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4231 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4243 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_4255 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_4261 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4263 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4275 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4287 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4299 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_4311 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_4317 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4319 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4331 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4343 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4355 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_4367 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_4373 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4375 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4387 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4399 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4411 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_4423 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_4429 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4431 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4443 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4455 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4467 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_4479 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_4485 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4487 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4499 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4511 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4523 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_4535 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_4541 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_4543 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_4549 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_4553 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_4557 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_4561 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_4565 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_4579 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1427 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1437 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2249 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_2273 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2275 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2287 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_2299 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_2303 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_2307 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_2316 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_2320 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_2328 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2331 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2343 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2355 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2367 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_2379 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_2385 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2387 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2399 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2411 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2423 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_2435 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_2441 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2443 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2455 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2467 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2479 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_2491 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_2497 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_2499 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_2507 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_2512 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2533 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_2545 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_2553 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2555 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2567 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2579 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2591 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_2603 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_2609 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_2611 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2623 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_2635 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_2643 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2654 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2667 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_2679 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_2687 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_2698 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_2702 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_2711 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_2719 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2723 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2735 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2747 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2759 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_2771 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_2777 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_2779 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_2791 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2795 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2807 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2819 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_2831 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_2835 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_2844 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2848 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2860 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2872 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_2884 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2891 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_2895 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_2898 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_2907 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2923 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_2935 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_2943 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_2947 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_2955 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_2959 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_2963 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_2975 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2979 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_2983 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_2991 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_2995 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_2999 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3003 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3007 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_3019 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3022 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3026 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3030 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3034 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3038 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3042 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3051 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_3055 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3059 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3063 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3067 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3071 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3075 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3079 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3091 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_3103 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_3111 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3115 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3127 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_3139 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3147 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3151 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3160 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_3164 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3171 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3183 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_3195 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3203 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3207 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_3216 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3224 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3227 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3239 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3251 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3263 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_3275 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_3281 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3283 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3295 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_3307 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3312 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3321 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3333 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_3337 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3339 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3351 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3355 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3359 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3368 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3380 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3392 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3395 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3407 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3419 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3431 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_3443 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_3449 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3451 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3463 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3475 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3487 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_3499 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_3505 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3507 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3519 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3531 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3543 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_3555 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_3561 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3563 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3575 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3587 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_3599 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3616 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3619 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3631 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3643 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3655 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_3667 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_3673 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3675 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3687 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3699 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3711 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_3723 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_3729 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3731 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3743 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_3755 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3772 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3784 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3787 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3799 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3811 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3823 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_3835 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_3841 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3843 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3855 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3867 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3879 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3883 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_3895 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3899 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3911 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3923 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3935 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_3947 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_3953 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3955 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3967 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3979 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3991 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_4003 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_4009 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4011 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4023 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4035 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4047 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_4059 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_4065 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4067 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4079 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4091 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4103 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_4115 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_4121 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4123 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4135 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4147 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4159 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_4171 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_4177 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4179 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4191 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4203 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4215 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_4227 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_4233 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4235 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4247 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4259 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4271 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_4283 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_4289 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4291 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4303 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4315 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4327 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_4339 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_4345 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4347 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4359 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4371 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4383 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_4395 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_4401 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4403 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4415 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4427 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4439 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_4451 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_4456 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_4459 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_4463 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_4466 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_4470 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_4474 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_4478 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_4486 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_4490 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_4494 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_4498 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_4502 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_4506 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_4510 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4515 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4527 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4539 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4551 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_4563 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_4569 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_4571 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_940 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1200 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1425 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1437 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_2249 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_2253 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_2257 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_2261 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_2265 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_2274 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_2278 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_2282 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_2286 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_2290 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_2294 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2303 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2315 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2327 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_2339 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_2348 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_2356 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_2359 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_2368 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2372 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2384 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2396 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_2408 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2415 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2427 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2439 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2451 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_2463 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_2469 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2471 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2483 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2495 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2507 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_2519 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_2525 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2527 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2539 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2551 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2563 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_2575 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_2581 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2583 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2595 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2607 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_2619 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_2636 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2639 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2651 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2663 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2675 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_2687 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_2693 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2707 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2719 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2731 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_2743 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_2749 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2751 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2763 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2775 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2787 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_2799 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_2805 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2807 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2819 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2831 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_2843 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2858 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2863 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2875 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2887 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_2899 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_2911 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_2917 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2919 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_2925 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_2929 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_2933 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_2945 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_2949 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_2957 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_2962 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_2971 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_2975 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2979 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2991 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3003 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_3015 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_3023 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3028 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3031 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3040 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3044 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_3056 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3064 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_3082 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3087 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3099 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3123 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_3135 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_3141 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3143 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3155 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3179 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_3191 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_3197 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3199 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3211 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3235 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_3247 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_3253 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3255 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3267 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3279 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3291 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_3303 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_3309 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3311 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3323 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3335 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3347 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_3359 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_3365 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_3367 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3372 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3381 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3397 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3409 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_3421 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3423 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3435 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3447 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3459 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_3471 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_3477 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3479 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3483 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3495 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3507 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3519 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_3531 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3535 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3547 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3559 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3571 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_3583 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_3589 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3591 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3603 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3615 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3627 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_3639 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_3645 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_3647 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3655 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3666 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3678 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3690 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3703 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3715 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3727 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3739 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_3751 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_3757 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3759 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3771 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3783 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_3795 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_3801 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_3811 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3815 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3827 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3839 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3851 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_3863 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_3869 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3871 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3883 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3895 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3907 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_3919 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_3925 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3927 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3939 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3951 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3963 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_3975 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_3981 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3983 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3995 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4007 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4019 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_4031 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_4037 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4039 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4051 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4063 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4075 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_4087 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_4093 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4095 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4107 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4119 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4131 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_4143 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_4149 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4151 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4163 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4175 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4187 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_4199 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_4205 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4207 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4219 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4231 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4243 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_4255 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_4261 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4263 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4275 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4287 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4299 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_4311 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_4317 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4319 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4331 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4343 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4355 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_4367 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_4373 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4375 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4387 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4399 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4411 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_4423 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_4429 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4431 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4443 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_4455 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4462 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4474 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4487 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4499 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4511 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4523 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_4535 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_4541 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4543 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4555 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4567 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_4579 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1384 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1396 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1441 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1453 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1457 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1463 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1480 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1490 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1494 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1498 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1502 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1506 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1510 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1513 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1522 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1526 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1531 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1535 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1539 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1541 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1545 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1548 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1552 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1556 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1560 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1564 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1569 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1573 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1595 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1601 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1607 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1619 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1625 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1637 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1645 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1648 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1653 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1662 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1667 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1671 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1675 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1679 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1681 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1685 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1694 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1698 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1704 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1709 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1713 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1716 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1720 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1724 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1730 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1749 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1761 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1765 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1777 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1790 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1793 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1802 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1806 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1818 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1821 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1825 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1835 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1847 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1849 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1857 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1860 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1875 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1877 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1881 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1889 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1896 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1905 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1916 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1920 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1924 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1928 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1933 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1949 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1952 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1956 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1961 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1965 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1969 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1972 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1976 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1985 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1989 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2002 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2006 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2012 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2017 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2025 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2029 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2033 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2039 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2057 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2085 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2097 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2101 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2105 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2108 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2112 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2116 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2120 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2124 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2129 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2133 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2136 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2140 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2144 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2148 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2152 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2157 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2166 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2180 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2185 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2189 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2193 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2197 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2201 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2205 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2210 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2213 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2217 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2221 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2265 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2282 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2294 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2321 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2325 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_2333 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2339 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2461 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2465 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2469 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2479 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2517 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2521 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2525 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2533 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2537 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2785 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2797 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_2801 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2809 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2826 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2993 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2997 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_3015 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_3023 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3025 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3037 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3049 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3065 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3093 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3121 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3149 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3177 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3205 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3233 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3245 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3249 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3261 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3273 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3289 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3301 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3317 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3329 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3345 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3357 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3373 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3389 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_3401 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3409 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3414 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3417 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3427 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3431 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3435 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3439 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_3443 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3445 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3449 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3453 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3457 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_3461 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3469 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_3473 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3479 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3483 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3492 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_3496 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3513 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3541 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3553 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3557 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3566 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3570 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3582 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3596 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_3608 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3625 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3653 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3681 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3709 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3737 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3749 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3765 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3777 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3781 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3793 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3805 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3821 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3849 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3861 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3865 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3877 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3889 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3905 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3917 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3933 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3961 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3973 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3989 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4017 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4045 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4073 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_4085 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4089 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4101 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_4113 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4117 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4129 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_4141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4145 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4157 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_4169 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4173 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4185 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_4197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4201 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4213 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_4225 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4229 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4241 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_4253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4257 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4269 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_4281 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4285 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4297 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_4309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4313 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4325 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_4337 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4341 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4353 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_4365 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4369 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4381 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_4393 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4397 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4409 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_4421 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4425 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4437 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_4449 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_4453 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_4459 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4462 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_4474 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4481 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4493 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_4505 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4509 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4521 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_4533 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4537 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4549 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_4561 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_4565 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_4579 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1455 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1457 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1467 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1471 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1480 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1484 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1488 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1492 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1496 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1500 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1504 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1508 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1513 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1517 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1525 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1529 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1533 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1537 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1545 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1549 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1552 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1556 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1560 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1576 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1588 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1600 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1612 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1632 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1644 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1652 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1656 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1660 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1664 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1668 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1672 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1676 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1681 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1685 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1689 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1694 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1702 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1706 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1712 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1715 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1727 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1749 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1761 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1767 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1776 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1787 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1791 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1797 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1809 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1820 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1832 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1836 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1844 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1905 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1917 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1920 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1924 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1928 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1932 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1936 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1940 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1944 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1948 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1952 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1956 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1961 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1965 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1969 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1973 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1977 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1981 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1985 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1996 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2000 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2004 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2008 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2012 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_2017 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2027 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2031 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2035 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2039 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2043 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2047 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2051 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2060 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2064 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2068 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2077 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2089 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_2101 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2109 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2112 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2116 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2120 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2124 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2129 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2133 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2136 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2140 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2144 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2148 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2152 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2156 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2160 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2164 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2168 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2172 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2176 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2180 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2185 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2192 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2198 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2202 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2212 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2216 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2220 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2229 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2575 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_2577 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_2585 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2590 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2599 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2615 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2627 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2725 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_2737 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2742 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2745 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2754 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2758 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2770 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2782 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_2794 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3005 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3017 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_3023 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3025 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3037 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3049 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3061 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3073 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_3079 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3093 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3117 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3129 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_3135 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3149 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3173 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3185 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_3191 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3229 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3241 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_3247 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3249 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3261 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3273 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3285 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3297 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_3303 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3317 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3329 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3341 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3353 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_3359 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3373 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3397 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3409 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_3415 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3429 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3453 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3465 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_3471 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3497 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3509 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3521 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_3527 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3541 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3565 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3577 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_3583 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3597 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3621 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3633 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_3639 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3641 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_3653 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_3657 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3660 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3664 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3668 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3672 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3681 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3685 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3689 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3697 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_3709 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3719 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3723 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3732 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_3744 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3765 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3777 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3789 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3801 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_3807 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3821 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3845 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3857 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_3863 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3865 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3877 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_3889 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3913 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_3919 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3933 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3957 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3969 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_3975 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3977 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3989 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4007 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4019 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4045 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4069 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_4081 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_4087 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4089 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4125 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_4137 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_4143 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4145 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4157 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4181 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_4193 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_4199 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4201 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4213 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4237 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_4249 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_4255 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4257 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4269 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4293 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_4305 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_4311 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4313 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4325 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4349 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_4361 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_4367 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4369 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_4381 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_4387 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_4390 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_4394 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_4398 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_4402 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_4406 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_4410 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_4414 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_4418 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_4422 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_4425 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_4429 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_4436 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_4440 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_4444 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_4448 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_4452 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_4456 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_4460 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_4466 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_4470 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_4474 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_4478 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_4481 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_4486 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4490 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4502 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4514 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_4526 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_4534 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4537 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4549 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4561 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_4573 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1441 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1453 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1462 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1471 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1476 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1480 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1492 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1496 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1500 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1504 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1508 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1512 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1516 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1520 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1526 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1530 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1534 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1651 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1653 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1661 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1664 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1668 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1672 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1676 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1680 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1696 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1763 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1765 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1775 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1781 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1821 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1833 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1931 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1933 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1940 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1944 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1948 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1952 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1956 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1960 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1964 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1968 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1972 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1976 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1980 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1984 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1989 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1993 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1996 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2000 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2006 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2012 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_2018 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_2022 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2026 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_2038 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2045 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2068 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2080 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2101 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_2113 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2119 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_2122 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_2126 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_2130 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_2134 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_2138 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_2142 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2146 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_2152 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2157 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2161 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_2164 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_2168 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2172 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_2177 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_2181 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_2185 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_2189 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2193 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2198 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_2210 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2629 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_2643 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_2647 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2997 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3009 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3021 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3033 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3045 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_3051 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3065 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3089 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3101 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_3107 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3121 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3145 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3157 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_3163 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3177 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3201 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3213 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_3219 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3233 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3245 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3257 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3269 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_3275 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3289 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3301 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3313 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3325 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_3331 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3345 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3357 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3369 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3381 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_3387 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3401 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3425 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3437 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_3443 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3457 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3481 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3493 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_3499 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3513 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3537 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3549 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_3555 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3569 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3593 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3605 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_3611 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3625 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3649 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3661 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_3667 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3681 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3705 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3717 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_3723 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3725 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_3737 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_3745 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3748 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3752 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3756 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3760 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3764 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3773 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_3777 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3781 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3785 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_3789 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_3793 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3796 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3805 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3809 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3813 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3817 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3821 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3825 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3829 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3849 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3861 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3873 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3885 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_3891 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3905 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3917 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3929 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3941 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_3947 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3961 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3973 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3985 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3997 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_4003 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4017 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4041 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_4053 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_4059 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4073 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4085 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4097 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_4109 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_4115 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4117 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4129 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4153 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_4165 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_4171 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4173 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4185 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4209 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_4221 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_4227 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4229 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4241 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4265 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_4277 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_4283 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4285 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4297 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4321 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_4333 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_4339 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4341 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4353 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4365 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4377 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_4389 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_4395 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4397 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4409 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4421 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4433 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_4445 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_4451 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4453 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4465 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4477 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4489 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_4501 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_4507 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4509 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4521 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4533 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4545 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_4557 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_4563 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4565 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_4577 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1469 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1488 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1492 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1496 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1500 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1504 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1508 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1513 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1517 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1520 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1524 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1536 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1548 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1560 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1649 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1661 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1669 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1673 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1817 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1829 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1837 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1843 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1929 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1941 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1949 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1954 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1958 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1961 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1965 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1968 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1972 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1976 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1982 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1986 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1991 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1996 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_2000 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_2004 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_2008 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2109 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2125 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2135 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2147 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2153 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_2156 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_2160 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_2164 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_2168 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2172 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2180 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2189 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2201 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3005 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3017 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_3023 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3025 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3037 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3049 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3061 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3073 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_3079 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3093 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3117 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3129 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_3135 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3149 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3173 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3185 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_3191 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3229 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3241 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_3247 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3249 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3261 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3273 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3285 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3297 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_3303 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3317 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3329 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3341 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3353 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_3359 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3373 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3397 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3409 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_3415 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3429 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3453 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3465 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_3471 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3497 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3509 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3521 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_3527 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3541 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3565 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3577 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_3583 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3597 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3621 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3633 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_3639 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3653 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3677 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3689 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_3695 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3709 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3733 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3745 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_3751 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3765 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3777 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3789 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3801 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_3807 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3821 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3845 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3857 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_3863 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3865 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3877 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3889 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3901 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3913 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_3919 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3933 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3957 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3969 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_3975 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3989 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4013 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_4025 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4045 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4069 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_4081 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_4087 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4089 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4125 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_4137 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_4143 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4145 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4157 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4181 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_4193 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_4199 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4201 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4213 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4237 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_4249 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_4255 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4257 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4269 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4293 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_4305 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_4311 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4313 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4325 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4349 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_4361 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_4367 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4369 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4381 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4393 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4405 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_4417 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_4423 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4425 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4437 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4449 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4461 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_4473 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_4479 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4481 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4493 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4505 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4517 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_4529 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_4535 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4537 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4549 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_4561 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_4579 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1493 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1496 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_1502 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1507 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1515 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1527 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1945 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1957 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1967 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_1971 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1976 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1984 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1993 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2005 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2155 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2165 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2177 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2189 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_2201 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2997 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3009 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3021 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3033 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3045 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3051 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3065 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3089 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3101 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3107 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3121 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3145 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3157 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3163 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3177 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3201 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3213 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3219 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3233 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3245 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3257 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3269 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3275 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3289 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3301 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3313 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3325 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3331 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3345 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3357 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3369 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3381 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3387 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3401 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3425 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3437 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3443 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3457 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3481 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3493 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3499 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3513 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3537 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3549 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3555 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3569 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3593 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3605 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3611 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3625 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3649 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3661 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3667 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3681 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3705 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3717 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3723 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3737 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3749 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3761 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3773 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3779 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3781 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3793 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3805 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3817 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3829 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3835 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3849 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3861 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3873 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3885 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3891 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3905 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3917 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3929 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3941 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3947 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3961 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3973 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3985 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3997 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_4003 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4017 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4041 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_4053 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_4059 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4073 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4085 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4097 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_4109 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_4115 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4117 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4129 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4153 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_4165 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_4171 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4173 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4185 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4209 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_4221 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_4227 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4229 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4241 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4265 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_4277 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_4283 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4285 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4297 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4321 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_4333 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_4339 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4341 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4353 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4377 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_4389 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_4395 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4397 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4409 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4421 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4433 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_4445 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_4451 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4453 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4465 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_4477 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4485 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_4497 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_4505 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_4509 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_4514 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_4518 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_4522 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4526 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4538 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4550 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_4562 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4565 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_4577 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3005 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3017 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3023 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3025 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3037 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3049 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3061 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3073 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3079 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3093 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3117 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3129 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3135 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3149 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3173 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3185 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3191 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3229 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3241 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3247 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3249 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3261 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3273 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3285 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3297 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3303 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3317 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3329 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3341 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3353 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3359 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3373 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3397 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3409 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3415 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3429 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3453 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3465 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3471 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3497 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3509 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3521 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3527 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3541 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3565 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3577 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3583 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3597 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3621 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3633 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3639 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3653 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3677 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3689 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3695 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3709 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3733 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3745 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3751 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3765 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3777 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3789 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3801 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3807 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3821 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3845 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3857 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3863 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3865 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3877 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3889 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3901 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3913 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3919 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3933 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3957 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3969 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3975 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3989 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4013 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_4025 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4045 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4069 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_4081 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_4087 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4089 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4125 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_4137 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_4143 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4145 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4157 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4181 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_4193 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_4199 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4201 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4213 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4237 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_4249 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_4255 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4257 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4269 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4293 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_4305 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_4311 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4313 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4325 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4349 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_4361 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_4367 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4369 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4381 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4393 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4405 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_4417 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_4423 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4425 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4437 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_4449 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_4457 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_4462 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_4466 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_4470 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_4474 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_4478 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_4481 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_4488 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_4492 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_4496 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_4500 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_4504 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_4508 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_4512 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_4518 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_4522 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_4526 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_4530 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_4534 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4537 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4549 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_4561 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_4565 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_4579 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2997 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3009 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3021 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3033 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3045 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_3051 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3065 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3089 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3101 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_3107 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3121 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3145 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3157 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_3163 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3177 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3201 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3213 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_3219 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3233 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3245 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3257 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3269 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_3275 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3289 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3301 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3313 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3325 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_3331 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3345 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3357 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3369 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3381 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_3387 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3401 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3425 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3437 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_3443 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3457 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3481 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3493 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_3499 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3513 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3537 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3549 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_3555 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3569 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3593 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3605 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_3611 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3625 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3649 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3661 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_3667 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3681 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3705 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3717 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_3723 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3737 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3749 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3761 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3773 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_3779 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3781 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3793 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3805 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3817 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3829 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_3835 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3849 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3861 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3873 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3885 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_3891 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3905 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3917 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3929 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3941 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_3947 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3961 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3973 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3985 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3997 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_4003 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4017 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4041 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_4053 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_4059 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4073 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4085 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4097 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_4109 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_4115 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4117 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4129 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4153 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_4165 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_4171 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4173 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4185 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4209 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_4221 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_4227 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4229 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4241 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4265 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_4277 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_4283 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4285 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4297 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4321 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_4333 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_4339 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4341 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4353 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4377 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_4389 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_4395 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4397 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4409 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4421 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4433 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_4445 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_4451 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4453 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4465 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4477 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4489 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_4501 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_4507 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_4509 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_4515 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_4518 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_4522 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4526 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4538 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4550 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_4562 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4565 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_4577 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3005 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3017 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3023 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3025 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3037 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3049 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3061 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3073 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3079 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3093 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3117 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3129 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3135 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3149 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3173 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3185 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3191 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3229 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3241 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3247 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3261 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3273 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3285 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3297 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3303 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3317 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3329 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3341 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3353 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3359 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3373 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3397 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3409 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3415 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3429 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3453 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3465 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3471 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3497 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3509 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3521 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3527 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3541 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3565 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3577 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3583 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3597 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3621 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3633 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3639 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3653 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3677 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3689 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3695 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3709 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3733 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3745 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3751 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3765 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3777 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3789 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3801 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3807 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3821 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3845 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3857 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3863 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3865 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3877 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3889 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3901 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3913 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3919 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3933 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3957 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3969 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3975 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3989 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4013 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_4025 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4045 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4069 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_4081 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_4087 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4089 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4125 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_4137 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_4143 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4145 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4157 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4181 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_4193 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_4199 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4201 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4213 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4237 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_4249 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_4255 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4257 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4269 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4293 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_4305 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_4311 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4313 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4325 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4349 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_4361 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_4367 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4369 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4381 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4393 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4405 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_4417 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_4423 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4425 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4437 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4449 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_4461 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_4469 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_4473 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_4479 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4481 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4493 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4505 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4517 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_4529 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_4535 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4537 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4549 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_4561 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_4565 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_4579 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2997 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3009 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3021 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3033 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3045 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_3051 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3065 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3089 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3101 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_3107 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3121 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3145 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3157 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_3163 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3177 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3201 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3213 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_3219 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3233 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3245 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3257 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3269 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_3275 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3289 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3301 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3313 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3325 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_3331 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3345 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3357 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3369 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3381 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_3387 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3401 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3425 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3437 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_3443 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3457 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3481 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3493 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_3499 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3513 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3537 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3549 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_3555 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3569 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3593 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3605 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_3611 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3625 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3649 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3661 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_3667 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3681 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3705 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3717 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_3723 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3737 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3749 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3761 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3773 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_3779 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3781 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3793 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3805 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3817 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3829 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_3835 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3849 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3861 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3873 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3885 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_3891 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3905 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3917 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3929 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3941 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_3947 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3961 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3973 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3985 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3997 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_4003 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4017 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4041 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_4053 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_4059 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4073 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4085 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4097 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_4109 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_4115 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4117 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4129 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4153 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_4165 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_4171 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4173 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4185 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4209 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_4221 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_4227 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4229 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4241 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4265 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_4277 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_4283 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4285 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4297 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4321 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_4333 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_4339 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4341 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4353 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4377 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_4389 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_4395 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4397 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4409 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4421 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4433 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_4445 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_4451 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4453 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4465 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4480 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4492 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_4504 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4509 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4521 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4533 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4545 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_4557 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_4563 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4565 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_4577 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3005 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3017 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_3023 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3025 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3037 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3049 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3061 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3073 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_3079 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3093 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3117 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3129 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_3135 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3149 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3173 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3185 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_3191 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3229 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3241 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_3247 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3261 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3273 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3285 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3297 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_3303 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3317 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3329 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3341 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3353 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_3359 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3373 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3397 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3409 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_3415 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3429 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3453 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3465 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_3471 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3497 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3509 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3521 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_3527 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3541 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3565 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3577 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_3583 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3597 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3621 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3633 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_3639 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3653 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3677 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3689 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_3695 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3709 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3733 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3745 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_3751 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3765 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3777 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3789 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3801 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_3807 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3821 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3845 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3857 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_3863 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3865 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3877 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3889 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3901 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3913 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_3919 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3933 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3957 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3969 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_3975 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3989 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4013 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_4025 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4045 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4069 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_4081 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_4087 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4089 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4125 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_4137 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_4143 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4145 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4157 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4181 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_4193 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_4199 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4201 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4213 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4237 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_4249 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_4255 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4257 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4269 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4293 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_4305 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_4311 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4313 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4325 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4349 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_4361 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_4367 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4369 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4381 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4393 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4405 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_4417 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_4423 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4425 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4437 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4449 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4461 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_4473 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_4479 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4481 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4493 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4505 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4517 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_4529 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_4535 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4537 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_4549 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_4557 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_4561 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_4565 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_4579 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2997 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3009 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3021 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3033 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3045 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_3051 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3065 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3089 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3101 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_3107 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3121 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3145 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3157 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_3163 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3177 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3201 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3213 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_3219 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3233 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3245 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3257 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3269 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_3275 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3289 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3301 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3313 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3325 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_3331 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3345 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3357 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3369 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3381 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_3387 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3401 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3425 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3437 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_3443 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3457 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3481 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3493 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_3499 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3513 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3537 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3549 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_3555 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3569 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3593 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3605 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_3611 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3625 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3649 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3661 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_3667 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3681 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3705 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3717 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_3723 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3737 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3749 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3761 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3773 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_3779 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3781 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3793 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3805 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3817 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3829 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_3835 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3849 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3861 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3873 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3885 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_3891 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3905 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3917 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3929 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3941 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_3947 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3961 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3973 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3985 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3997 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_4003 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4017 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4041 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_4053 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_4059 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4073 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4085 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4097 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_4109 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_4115 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4117 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4129 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4153 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_4165 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_4171 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4173 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4185 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4209 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_4221 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_4227 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4229 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4241 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4265 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_4277 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_4283 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4285 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4297 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4321 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_4333 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_4339 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4341 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4353 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4365 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4377 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_4389 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_4395 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4397 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4409 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4421 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4433 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_4445 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_4451 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4453 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4465 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4477 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4489 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_4501 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_4507 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4509 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4521 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4533 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4545 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_4557 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_4563 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4565 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_4577 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3005 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3017 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_3023 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3025 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3037 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3049 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3061 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3073 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_3079 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3093 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3117 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3129 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_3135 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3149 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3173 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3185 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_3191 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3229 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3241 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_3247 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3249 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3261 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3273 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3285 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3297 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_3303 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3317 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3329 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3341 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3353 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_3359 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3373 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3397 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3409 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_3415 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3429 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3453 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3465 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_3471 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3497 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3509 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3521 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_3527 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3541 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3565 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3577 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_3583 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3597 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3621 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3633 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_3639 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3653 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3677 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3689 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_3695 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3709 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3733 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3745 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_3751 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3765 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3777 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3789 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3801 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_3807 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3821 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3845 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3857 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_3863 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3865 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3877 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3889 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3901 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3913 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_3919 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3933 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3957 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3969 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_3975 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3989 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4013 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_4025 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4045 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4069 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_4081 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_4087 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4089 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4125 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_4137 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_4143 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4145 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4157 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4181 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_4193 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_4199 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4201 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4213 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4237 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_4249 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_4255 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4257 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4269 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4293 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_4305 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_4311 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4313 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4325 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4349 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_4361 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_4367 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4369 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4381 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4393 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4405 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_4417 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_4423 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4425 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4437 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4449 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4461 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_4473 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_4479 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4481 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4493 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4505 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4517 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_4529 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_4535 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4537 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4549 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4561 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_4573 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2997 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3009 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3021 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3033 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3045 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_3051 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3065 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3089 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3101 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_3107 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3121 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3145 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3157 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_3163 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3177 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3201 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3213 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_3219 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3233 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3245 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3257 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3269 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_3275 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3289 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3301 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3313 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3325 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_3331 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3345 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3357 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3369 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3381 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_3387 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3401 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3425 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3437 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_3443 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3457 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3481 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3493 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_3499 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3513 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3537 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3549 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_3555 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3569 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3593 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3605 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_3611 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3625 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3649 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3661 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_3667 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3681 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3705 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3717 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_3723 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3737 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3749 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3761 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3773 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_3779 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3781 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3793 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3805 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3817 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3829 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_3835 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3849 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3861 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3873 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3885 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_3891 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3905 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3917 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3929 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3941 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_3947 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3961 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3973 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3985 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3997 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_4003 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4017 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4041 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_4053 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_4059 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4073 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4085 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4097 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_4109 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_4115 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4117 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4129 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4153 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_4165 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_4171 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4173 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4185 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4209 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_4221 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_4227 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4229 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4241 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4265 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_4277 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_4283 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4285 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4297 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4321 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_4333 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_4339 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4341 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4353 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4365 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4377 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_4389 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_4395 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4397 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4409 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4421 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4433 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_4445 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_4451 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4453 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4465 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4477 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4489 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_4501 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_4507 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_4509 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_4514 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_4518 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_4522 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4526 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4538 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_4550 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_4558 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_4562 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_4565 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_4579 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3005 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3017 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_3023 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3025 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3037 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3049 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3061 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3073 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_3079 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3093 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3117 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3129 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_3135 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3149 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3173 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3185 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_3191 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3229 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3241 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_3247 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3249 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3261 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3273 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3285 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3297 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_3303 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3317 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3329 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3341 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3353 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_3359 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3373 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3397 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3409 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_3415 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3429 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3453 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3465 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_3471 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3497 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3509 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3521 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_3527 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3541 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3565 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3577 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_3583 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3597 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3621 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3633 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_3639 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3653 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3677 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3689 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_3695 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3709 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3733 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3745 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_3751 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3765 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3777 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3789 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3801 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_3807 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3821 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3845 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3857 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_3863 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3865 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3877 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3889 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3901 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3913 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_3919 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3933 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3957 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3969 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_3975 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3989 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4013 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_4025 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4045 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4069 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_4081 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_4087 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4089 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4125 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_4137 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_4143 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4145 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4157 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4181 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_4193 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_4199 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4201 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4213 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4237 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_4249 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_4255 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4257 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4269 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4293 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_4305 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_4311 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4313 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4325 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4349 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_4361 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_4367 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4369 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4381 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4393 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4405 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_4417 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_4423 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4425 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4437 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_4449 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_4457 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_4462 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_4466 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_4470 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_4474 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_4478 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_4481 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_4488 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_4492 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_4496 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_4500 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_4504 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_4508 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_4512 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_4518 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_4522 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_4526 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_4530 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_4534 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4537 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4549 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4561 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_4573 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2997 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3009 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3021 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3033 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3045 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_3051 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3065 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3089 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3101 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_3107 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3121 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3145 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3157 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_3163 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3177 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3201 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3213 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_3219 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3233 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3245 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3257 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3269 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_3275 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3289 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3301 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3313 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3325 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_3331 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3345 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3357 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3369 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3381 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_3387 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3401 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3425 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3437 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_3443 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3457 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3481 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3493 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_3499 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3513 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3537 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3549 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_3555 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3569 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3593 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3605 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_3611 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3625 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3649 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3661 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_3667 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3681 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3705 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3717 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_3723 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3737 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3749 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3761 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3773 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_3779 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3781 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3793 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3805 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3817 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3829 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_3835 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3849 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3861 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3873 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3885 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_3891 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3905 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3917 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3929 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3941 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_3947 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3961 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3973 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3985 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3997 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_4003 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4017 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4041 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_4053 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_4059 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4073 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4085 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4097 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_4109 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_4115 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4117 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4129 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4153 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_4165 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_4171 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4173 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4185 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4209 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_4221 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_4227 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4229 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4241 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4265 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_4277 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_4283 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4285 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4297 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4321 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_4333 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_4339 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4341 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4353 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4365 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4377 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_4389 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_4395 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4397 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4409 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4421 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4433 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_4445 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_4451 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4453 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4465 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4477 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4489 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_4501 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_4507 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_4509 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_4515 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_4518 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_4522 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4526 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4538 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4550 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_4562 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_4565 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_4579 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3005 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3017 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_3023 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3025 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3037 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3049 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3061 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3073 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_3079 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3093 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3117 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3129 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_3135 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3149 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3173 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3185 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_3191 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3229 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3241 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_3247 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3261 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3273 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3285 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3297 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_3303 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3317 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3329 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3341 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3353 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_3359 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3373 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3397 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3409 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_3415 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3429 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3453 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3465 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_3471 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3497 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3509 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3521 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_3527 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3541 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3565 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3577 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_3583 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3597 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3621 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3633 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_3639 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3653 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3677 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3689 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_3695 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3709 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3733 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3745 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_3751 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3765 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3777 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3789 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3801 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_3807 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3821 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3845 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3857 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_3863 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3865 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3877 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3889 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3901 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3913 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_3919 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3933 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3957 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3969 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_3975 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3989 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4013 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_4025 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4045 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4069 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_4081 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_4087 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4089 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4125 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_4137 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_4143 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4145 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4157 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4181 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_4193 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_4199 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4201 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4213 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4237 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_4249 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_4255 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4257 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4269 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4293 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_4305 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_4311 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4313 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4325 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4349 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_4361 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_4367 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4369 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4381 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4393 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4405 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_4417 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_4423 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4425 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4437 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4449 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4461 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_4473 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_4479 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4481 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4493 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4505 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4517 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_4529 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_4535 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4537 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4549 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4561 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_4573 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2997 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3009 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3021 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3033 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3045 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3051 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3065 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3089 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3101 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3107 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3121 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3145 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3157 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3163 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3177 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3201 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3213 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3219 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3233 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3245 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3257 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3269 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3275 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3289 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3301 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3313 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3325 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3331 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3345 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3357 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3369 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3381 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3387 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3401 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3425 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3437 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3443 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3457 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3481 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3493 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3499 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3513 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3537 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3549 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3555 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3569 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3593 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3605 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3611 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3625 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3649 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3661 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3667 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3681 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3705 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3717 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3723 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3737 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3749 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3761 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3773 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3779 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3781 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3793 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3805 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3817 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3829 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3835 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3849 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3861 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3873 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3885 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3891 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3905 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3917 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3929 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3941 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3947 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3961 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3973 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3985 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3997 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_4003 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4017 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4041 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_4053 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_4059 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4073 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4085 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4097 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_4109 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_4115 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4117 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4129 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4153 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_4165 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_4171 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4173 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4185 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4209 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_4221 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_4227 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4229 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4241 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4265 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_4277 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_4283 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4285 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4297 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4321 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_4333 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_4339 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4341 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4353 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4377 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_4389 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_4395 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4397 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4409 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4421 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4433 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_4445 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_4451 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4453 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4465 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4477 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4489 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_4501 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_4507 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4509 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4521 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4533 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4545 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_4557 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_4563 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_4565 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_4579 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3005 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_3017 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_3023 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3025 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3037 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3049 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3061 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_3073 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_3079 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3093 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3117 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_3129 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_3135 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3149 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3173 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_3185 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_3191 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3229 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_3241 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_3247 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3249 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3261 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3273 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3285 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_3297 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_3303 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3317 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3329 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3341 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_3353 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_3359 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3373 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3397 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_3409 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_3415 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3429 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3453 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_3465 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_3471 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3497 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3509 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_3521 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_3527 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3541 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3565 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_3577 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_3583 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3597 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3621 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_3633 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_3639 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3653 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3677 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_3689 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_3695 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3709 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3733 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_3745 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_3751 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3765 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3777 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3789 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_3801 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_3807 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3821 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3845 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_3857 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_3863 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3865 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3877 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3889 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3901 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_3913 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_3919 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3933 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3957 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_3969 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_3975 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3989 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4013 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_4025 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4045 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4069 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_4081 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_4087 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4089 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4125 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_4137 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_4143 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4145 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4157 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4181 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_4193 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_4199 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4201 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4213 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4237 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_4249 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_4255 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4257 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4269 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4293 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_4305 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_4311 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4313 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4325 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4349 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_4361 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_4367 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4369 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4381 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4393 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4405 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_4417 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_4423 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4425 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4437 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4449 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4461 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_4473 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_4479 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_4481 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4486 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4498 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4510 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4522 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_4534 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4537 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4549 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4561 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_4573 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2997 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3009 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3021 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3033 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3045 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3051 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3065 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3089 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3101 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3107 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3121 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3145 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3157 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3163 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3177 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3201 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3213 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3219 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3233 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3245 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3257 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3269 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3275 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3289 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3301 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3313 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3325 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3331 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3345 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3357 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3369 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3381 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3387 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3401 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3425 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3437 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3443 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3457 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3481 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3493 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3499 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3513 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3537 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3549 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3555 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3569 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3593 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3605 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3611 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3625 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3649 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3661 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3667 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3681 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3705 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3717 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3723 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3737 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3749 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3761 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3773 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3779 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3781 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3793 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3805 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3817 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3829 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3835 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3849 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3861 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3873 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3885 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3891 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3905 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3917 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3929 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3941 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3947 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3961 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3973 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3985 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3997 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_4003 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4017 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4041 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_4053 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_4059 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4073 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4085 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4097 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_4109 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_4115 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4117 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4129 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4153 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_4165 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_4171 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4173 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4185 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4209 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_4221 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_4227 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4229 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4241 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4265 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_4277 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_4283 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4285 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4297 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4321 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_4333 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_4339 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4341 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4353 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4377 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_4389 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_4395 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4397 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4409 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4421 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4433 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_4445 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_4451 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4453 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4465 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_4477 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4484 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4496 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4509 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4521 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4533 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4545 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_4557 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_4563 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_4565 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_4579 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3005 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3017 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_3023 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3025 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3037 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3049 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3061 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3073 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_3079 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3093 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3117 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3129 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_3135 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3149 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3173 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3185 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_3191 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3229 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3241 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_3247 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3249 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3261 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3273 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3285 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3297 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_3303 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3317 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3329 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3341 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3353 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_3359 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3373 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3397 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3409 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_3415 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3429 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3453 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3465 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_3471 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3497 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3509 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3521 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_3527 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3541 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3565 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3577 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_3583 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3597 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3621 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3633 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_3639 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3653 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3677 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3689 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_3695 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3709 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3733 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3745 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_3751 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3765 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3777 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3789 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3801 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_3807 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3821 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3845 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3857 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_3863 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3865 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3877 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3889 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3901 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3913 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_3919 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3933 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3957 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3969 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_3975 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3989 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4013 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_4025 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4045 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4069 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_4081 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_4087 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4089 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4125 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_4137 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_4143 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4145 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4157 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4181 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_4193 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_4199 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4201 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4213 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4237 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_4249 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_4255 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4257 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4269 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4293 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_4305 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_4311 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4313 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4325 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4349 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_4361 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_4367 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4369 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4381 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4393 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4405 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_4417 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_4423 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4425 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4437 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4449 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4461 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_4473 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_4479 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4481 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4493 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4505 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4517 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_4529 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_4535 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4537 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4549 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4561 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_4573 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2997 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3009 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3021 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3033 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3045 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_3051 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3065 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3089 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3101 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_3107 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3121 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3145 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3157 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_3163 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3177 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3201 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3213 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_3219 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3233 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3245 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3257 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3269 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_3275 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3289 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3301 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3313 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3325 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_3331 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3345 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3357 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3369 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3381 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_3387 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3401 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3425 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3437 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_3443 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3457 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3481 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3493 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_3499 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3513 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3537 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3549 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_3555 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3569 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3593 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3605 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_3611 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3625 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3649 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3661 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_3667 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3681 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3705 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3717 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_3723 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3737 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3749 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3761 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3773 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_3779 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3781 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3793 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3805 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3817 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3829 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_3835 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3849 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3861 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3873 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3885 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_3891 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3905 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3917 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3929 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3941 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_3947 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3961 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3973 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3985 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3997 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_4003 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4017 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4041 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_4053 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_4059 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4073 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4085 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4097 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_4109 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_4115 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4117 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4129 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4153 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_4165 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_4171 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4173 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4185 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4209 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_4221 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_4227 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4229 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4241 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4265 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_4277 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_4283 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4285 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4297 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4321 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_4333 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_4339 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4341 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4353 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4377 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_4389 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_4395 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4397 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4409 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4421 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4433 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_4445 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_4451 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4453 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4465 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4477 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4489 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_4501 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_4507 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4509 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4521 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4533 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4545 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_4557 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_4563 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4565 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_4577 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3005 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3017 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_3023 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3025 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3037 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3049 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3061 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3073 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_3079 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3093 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3117 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3129 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_3135 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3149 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3173 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3185 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_3191 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3229 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3241 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_3247 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3261 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3273 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3285 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3297 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_3303 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3317 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3329 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3341 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3353 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_3359 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3373 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3397 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3409 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_3415 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3429 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3453 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3465 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_3471 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3497 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3509 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3521 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_3527 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3541 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3565 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3577 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_3583 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3597 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3621 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3633 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_3639 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3653 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3677 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3689 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_3695 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3709 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3733 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3745 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_3751 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3765 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3777 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3789 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3801 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_3807 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3821 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3845 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3857 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_3863 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3865 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3877 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3889 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3901 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3913 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_3919 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3933 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3957 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3969 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_3975 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3989 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4013 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_4025 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4045 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4069 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_4081 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_4087 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4089 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4125 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_4137 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_4143 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4145 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4157 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4181 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_4193 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_4199 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4201 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4213 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4237 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_4249 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_4255 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4257 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4269 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4293 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_4305 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_4311 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4313 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4325 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4349 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_4361 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_4367 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4369 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4381 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4393 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4405 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_4417 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_4423 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4425 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4437 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4449 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4461 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_4473 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_4479 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4481 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4493 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4505 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4517 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_4529 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_4535 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4537 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4549 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4561 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_4579 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2997 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3009 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3021 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3033 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_3045 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_3051 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3065 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3089 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_3101 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_3107 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3121 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3145 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_3157 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_3163 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3177 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3201 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_3213 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_3219 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3233 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3245 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3257 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_3269 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_3275 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3289 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3301 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3313 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_3325 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_3331 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3345 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3357 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3369 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_3381 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_3387 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3401 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3425 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_3437 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_3443 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3457 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3481 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_3493 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_3499 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3513 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3537 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_3549 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_3555 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3569 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3593 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_3605 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_3611 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3625 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3649 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_3661 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_3667 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3681 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3705 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_3717 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_3723 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3737 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3749 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3761 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_3773 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_3779 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3781 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3793 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3805 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3817 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_3829 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_3835 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3849 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3861 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3873 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_3885 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_3891 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3905 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3917 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3929 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_3941 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_3947 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3961 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3973 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3985 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_3997 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_4003 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4017 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4041 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_4053 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_4059 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4073 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4085 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4097 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_4109 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_4115 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4117 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4129 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4153 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_4165 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_4171 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4173 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4185 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4209 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_4221 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_4227 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4229 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4241 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4265 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_4277 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_4283 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4285 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4297 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4321 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_4333 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_4339 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4341 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4353 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4377 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_4389 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_4395 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4397 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4409 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4421 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4433 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_4445 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_4451 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4453 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4465 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4477 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4489 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_4501 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_4507 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4509 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4521 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4533 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4545 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_4557 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_4563 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4565 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_4577 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1749 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1774 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1786 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3005 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3017 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_3023 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3025 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3037 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3049 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3061 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3073 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_3079 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3093 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3117 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3129 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_3135 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3149 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3173 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3185 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_3191 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3229 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3241 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_3247 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3249 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3261 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3273 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3285 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3297 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_3303 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3317 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3329 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3341 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3353 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_3359 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3373 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3397 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3409 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_3415 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3429 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3453 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3465 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_3471 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3497 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3509 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3521 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_3527 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3541 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3565 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3577 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_3583 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3597 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3621 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3633 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_3639 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3653 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3677 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3689 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_3695 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3709 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3733 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3745 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_3751 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3765 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3777 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3789 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3801 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_3807 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3821 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3845 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3857 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_3863 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3865 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3877 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3889 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3901 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3913 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_3919 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3933 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3957 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3969 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_3975 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3989 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4013 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_4025 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4045 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4069 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_4081 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_4087 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4089 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4125 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_4137 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_4143 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4145 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4157 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4181 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_4193 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_4199 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4201 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4213 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4237 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_4249 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_4255 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4257 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4269 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4293 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_4305 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_4311 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4313 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4325 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4349 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_4361 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_4367 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4369 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4381 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4393 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4405 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_4417 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_4423 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4425 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4437 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4449 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4461 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_4473 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_4479 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4481 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4493 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4505 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4517 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_4529 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_4535 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4537 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4549 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4561 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_4579 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_976 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1000 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1054 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1066 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1108 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1219 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1275 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1283 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1337 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1351 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1385 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1405 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1427 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1437 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1450 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1462 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1483 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1491 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1504 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1516 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1531 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1539 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1541 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1545 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1558 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1570 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1585 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1593 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1612 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1624 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1639 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1651 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1667 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1705 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1723 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1747 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1759 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1763 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1783 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1795 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1810 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1818 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1837 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1864 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1891 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1918 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1930 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1947 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1972 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1984 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1989 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_2003 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_2011 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2026 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_2038 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_2045 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_2059 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_2067 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_2080 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_2084 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_2098 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2101 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_2113 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_2121 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_2134 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2152 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2157 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_2169 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_2175 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_2188 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_2206 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2233 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_2245 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_2260 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2287 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2299 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2311 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_2323 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2325 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2341 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_2357 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_2377 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_2381 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_2389 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2404 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_2416 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2431 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_2435 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_2437 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_2445 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2458 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_2470 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_2491 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_2493 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_2499 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2512 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_2524 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_2539 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_2547 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2549 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_2553 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_2566 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_2570 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_2578 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_2593 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_2601 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_2605 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_2620 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_2624 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_2632 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2647 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_2659 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_2661 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2675 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_2679 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2692 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2704 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_2717 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2731 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2747 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2759 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_2771 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_2773 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2787 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2803 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2815 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_2827 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_2829 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2843 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_2859 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_2867 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_2881 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_2885 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_2893 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2908 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_2920 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2935 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_2939 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_2941 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_2949 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2962 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_2974 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_2995 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_2997 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_3003 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3016 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3032 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_3044 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3053 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_3057 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3070 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_3086 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3106 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3133 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_3145 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3160 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_3165 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3173 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3187 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_3199 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_3214 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3241 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_3253 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_3268 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3295 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_3307 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_3322 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3330 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3349 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3376 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3389 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_3403 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3421 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_3433 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_3441 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3445 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3459 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3475 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3487 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_3499 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3513 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3517 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3531 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3543 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_3555 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3557 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3571 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_3587 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_3595 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3610 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3637 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_3649 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3664 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_3669 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3677 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3691 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_3703 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_3718 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_3725 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3743 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3747 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3761 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_3773 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_3779 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_3781 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3799 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3815 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_3827 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_3835 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3837 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3853 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_3869 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_3889 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_3893 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_3901 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3916 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_3928 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3943 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_3947 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_3949 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_3957 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3970 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_3982 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_3997 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_4003 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_4005 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_4011 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_4024 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_4036 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_4051 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_4059 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_4061 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_4065 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_4078 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_4090 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_4105 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_4113 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_4117 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_4132 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_4144 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_4159 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_4171 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_4173 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_4187 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_4191 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_4204 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_4216 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_4229 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_4243 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_4259 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_4271 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_4283 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_4285 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_4299 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_4315 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_4327 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_4339 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_4341 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_4355 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_4371 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_4379 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_4393 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_4397 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_4405 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_4420 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_4432 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_4447 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_4451 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_4453 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_4461 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_4474 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_4486 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_4501 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_4507 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_4509 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_4521 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_4533 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_4545 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_4557 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_4563 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_4565 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_4577 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1357 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1370 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1373 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1381 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1396 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1413 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1426 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1441 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1469 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1482 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1497 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1510 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1513 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1525 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1538 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1541 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1553 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1566 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1569 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1581 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1594 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1597 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1621 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1625 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1633 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1648 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1653 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1661 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1675 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1679 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1681 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1702 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1709 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1735 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1737 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1743 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1765 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1777 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1790 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1793 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1805 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1818 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1821 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1833 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1846 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1849 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1861 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1874 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1877 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1889 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1902 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1905 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1917 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1930 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1933 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1945 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1958 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1961 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1973 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1986 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1989 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2001 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2014 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2017 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2029 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2042 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2045 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2057 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2070 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2073 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2085 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2098 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2101 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2129 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2141 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2154 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_2157 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2165 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_2179 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2185 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2197 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2210 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2213 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2225 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2238 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_2241 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2249 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2252 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2266 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2269 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2281 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2294 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_2297 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2301 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_2314 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2322 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2339 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2351 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2368 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2395 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2407 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2423 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2435 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2451 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2463 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2479 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2491 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2507 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2519 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2535 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2547 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2563 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2575 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2591 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2603 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2619 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2631 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2633 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2647 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_2651 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2659 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2675 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2687 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2703 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2715 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2731 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2743 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2759 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2771 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2787 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2799 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2815 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2827 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2843 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2855 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2871 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2883 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2899 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2911 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2927 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2939 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2955 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2967 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_2983 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2995 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2997 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3011 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3023 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_3025 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_3043 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3051 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3067 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3079 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_3081 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_3097 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_3105 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3124 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3151 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3163 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3179 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3191 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3207 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3219 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3235 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3247 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3249 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3263 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3275 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3291 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3303 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3319 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3331 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3347 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3359 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3375 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3387 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3403 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3415 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3431 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3443 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3459 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3471 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3487 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3499 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3501 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3515 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_3519 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3527 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3543 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3555 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3571 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3583 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3599 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3611 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3627 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3639 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3641 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3655 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_3659 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3667 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3683 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3695 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3711 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3723 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3739 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3751 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_3753 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3759 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_3772 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3781 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3795 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3807 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_3809 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3813 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_3826 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3834 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3851 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3863 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_3865 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3880 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3907 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3919 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3935 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3947 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3963 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3975 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3991 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_4003 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_4019 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_4031 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_4047 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_4059 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_4075 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_4087 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_4089 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_4103 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_4115 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_4117 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_4131 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_4143 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_4145 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_4159 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_4171 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_4173 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_4187 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_4199 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_4201 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_4215 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_4227 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_4229 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_4243 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_4255 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_4257 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_4271 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_4283 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_4285 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_4299 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_4311 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_4313 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_4327 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_4339 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_4341 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_4355 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_4367 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_4369 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_4383 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_4395 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_4397 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_4411 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_4423 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_4425 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_4439 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_4451 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_4453 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_4467 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_4479 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_4481 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_4495 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_4507 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_4509 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_4523 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_4535 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_4537 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_4549 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_4561 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_4565 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_4579 ();
endmodule

