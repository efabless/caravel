magic
tech sky130A
timestamp 1641854866
<< checkpaint >>
rect -33284 -139989 326776 380071
<< metal2 >>
rect 4043 351760 4099 352480
rect 12139 351760 12195 352480
rect 20235 351760 20291 352480
rect 28377 351760 28433 352480
rect 36473 351760 36529 352480
rect 44569 351760 44625 352480
rect 52711 351760 52767 352480
rect 60807 351760 60863 352480
rect 68903 351760 68959 352480
rect 77045 351760 77101 352480
rect 85141 351760 85197 352480
rect 93237 351760 93293 352480
rect 101379 351760 101435 352480
rect 109475 351760 109531 352480
rect 117571 351760 117627 352480
rect 125713 351760 125769 352480
rect 133809 351760 133865 352480
rect 141905 351760 141961 352480
rect 150047 351760 150103 352480
rect 158143 351760 158199 352480
rect 166239 351760 166295 352480
rect 174381 351760 174437 352480
rect 182477 351760 182533 352480
rect 190573 351760 190629 352480
rect 198715 351760 198771 352480
rect 206811 351760 206867 352480
rect 214907 351760 214963 352480
rect 223049 351760 223105 352480
rect 231145 351760 231201 352480
rect 239241 351760 239297 352480
rect 247383 351760 247439 352480
rect 255479 351760 255535 352480
rect 263575 351760 263631 352480
rect 271717 351760 271773 352480
rect 279813 351760 279869 352480
rect 287909 351760 287965 352480
rect 227179 -480 227235 240
rect 227731 -480 227787 240
rect 228329 -480 228385 240
rect 228927 -480 228983 240
rect 229525 -480 229581 240
rect 230123 -480 230179 240
rect 230721 -480 230777 240
rect 231273 -480 231329 240
rect 231871 -480 231927 240
rect 232469 -480 232525 240
rect 233067 -480 233123 240
rect 233665 -480 233721 240
rect 234263 -480 234319 240
rect 234861 -480 234917 240
rect 235413 -480 235469 240
rect 236011 -480 236067 240
rect 236609 -480 236665 240
rect 237207 -480 237263 240
rect 237805 -480 237861 240
rect 238403 -480 238459 240
rect 239001 -480 239057 240
rect 239553 -480 239609 240
rect 240151 -480 240207 240
rect 240749 -480 240805 240
rect 241347 -480 241403 240
rect 241945 -480 242001 240
rect 242543 -480 242599 240
rect 243095 -480 243151 240
rect 243693 -480 243749 240
rect 244291 -480 244347 240
rect 244889 -480 244945 240
rect 245487 -480 245543 240
rect 246085 -480 246141 240
rect 246683 -480 246739 240
rect 247235 -480 247291 240
rect 247833 -480 247889 240
rect 248431 -480 248487 240
rect 249029 -480 249085 240
rect 249627 -480 249683 240
rect 250225 -480 250281 240
rect 250823 -480 250879 240
rect 251375 -480 251431 240
rect 251973 -480 252029 240
rect 252571 -480 252627 240
rect 253169 -480 253225 240
rect 253767 -480 253823 240
rect 254365 -480 254421 240
rect 254917 -480 254973 240
rect 255515 -480 255571 240
rect 256113 -480 256169 240
rect 256711 -480 256767 240
rect 257309 -480 257365 240
rect 257907 -480 257963 240
rect 258505 -480 258561 240
rect 259057 -480 259113 240
rect 259655 -480 259711 240
rect 260253 -480 260309 240
rect 260851 -480 260907 240
rect 261449 -480 261505 240
rect 262047 -480 262103 240
rect 262645 -480 262701 240
rect 263197 -480 263253 240
rect 263795 -480 263851 240
rect 264393 -480 264449 240
rect 264991 -480 265047 240
rect 265589 -480 265645 240
rect 266187 -480 266243 240
rect 266739 -480 266795 240
rect 267337 -480 267393 240
rect 267935 -480 267991 240
rect 268533 -480 268589 240
rect 269131 -480 269187 240
rect 269729 -480 269785 240
rect 270327 -480 270383 240
rect 270879 -480 270935 240
rect 271477 -480 271533 240
rect 272075 -480 272131 240
rect 272673 -480 272729 240
rect 273271 -480 273327 240
rect 273869 -480 273925 240
rect 274467 -480 274523 240
rect 275019 -480 275075 240
rect 275617 -480 275673 240
rect 276215 -480 276271 240
rect 276813 -480 276869 240
rect 277411 -480 277467 240
rect 278009 -480 278065 240
rect 278561 -480 278617 240
rect 279159 -480 279215 240
rect 279757 -480 279813 240
rect 280355 -480 280411 240
rect 280953 -480 281009 240
rect 281551 -480 281607 240
rect 282149 -480 282205 240
rect 282701 -480 282757 240
rect 283299 -480 283355 240
rect 283897 -480 283953 240
rect 284495 -480 284551 240
rect 285093 -480 285149 240
rect 285691 -480 285747 240
rect 286289 -480 286345 240
rect 286841 -480 286897 240
rect 287439 -480 287495 240
rect 288037 -480 288093 240
rect 288635 -480 288691 240
rect 289233 -480 289289 240
rect 289887 -480 289943 240
rect 290485 -480 290541 240
rect 291083 -480 291139 240
rect 291681 -480 291737 240
<< metal3 >>
rect -480 348610 240 348730
rect 291760 348542 292480 348662
rect -480 342082 240 342202
rect 291760 341878 292480 341998
rect -480 335554 240 335674
rect 291760 335282 292480 335402
rect -480 329026 240 329146
rect 291760 328618 292480 328738
rect -480 322498 240 322618
rect 291760 321954 292480 322074
rect -480 315970 240 316090
rect 291760 315358 292480 315478
rect -480 309510 240 309630
rect 291760 308694 292480 308814
rect -480 302982 240 303102
rect 291760 302030 292480 302150
rect -480 296454 240 296574
rect 291760 295434 292480 295554
rect -480 289926 240 290046
rect 291760 288770 292480 288890
rect -480 283398 240 283518
rect 291760 282106 292480 282226
rect -480 276870 240 276990
rect 291760 275510 292480 275630
rect -480 270342 240 270462
rect 291760 268846 292480 268966
rect -480 263882 240 264002
rect 291760 262182 292480 262302
rect -480 257354 240 257474
rect 291760 255586 292480 255706
rect -480 250826 240 250946
rect 291760 248922 292480 249042
rect -480 244298 240 244418
rect 291760 242258 292480 242378
rect -480 237770 240 237890
rect 291760 235662 292480 235782
rect -480 231242 240 231362
rect 291760 228998 292480 229118
rect -480 224714 240 224834
rect 291760 222334 292480 222454
rect -480 218254 240 218374
rect 291760 215738 292480 215858
rect -480 211726 240 211846
rect 291760 209074 292480 209194
rect -480 205198 240 205318
rect 291760 202410 292480 202530
rect -480 198670 240 198790
rect 291760 195814 292480 195934
rect -480 192142 240 192262
rect 291760 189150 292480 189270
rect -480 185614 240 185734
rect 291760 182486 292480 182606
rect -480 179154 240 179274
rect 291760 175890 292480 176010
rect -480 172626 240 172746
rect 291760 169226 292480 169346
rect -480 166098 240 166218
rect 291760 162562 292480 162682
rect -480 159570 240 159690
rect 291760 155966 292480 156086
rect -480 153042 240 153162
rect 291760 149302 292480 149422
rect -480 146514 240 146634
rect 291760 142638 292480 142758
rect -480 139986 240 140106
rect 291760 136042 292480 136162
rect -480 133526 240 133646
rect 291760 129378 292480 129498
rect -480 126998 240 127118
rect 291760 122714 292480 122834
rect -480 120470 240 120590
rect 291760 116118 292480 116238
rect -480 113942 240 114062
rect 291760 109454 292480 109574
rect -480 107414 240 107534
rect 291760 102790 292480 102910
rect -480 100886 240 101006
rect 291760 96194 292480 96314
rect -480 94358 240 94478
rect 291760 89530 292480 89650
rect -480 87898 240 88018
rect 291760 82866 292480 82986
rect -480 81370 240 81490
rect 291760 76270 292480 76390
rect -480 74842 240 74962
rect 291760 69606 292480 69726
rect -480 68314 240 68434
rect 291760 62942 292480 63062
rect -480 61786 240 61906
rect 291760 56346 292480 56466
rect -480 55258 240 55378
rect 291760 49682 292480 49802
rect -480 48730 240 48850
rect 291760 43018 292480 43138
rect -480 42270 240 42390
rect 291760 36422 292480 36542
rect -480 35742 240 35862
rect 291760 29758 292480 29878
rect -480 29214 240 29334
rect 291760 23094 292480 23214
rect -480 22686 240 22806
rect 291760 16498 292480 16618
rect -480 16158 240 16278
rect 291760 9834 292480 9954
rect -480 9630 240 9750
rect -480 3170 240 3290
rect 291760 3238 292480 3358
<< metal4 >>
rect -4363 355779 -4053 355795
rect -4363 355661 -4347 355779
rect -4229 355661 -4187 355779
rect -4069 355661 -4053 355779
rect -4363 355619 -4053 355661
rect -4363 355501 -4347 355619
rect -4229 355501 -4187 355619
rect -4069 355501 -4053 355619
rect -4363 -3533 -4053 355501
rect 296015 355779 296325 355795
rect 296015 355661 296031 355779
rect 296149 355661 296191 355779
rect 296309 355661 296325 355779
rect 296015 355619 296325 355661
rect 296015 355501 296031 355619
rect 296149 355501 296191 355619
rect 296309 355501 296325 355619
rect -3883 355299 -3573 355315
rect -3883 355181 -3867 355299
rect -3749 355181 -3707 355299
rect -3589 355181 -3573 355299
rect -3883 355139 -3573 355181
rect -3883 355021 -3867 355139
rect -3749 355021 -3707 355139
rect -3589 355021 -3573 355139
rect -3883 -3053 -3573 355021
rect 295535 355299 295845 355315
rect 295535 355181 295551 355299
rect 295669 355181 295711 355299
rect 295829 355181 295845 355299
rect 295535 355139 295845 355181
rect 295535 355021 295551 355139
rect 295669 355021 295711 355139
rect 295829 355021 295845 355139
rect -3403 354819 -3093 354835
rect -3403 354701 -3387 354819
rect -3269 354701 -3227 354819
rect -3109 354701 -3093 354819
rect -3403 354659 -3093 354701
rect -3403 354541 -3387 354659
rect -3269 354541 -3227 354659
rect -3109 354541 -3093 354659
rect -3403 -2573 -3093 354541
rect 295055 354819 295365 354835
rect 295055 354701 295071 354819
rect 295189 354701 295231 354819
rect 295349 354701 295365 354819
rect 295055 354659 295365 354701
rect 295055 354541 295071 354659
rect 295189 354541 295231 354659
rect 295349 354541 295365 354659
rect -2923 354339 -2613 354355
rect -2923 354221 -2907 354339
rect -2789 354221 -2747 354339
rect -2629 354221 -2613 354339
rect -2923 354179 -2613 354221
rect -2923 354061 -2907 354179
rect -2789 354061 -2747 354179
rect -2629 354061 -2613 354179
rect -2923 -2093 -2613 354061
rect 294575 354339 294885 354355
rect 294575 354221 294591 354339
rect 294709 354221 294751 354339
rect 294869 354221 294885 354339
rect 294575 354179 294885 354221
rect 294575 354061 294591 354179
rect 294709 354061 294751 354179
rect 294869 354061 294885 354179
rect -2443 353859 -2133 353875
rect -2443 353741 -2427 353859
rect -2309 353741 -2267 353859
rect -2149 353741 -2133 353859
rect -2443 353699 -2133 353741
rect -2443 353581 -2427 353699
rect -2309 353581 -2267 353699
rect -2149 353581 -2133 353699
rect -2443 -1613 -2133 353581
rect 294095 353859 294405 353875
rect 294095 353741 294111 353859
rect 294229 353741 294271 353859
rect 294389 353741 294405 353859
rect 294095 353699 294405 353741
rect 294095 353581 294111 353699
rect 294229 353581 294271 353699
rect 294389 353581 294405 353699
rect -1963 353379 -1653 353395
rect -1963 353261 -1947 353379
rect -1829 353261 -1787 353379
rect -1669 353261 -1653 353379
rect -1963 353219 -1653 353261
rect -1963 353101 -1947 353219
rect -1829 353101 -1787 353219
rect -1669 353101 -1653 353219
rect -1963 -1133 -1653 353101
rect 293615 353379 293925 353395
rect 293615 353261 293631 353379
rect 293749 353261 293791 353379
rect 293909 353261 293925 353379
rect 293615 353219 293925 353261
rect 293615 353101 293631 353219
rect 293749 353101 293791 353219
rect 293909 353101 293925 353219
rect -1483 352899 -1173 352915
rect -1483 352781 -1467 352899
rect -1349 352781 -1307 352899
rect -1189 352781 -1173 352899
rect -1483 352739 -1173 352781
rect -1483 352621 -1467 352739
rect -1349 352621 -1307 352739
rect -1189 352621 -1173 352739
rect -1483 -653 -1173 352621
rect 293135 352899 293445 352915
rect 293135 352781 293151 352899
rect 293269 352781 293311 352899
rect 293429 352781 293445 352899
rect 293135 352739 293445 352781
rect 293135 352621 293151 352739
rect 293269 352621 293311 352739
rect 293429 352621 293445 352739
rect -1003 352419 -693 352435
rect -1003 352301 -987 352419
rect -869 352301 -827 352419
rect -709 352301 -693 352419
rect -1003 352259 -693 352301
rect -1003 352141 -987 352259
rect -869 352141 -827 352259
rect -709 352141 -693 352259
rect -1003 -173 -693 352141
rect -1003 -291 -987 -173
rect -869 -291 -827 -173
rect -709 -291 -693 -173
rect -1003 -333 -693 -291
rect -1003 -451 -987 -333
rect -869 -451 -827 -333
rect -709 -451 -693 -333
rect -1003 -467 -693 -451
rect 292655 352419 292965 352435
rect 292655 352301 292671 352419
rect 292789 352301 292831 352419
rect 292949 352301 292965 352419
rect 292655 352259 292965 352301
rect 292655 352141 292671 352259
rect 292789 352141 292831 352259
rect 292949 352141 292965 352259
rect 292655 -173 292965 352141
rect 292655 -291 292671 -173
rect 292789 -291 292831 -173
rect 292949 -291 292965 -173
rect 292655 -333 292965 -291
rect 292655 -451 292671 -333
rect 292789 -451 292831 -333
rect 292949 -451 292965 -333
rect 292655 -467 292965 -451
rect -1483 -771 -1467 -653
rect -1349 -771 -1307 -653
rect -1189 -771 -1173 -653
rect -1483 -813 -1173 -771
rect -1483 -931 -1467 -813
rect -1349 -931 -1307 -813
rect -1189 -931 -1173 -813
rect -1483 -947 -1173 -931
rect 293135 -653 293445 352621
rect 293135 -771 293151 -653
rect 293269 -771 293311 -653
rect 293429 -771 293445 -653
rect 293135 -813 293445 -771
rect 293135 -931 293151 -813
rect 293269 -931 293311 -813
rect 293429 -931 293445 -813
rect 293135 -947 293445 -931
rect -1963 -1251 -1947 -1133
rect -1829 -1251 -1787 -1133
rect -1669 -1251 -1653 -1133
rect -1963 -1293 -1653 -1251
rect -1963 -1411 -1947 -1293
rect -1829 -1411 -1787 -1293
rect -1669 -1411 -1653 -1293
rect -1963 -1427 -1653 -1411
rect 293615 -1133 293925 353101
rect 293615 -1251 293631 -1133
rect 293749 -1251 293791 -1133
rect 293909 -1251 293925 -1133
rect 293615 -1293 293925 -1251
rect 293615 -1411 293631 -1293
rect 293749 -1411 293791 -1293
rect 293909 -1411 293925 -1293
rect 293615 -1427 293925 -1411
rect -2443 -1731 -2427 -1613
rect -2309 -1731 -2267 -1613
rect -2149 -1731 -2133 -1613
rect -2443 -1773 -2133 -1731
rect -2443 -1891 -2427 -1773
rect -2309 -1891 -2267 -1773
rect -2149 -1891 -2133 -1773
rect -2443 -1907 -2133 -1891
rect 294095 -1613 294405 353581
rect 294095 -1731 294111 -1613
rect 294229 -1731 294271 -1613
rect 294389 -1731 294405 -1613
rect 294095 -1773 294405 -1731
rect 294095 -1891 294111 -1773
rect 294229 -1891 294271 -1773
rect 294389 -1891 294405 -1773
rect 294095 -1907 294405 -1891
rect -2923 -2211 -2907 -2093
rect -2789 -2211 -2747 -2093
rect -2629 -2211 -2613 -2093
rect -2923 -2253 -2613 -2211
rect -2923 -2371 -2907 -2253
rect -2789 -2371 -2747 -2253
rect -2629 -2371 -2613 -2253
rect -2923 -2387 -2613 -2371
rect 294575 -2093 294885 354061
rect 294575 -2211 294591 -2093
rect 294709 -2211 294751 -2093
rect 294869 -2211 294885 -2093
rect 294575 -2253 294885 -2211
rect 294575 -2371 294591 -2253
rect 294709 -2371 294751 -2253
rect 294869 -2371 294885 -2253
rect 294575 -2387 294885 -2371
rect -3403 -2691 -3387 -2573
rect -3269 -2691 -3227 -2573
rect -3109 -2691 -3093 -2573
rect -3403 -2733 -3093 -2691
rect -3403 -2851 -3387 -2733
rect -3269 -2851 -3227 -2733
rect -3109 -2851 -3093 -2733
rect -3403 -2867 -3093 -2851
rect 295055 -2573 295365 354541
rect 295055 -2691 295071 -2573
rect 295189 -2691 295231 -2573
rect 295349 -2691 295365 -2573
rect 295055 -2733 295365 -2691
rect 295055 -2851 295071 -2733
rect 295189 -2851 295231 -2733
rect 295349 -2851 295365 -2733
rect 295055 -2867 295365 -2851
rect -3883 -3171 -3867 -3053
rect -3749 -3171 -3707 -3053
rect -3589 -3171 -3573 -3053
rect -3883 -3213 -3573 -3171
rect -3883 -3331 -3867 -3213
rect -3749 -3331 -3707 -3213
rect -3589 -3331 -3573 -3213
rect -3883 -3347 -3573 -3331
rect 295535 -3053 295845 355021
rect 295535 -3171 295551 -3053
rect 295669 -3171 295711 -3053
rect 295829 -3171 295845 -3053
rect 295535 -3213 295845 -3171
rect 295535 -3331 295551 -3213
rect 295669 -3331 295711 -3213
rect 295829 -3331 295845 -3213
rect 295535 -3347 295845 -3331
rect -4363 -3651 -4347 -3533
rect -4229 -3651 -4187 -3533
rect -4069 -3651 -4053 -3533
rect -4363 -3693 -4053 -3651
rect -4363 -3811 -4347 -3693
rect -4229 -3811 -4187 -3693
rect -4069 -3811 -4053 -3693
rect -4363 -3827 -4053 -3811
rect 296015 -3533 296325 355501
rect 296015 -3651 296031 -3533
rect 296149 -3651 296191 -3533
rect 296309 -3651 296325 -3533
rect 296015 -3693 296325 -3651
rect 296015 -3811 296031 -3693
rect 296149 -3811 296191 -3693
rect 296309 -3811 296325 -3693
rect 296015 -3827 296325 -3811
<< via4 >>
rect -4347 355661 -4229 355779
rect -4187 355661 -4069 355779
rect -4347 355501 -4229 355619
rect -4187 355501 -4069 355619
rect 296031 355661 296149 355779
rect 296191 355661 296309 355779
rect 296031 355501 296149 355619
rect 296191 355501 296309 355619
rect -3867 355181 -3749 355299
rect -3707 355181 -3589 355299
rect -3867 355021 -3749 355139
rect -3707 355021 -3589 355139
rect 295551 355181 295669 355299
rect 295711 355181 295829 355299
rect 295551 355021 295669 355139
rect 295711 355021 295829 355139
rect -3387 354701 -3269 354819
rect -3227 354701 -3109 354819
rect -3387 354541 -3269 354659
rect -3227 354541 -3109 354659
rect 295071 354701 295189 354819
rect 295231 354701 295349 354819
rect 295071 354541 295189 354659
rect 295231 354541 295349 354659
rect -2907 354221 -2789 354339
rect -2747 354221 -2629 354339
rect -2907 354061 -2789 354179
rect -2747 354061 -2629 354179
rect 294591 354221 294709 354339
rect 294751 354221 294869 354339
rect 294591 354061 294709 354179
rect 294751 354061 294869 354179
rect -2427 353741 -2309 353859
rect -2267 353741 -2149 353859
rect -2427 353581 -2309 353699
rect -2267 353581 -2149 353699
rect 294111 353741 294229 353859
rect 294271 353741 294389 353859
rect 294111 353581 294229 353699
rect 294271 353581 294389 353699
rect -1947 353261 -1829 353379
rect -1787 353261 -1669 353379
rect -1947 353101 -1829 353219
rect -1787 353101 -1669 353219
rect 293631 353261 293749 353379
rect 293791 353261 293909 353379
rect 293631 353101 293749 353219
rect 293791 353101 293909 353219
rect -1467 352781 -1349 352899
rect -1307 352781 -1189 352899
rect -1467 352621 -1349 352739
rect -1307 352621 -1189 352739
rect 293151 352781 293269 352899
rect 293311 352781 293429 352899
rect 293151 352621 293269 352739
rect 293311 352621 293429 352739
rect -987 352301 -869 352419
rect -827 352301 -709 352419
rect -987 352141 -869 352259
rect -827 352141 -709 352259
rect -987 -291 -869 -173
rect -827 -291 -709 -173
rect -987 -451 -869 -333
rect -827 -451 -709 -333
rect 292671 352301 292789 352419
rect 292831 352301 292949 352419
rect 292671 352141 292789 352259
rect 292831 352141 292949 352259
rect 292671 -291 292789 -173
rect 292831 -291 292949 -173
rect 292671 -451 292789 -333
rect 292831 -451 292949 -333
rect -1467 -771 -1349 -653
rect -1307 -771 -1189 -653
rect -1467 -931 -1349 -813
rect -1307 -931 -1189 -813
rect 293151 -771 293269 -653
rect 293311 -771 293429 -653
rect 293151 -931 293269 -813
rect 293311 -931 293429 -813
rect -1947 -1251 -1829 -1133
rect -1787 -1251 -1669 -1133
rect -1947 -1411 -1829 -1293
rect -1787 -1411 -1669 -1293
rect 293631 -1251 293749 -1133
rect 293791 -1251 293909 -1133
rect 293631 -1411 293749 -1293
rect 293791 -1411 293909 -1293
rect -2427 -1731 -2309 -1613
rect -2267 -1731 -2149 -1613
rect -2427 -1891 -2309 -1773
rect -2267 -1891 -2149 -1773
rect 294111 -1731 294229 -1613
rect 294271 -1731 294389 -1613
rect 294111 -1891 294229 -1773
rect 294271 -1891 294389 -1773
rect -2907 -2211 -2789 -2093
rect -2747 -2211 -2629 -2093
rect -2907 -2371 -2789 -2253
rect -2747 -2371 -2629 -2253
rect 294591 -2211 294709 -2093
rect 294751 -2211 294869 -2093
rect 294591 -2371 294709 -2253
rect 294751 -2371 294869 -2253
rect -3387 -2691 -3269 -2573
rect -3227 -2691 -3109 -2573
rect -3387 -2851 -3269 -2733
rect -3227 -2851 -3109 -2733
rect 295071 -2691 295189 -2573
rect 295231 -2691 295349 -2573
rect 295071 -2851 295189 -2733
rect 295231 -2851 295349 -2733
rect -3867 -3171 -3749 -3053
rect -3707 -3171 -3589 -3053
rect -3867 -3331 -3749 -3213
rect -3707 -3331 -3589 -3213
rect 295551 -3171 295669 -3053
rect 295711 -3171 295829 -3053
rect 295551 -3331 295669 -3213
rect 295711 -3331 295829 -3213
rect -4347 -3651 -4229 -3533
rect -4187 -3651 -4069 -3533
rect -4347 -3811 -4229 -3693
rect -4187 -3811 -4069 -3693
rect 296031 -3651 296149 -3533
rect 296191 -3651 296309 -3533
rect 296031 -3811 296149 -3693
rect 296191 -3811 296309 -3693
<< metal5 >>
rect -4363 355779 296325 355795
rect -4363 355661 -4347 355779
rect -4229 355661 -4187 355779
rect -4069 355661 296031 355779
rect 296149 355661 296191 355779
rect 296309 355661 296325 355779
rect -4363 355619 296325 355661
rect -4363 355501 -4347 355619
rect -4229 355501 -4187 355619
rect -4069 355501 296031 355619
rect 296149 355501 296191 355619
rect 296309 355501 296325 355619
rect -4363 355485 296325 355501
rect -3883 355299 295845 355315
rect -3883 355181 -3867 355299
rect -3749 355181 -3707 355299
rect -3589 355181 295551 355299
rect 295669 355181 295711 355299
rect 295829 355181 295845 355299
rect -3883 355139 295845 355181
rect -3883 355021 -3867 355139
rect -3749 355021 -3707 355139
rect -3589 355021 295551 355139
rect 295669 355021 295711 355139
rect 295829 355021 295845 355139
rect -3883 355005 295845 355021
rect -3403 354819 295365 354835
rect -3403 354701 -3387 354819
rect -3269 354701 -3227 354819
rect -3109 354701 295071 354819
rect 295189 354701 295231 354819
rect 295349 354701 295365 354819
rect -3403 354659 295365 354701
rect -3403 354541 -3387 354659
rect -3269 354541 -3227 354659
rect -3109 354541 295071 354659
rect 295189 354541 295231 354659
rect 295349 354541 295365 354659
rect -3403 354525 295365 354541
rect -2923 354339 294885 354355
rect -2923 354221 -2907 354339
rect -2789 354221 -2747 354339
rect -2629 354221 294591 354339
rect 294709 354221 294751 354339
rect 294869 354221 294885 354339
rect -2923 354179 294885 354221
rect -2923 354061 -2907 354179
rect -2789 354061 -2747 354179
rect -2629 354061 294591 354179
rect 294709 354061 294751 354179
rect 294869 354061 294885 354179
rect -2923 354045 294885 354061
rect -2443 353859 294405 353875
rect -2443 353741 -2427 353859
rect -2309 353741 -2267 353859
rect -2149 353741 294111 353859
rect 294229 353741 294271 353859
rect 294389 353741 294405 353859
rect -2443 353699 294405 353741
rect -2443 353581 -2427 353699
rect -2309 353581 -2267 353699
rect -2149 353581 294111 353699
rect 294229 353581 294271 353699
rect 294389 353581 294405 353699
rect -2443 353565 294405 353581
rect -1963 353379 293925 353395
rect -1963 353261 -1947 353379
rect -1829 353261 -1787 353379
rect -1669 353261 293631 353379
rect 293749 353261 293791 353379
rect 293909 353261 293925 353379
rect -1963 353219 293925 353261
rect -1963 353101 -1947 353219
rect -1829 353101 -1787 353219
rect -1669 353101 293631 353219
rect 293749 353101 293791 353219
rect 293909 353101 293925 353219
rect -1963 353085 293925 353101
rect -1483 352899 293445 352915
rect -1483 352781 -1467 352899
rect -1349 352781 -1307 352899
rect -1189 352781 293151 352899
rect 293269 352781 293311 352899
rect 293429 352781 293445 352899
rect -1483 352739 293445 352781
rect -1483 352621 -1467 352739
rect -1349 352621 -1307 352739
rect -1189 352621 293151 352739
rect 293269 352621 293311 352739
rect 293429 352621 293445 352739
rect -1483 352605 293445 352621
rect -1003 352419 292965 352435
rect -1003 352301 -987 352419
rect -869 352301 -827 352419
rect -709 352301 292671 352419
rect 292789 352301 292831 352419
rect 292949 352301 292965 352419
rect -1003 352259 292965 352301
rect -1003 352141 -987 352259
rect -869 352141 -827 352259
rect -709 352141 292671 352259
rect 292789 352141 292831 352259
rect 292949 352141 292965 352259
rect -1003 352125 292965 352141
rect -1003 -173 292965 -157
rect -1003 -291 -987 -173
rect -869 -291 -827 -173
rect -709 -291 292671 -173
rect 292789 -291 292831 -173
rect 292949 -291 292965 -173
rect -1003 -333 292965 -291
rect -1003 -451 -987 -333
rect -869 -451 -827 -333
rect -709 -451 292671 -333
rect 292789 -451 292831 -333
rect 292949 -451 292965 -333
rect -1003 -467 292965 -451
rect -1483 -653 293445 -637
rect -1483 -771 -1467 -653
rect -1349 -771 -1307 -653
rect -1189 -771 293151 -653
rect 293269 -771 293311 -653
rect 293429 -771 293445 -653
rect -1483 -813 293445 -771
rect -1483 -931 -1467 -813
rect -1349 -931 -1307 -813
rect -1189 -931 293151 -813
rect 293269 -931 293311 -813
rect 293429 -931 293445 -813
rect -1483 -947 293445 -931
rect -1963 -1133 293925 -1117
rect -1963 -1251 -1947 -1133
rect -1829 -1251 -1787 -1133
rect -1669 -1251 293631 -1133
rect 293749 -1251 293791 -1133
rect 293909 -1251 293925 -1133
rect -1963 -1293 293925 -1251
rect -1963 -1411 -1947 -1293
rect -1829 -1411 -1787 -1293
rect -1669 -1411 293631 -1293
rect 293749 -1411 293791 -1293
rect 293909 -1411 293925 -1293
rect -1963 -1427 293925 -1411
rect -2443 -1613 294405 -1597
rect -2443 -1731 -2427 -1613
rect -2309 -1731 -2267 -1613
rect -2149 -1731 294111 -1613
rect 294229 -1731 294271 -1613
rect 294389 -1731 294405 -1613
rect -2443 -1773 294405 -1731
rect -2443 -1891 -2427 -1773
rect -2309 -1891 -2267 -1773
rect -2149 -1891 294111 -1773
rect 294229 -1891 294271 -1773
rect 294389 -1891 294405 -1773
rect -2443 -1907 294405 -1891
rect -2923 -2093 294885 -2077
rect -2923 -2211 -2907 -2093
rect -2789 -2211 -2747 -2093
rect -2629 -2211 294591 -2093
rect 294709 -2211 294751 -2093
rect 294869 -2211 294885 -2093
rect -2923 -2253 294885 -2211
rect -2923 -2371 -2907 -2253
rect -2789 -2371 -2747 -2253
rect -2629 -2371 294591 -2253
rect 294709 -2371 294751 -2253
rect 294869 -2371 294885 -2253
rect -2923 -2387 294885 -2371
rect -3403 -2573 295365 -2557
rect -3403 -2691 -3387 -2573
rect -3269 -2691 -3227 -2573
rect -3109 -2691 295071 -2573
rect 295189 -2691 295231 -2573
rect 295349 -2691 295365 -2573
rect -3403 -2733 295365 -2691
rect -3403 -2851 -3387 -2733
rect -3269 -2851 -3227 -2733
rect -3109 -2851 295071 -2733
rect 295189 -2851 295231 -2733
rect 295349 -2851 295365 -2733
rect -3403 -2867 295365 -2851
rect -3883 -3053 295845 -3037
rect -3883 -3171 -3867 -3053
rect -3749 -3171 -3707 -3053
rect -3589 -3171 295551 -3053
rect 295669 -3171 295711 -3053
rect 295829 -3171 295845 -3053
rect -3883 -3213 295845 -3171
rect -3883 -3331 -3867 -3213
rect -3749 -3331 -3707 -3213
rect -3589 -3331 295551 -3213
rect 295669 -3331 295711 -3213
rect 295829 -3331 295845 -3213
rect -3883 -3347 295845 -3331
rect -4363 -3533 296325 -3517
rect -4363 -3651 -4347 -3533
rect -4229 -3651 -4187 -3533
rect -4069 -3651 296031 -3533
rect 296149 -3651 296191 -3533
rect 296309 -3651 296325 -3533
rect -4363 -3693 296325 -3651
rect -4363 -3811 -4347 -3693
rect -4229 -3811 -4187 -3693
rect -4069 -3811 296031 -3693
rect 296149 -3811 296191 -3693
rect 296309 -3811 296325 -3693
rect -4363 -3827 296325 -3811
<< labels >>
flabel metal3 s 291760 142638 292480 142758 0 FreeSans 400 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 223049 351760 223105 352480 0 FreeSans 400 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 190573 351760 190629 352480 0 FreeSans 400 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 158143 351760 158199 352480 0 FreeSans 400 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 125713 351760 125769 352480 0 FreeSans 400 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 93237 351760 93293 352480 0 FreeSans 400 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 60807 351760 60863 352480 0 FreeSans 400 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 28377 351760 28433 352480 0 FreeSans 400 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -480 348610 240 348730 0 FreeSans 400 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -480 322498 240 322618 0 FreeSans 400 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -480 296454 240 296574 0 FreeSans 400 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 291760 169226 292480 169346 0 FreeSans 400 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -480 270342 240 270462 0 FreeSans 400 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -480 244298 240 244418 0 FreeSans 400 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -480 218254 240 218374 0 FreeSans 400 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -480 192142 240 192262 0 FreeSans 400 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -480 166098 240 166218 0 FreeSans 400 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -480 139986 240 140106 0 FreeSans 400 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -480 113942 240 114062 0 FreeSans 400 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -480 87898 240 88018 0 FreeSans 400 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -480 61786 240 61906 0 FreeSans 400 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 291760 195814 292480 195934 0 FreeSans 400 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 291760 222334 292480 222454 0 FreeSans 400 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 291760 248922 292480 249042 0 FreeSans 400 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 291760 275510 292480 275630 0 FreeSans 400 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 291760 302030 292480 302150 0 FreeSans 400 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 291760 328618 292480 328738 0 FreeSans 400 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 287909 351760 287965 352480 0 FreeSans 400 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 255479 351760 255535 352480 0 FreeSans 400 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 291760 3238 292480 3358 0 FreeSans 400 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 291760 228998 292480 229118 0 FreeSans 400 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 291760 255586 292480 255706 0 FreeSans 400 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 291760 282106 292480 282226 0 FreeSans 400 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 291760 308694 292480 308814 0 FreeSans 400 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 291760 335282 292480 335402 0 FreeSans 400 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 279813 351760 279869 352480 0 FreeSans 400 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 247383 351760 247439 352480 0 FreeSans 400 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 214907 351760 214963 352480 0 FreeSans 400 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 182477 351760 182533 352480 0 FreeSans 400 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 150047 351760 150103 352480 0 FreeSans 400 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 291760 23094 292480 23214 0 FreeSans 400 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 117571 351760 117627 352480 0 FreeSans 400 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 85141 351760 85197 352480 0 FreeSans 400 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 52711 351760 52767 352480 0 FreeSans 400 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 20235 351760 20291 352480 0 FreeSans 400 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -480 342082 240 342202 0 FreeSans 400 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -480 315970 240 316090 0 FreeSans 400 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -480 289926 240 290046 0 FreeSans 400 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -480 263882 240 264002 0 FreeSans 400 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -480 237770 240 237890 0 FreeSans 400 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -480 211726 240 211846 0 FreeSans 400 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 291760 43018 292480 43138 0 FreeSans 400 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -480 185614 240 185734 0 FreeSans 400 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -480 159570 240 159690 0 FreeSans 400 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -480 133526 240 133646 0 FreeSans 400 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -480 107414 240 107534 0 FreeSans 400 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -480 81370 240 81490 0 FreeSans 400 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -480 55258 240 55378 0 FreeSans 400 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -480 35742 240 35862 0 FreeSans 400 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -480 16158 240 16278 0 FreeSans 400 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 291760 62942 292480 63062 0 FreeSans 400 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 291760 82866 292480 82986 0 FreeSans 400 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 291760 102790 292480 102910 0 FreeSans 400 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 291760 122714 292480 122834 0 FreeSans 400 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 291760 149302 292480 149422 0 FreeSans 400 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 291760 175890 292480 176010 0 FreeSans 400 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 291760 202410 292480 202530 0 FreeSans 400 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 291760 16498 292480 16618 0 FreeSans 400 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 291760 242258 292480 242378 0 FreeSans 400 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 291760 268846 292480 268966 0 FreeSans 400 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 291760 295434 292480 295554 0 FreeSans 400 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 291760 321954 292480 322074 0 FreeSans 400 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 291760 348542 292480 348662 0 FreeSans 400 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 263575 351760 263631 352480 0 FreeSans 400 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 231145 351760 231201 352480 0 FreeSans 400 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 198715 351760 198771 352480 0 FreeSans 400 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 166239 351760 166295 352480 0 FreeSans 400 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 133809 351760 133865 352480 0 FreeSans 400 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 291760 36422 292480 36542 0 FreeSans 400 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 101379 351760 101435 352480 0 FreeSans 400 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 68903 351760 68959 352480 0 FreeSans 400 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 36473 351760 36529 352480 0 FreeSans 400 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 4043 351760 4099 352480 0 FreeSans 400 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -480 329026 240 329146 0 FreeSans 400 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -480 302982 240 303102 0 FreeSans 400 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -480 276870 240 276990 0 FreeSans 400 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -480 250826 240 250946 0 FreeSans 400 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -480 224714 240 224834 0 FreeSans 400 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -480 198670 240 198790 0 FreeSans 400 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 291760 56346 292480 56466 0 FreeSans 400 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -480 172626 240 172746 0 FreeSans 400 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -480 146514 240 146634 0 FreeSans 400 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -480 120470 240 120590 0 FreeSans 400 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -480 94358 240 94478 0 FreeSans 400 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -480 68314 240 68434 0 FreeSans 400 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -480 42270 240 42390 0 FreeSans 400 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -480 22686 240 22806 0 FreeSans 400 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -480 3170 240 3290 0 FreeSans 400 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 291760 76270 292480 76390 0 FreeSans 400 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 291760 96194 292480 96314 0 FreeSans 400 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 291760 116118 292480 116238 0 FreeSans 400 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 291760 136042 292480 136162 0 FreeSans 400 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 291760 162562 292480 162682 0 FreeSans 400 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 291760 189150 292480 189270 0 FreeSans 400 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 291760 215738 292480 215858 0 FreeSans 400 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 291760 9834 292480 9954 0 FreeSans 400 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 291760 235662 292480 235782 0 FreeSans 400 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 291760 262182 292480 262302 0 FreeSans 400 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 291760 288770 292480 288890 0 FreeSans 400 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 291760 315358 292480 315478 0 FreeSans 400 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 291760 341878 292480 341998 0 FreeSans 400 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 271717 351760 271773 352480 0 FreeSans 400 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 239241 351760 239297 352480 0 FreeSans 400 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 206811 351760 206867 352480 0 FreeSans 400 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 174381 351760 174437 352480 0 FreeSans 400 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 141905 351760 141961 352480 0 FreeSans 400 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 291760 29758 292480 29878 0 FreeSans 400 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 109475 351760 109531 352480 0 FreeSans 400 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 77045 351760 77101 352480 0 FreeSans 400 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 44569 351760 44625 352480 0 FreeSans 400 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 12139 351760 12195 352480 0 FreeSans 400 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -480 335554 240 335674 0 FreeSans 400 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -480 309510 240 309630 0 FreeSans 400 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -480 283398 240 283518 0 FreeSans 400 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -480 257354 240 257474 0 FreeSans 400 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -480 231242 240 231362 0 FreeSans 400 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -480 205198 240 205318 0 FreeSans 400 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 291760 49682 292480 49802 0 FreeSans 400 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -480 179154 240 179274 0 FreeSans 400 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -480 153042 240 153162 0 FreeSans 400 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -480 126998 240 127118 0 FreeSans 400 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -480 100886 240 101006 0 FreeSans 400 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -480 74842 240 74962 0 FreeSans 400 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -480 48730 240 48850 0 FreeSans 400 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -480 29214 240 29334 0 FreeSans 400 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -480 9630 240 9750 0 FreeSans 400 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 291760 69606 292480 69726 0 FreeSans 400 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 291760 89530 292480 89650 0 FreeSans 400 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 291760 109454 292480 109574 0 FreeSans 400 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 291760 129378 292480 129498 0 FreeSans 400 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 291760 155966 292480 156086 0 FreeSans 400 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 291760 182486 292480 182606 0 FreeSans 400 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 291760 209074 292480 209194 0 FreeSans 400 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 289887 -480 289943 240 0 FreeSans 400 270 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 290485 -480 290541 240 0 FreeSans 400 270 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 291083 -480 291139 240 0 FreeSans 400 270 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 291681 -480 291737 240 0 FreeSans 400 270 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal5 -495 -3784 20 -3569 0 FreeSans 1600 0 0 0 vssa2
port 645 nsew
flabel metal5 -491 -3283 24 -3068 0 FreeSans 1600 0 0 0 vdda2
port 646 nsew
flabel metal5 -478 -2819 37 -2604 0 FreeSans 1600 0 0 0 vssa1
port 647 nsew
flabel metal5 -485 -2352 30 -2137 0 FreeSans 1600 0 0 0 vdda1
port 648 nsew
flabel metal5 -468 -1861 47 -1646 0 FreeSans 1600 0 0 0 vssd2
port 649 nsew
flabel metal5 -441 -1370 74 -1155 0 FreeSans 1600 0 0 0 vccd2
port 650 nsew
flabel metal5 -458 -903 57 -688 0 FreeSans 1600 0 0 0 vssd1
port 651 nsew
flabel metal5 -424 -429 91 -214 0 FreeSans 1600 0 0 0 vccd1
port 652 nsew
flabel metal2 s 227179 -480 227235 240 0 FreeSans 400 270 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 227731 -480 227787 240 0 FreeSans 400 270 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 228329 -480 228385 240 0 FreeSans 400 270 0 0 wb_ack_o
port 541 nsew signal tristate
flabel metal2 s 230721 -480 230777 240 0 FreeSans 400 270 0 0 wb_adr_i[0]
port 542 nsew signal input
flabel metal2 s 250823 -480 250879 240 0 FreeSans 400 270 0 0 wb_adr_i[10]
port 543 nsew signal input
flabel metal2 s 252571 -480 252627 240 0 FreeSans 400 270 0 0 wb_adr_i[11]
port 544 nsew signal input
flabel metal2 s 254365 -480 254421 240 0 FreeSans 400 270 0 0 wb_adr_i[12]
port 545 nsew signal input
flabel metal2 s 256113 -480 256169 240 0 FreeSans 400 270 0 0 wb_adr_i[13]
port 546 nsew signal input
flabel metal2 s 257907 -480 257963 240 0 FreeSans 400 270 0 0 wb_adr_i[14]
port 547 nsew signal input
flabel metal2 s 259655 -480 259711 240 0 FreeSans 400 270 0 0 wb_adr_i[15]
port 548 nsew signal input
flabel metal2 s 261449 -480 261505 240 0 FreeSans 400 270 0 0 wb_adr_i[16]
port 549 nsew signal input
flabel metal2 s 263197 -480 263253 240 0 FreeSans 400 270 0 0 wb_adr_i[17]
port 550 nsew signal input
flabel metal2 s 264991 -480 265047 240 0 FreeSans 400 270 0 0 wb_adr_i[18]
port 551 nsew signal input
flabel metal2 s 266739 -480 266795 240 0 FreeSans 400 270 0 0 wb_adr_i[19]
port 552 nsew signal input
flabel metal2 s 233067 -480 233123 240 0 FreeSans 400 270 0 0 wb_adr_i[1]
port 553 nsew signal input
flabel metal2 s 268533 -480 268589 240 0 FreeSans 400 270 0 0 wb_adr_i[20]
port 554 nsew signal input
flabel metal2 s 270327 -480 270383 240 0 FreeSans 400 270 0 0 wb_adr_i[21]
port 555 nsew signal input
flabel metal2 s 272075 -480 272131 240 0 FreeSans 400 270 0 0 wb_adr_i[22]
port 556 nsew signal input
flabel metal2 s 273869 -480 273925 240 0 FreeSans 400 270 0 0 wb_adr_i[23]
port 557 nsew signal input
flabel metal2 s 275617 -480 275673 240 0 FreeSans 400 270 0 0 wb_adr_i[24]
port 558 nsew signal input
flabel metal2 s 277411 -480 277467 240 0 FreeSans 400 270 0 0 wb_adr_i[25]
port 559 nsew signal input
flabel metal2 s 279159 -480 279215 240 0 FreeSans 400 270 0 0 wb_adr_i[26]
port 560 nsew signal input
flabel metal2 s 280953 -480 281009 240 0 FreeSans 400 270 0 0 wb_adr_i[27]
port 561 nsew signal input
flabel metal2 s 282701 -480 282757 240 0 FreeSans 400 270 0 0 wb_adr_i[28]
port 562 nsew signal input
flabel metal2 s 284495 -480 284551 240 0 FreeSans 400 270 0 0 wb_adr_i[29]
port 563 nsew signal input
flabel metal2 s 235413 -480 235469 240 0 FreeSans 400 270 0 0 wb_adr_i[2]
port 564 nsew signal input
flabel metal2 s 286289 -480 286345 240 0 FreeSans 400 270 0 0 wb_adr_i[30]
port 565 nsew signal input
flabel metal2 s 288037 -480 288093 240 0 FreeSans 400 270 0 0 wb_adr_i[31]
port 566 nsew signal input
flabel metal2 s 237805 -480 237861 240 0 FreeSans 400 270 0 0 wb_adr_i[3]
port 567 nsew signal input
flabel metal2 s 240151 -480 240207 240 0 FreeSans 400 270 0 0 wb_adr_i[4]
port 568 nsew signal input
flabel metal2 s 241945 -480 242001 240 0 FreeSans 400 270 0 0 wb_adr_i[5]
port 569 nsew signal input
flabel metal2 s 243693 -480 243749 240 0 FreeSans 400 270 0 0 wb_adr_i[6]
port 570 nsew signal input
flabel metal2 s 245487 -480 245543 240 0 FreeSans 400 270 0 0 wb_adr_i[7]
port 571 nsew signal input
flabel metal2 s 247235 -480 247291 240 0 FreeSans 400 270 0 0 wb_adr_i[8]
port 572 nsew signal input
flabel metal2 s 249029 -480 249085 240 0 FreeSans 400 270 0 0 wb_adr_i[9]
port 573 nsew signal input
flabel metal2 s 228927 -480 228983 240 0 FreeSans 400 270 0 0 wb_cyc_i
port 574 nsew signal input
flabel metal2 s 231273 -480 231329 240 0 FreeSans 400 270 0 0 wb_dat_i[0]
port 575 nsew signal input
flabel metal2 s 251375 -480 251431 240 0 FreeSans 400 270 0 0 wb_dat_i[10]
port 576 nsew signal input
flabel metal2 s 253169 -480 253225 240 0 FreeSans 400 270 0 0 wb_dat_i[11]
port 577 nsew signal input
flabel metal2 s 254917 -480 254973 240 0 FreeSans 400 270 0 0 wb_dat_i[12]
port 578 nsew signal input
flabel metal2 s 256711 -480 256767 240 0 FreeSans 400 270 0 0 wb_dat_i[13]
port 579 nsew signal input
flabel metal2 s 258505 -480 258561 240 0 FreeSans 400 270 0 0 wb_dat_i[14]
port 580 nsew signal input
flabel metal2 s 260253 -480 260309 240 0 FreeSans 400 270 0 0 wb_dat_i[15]
port 581 nsew signal input
flabel metal2 s 262047 -480 262103 240 0 FreeSans 400 270 0 0 wb_dat_i[16]
port 582 nsew signal input
flabel metal2 s 263795 -480 263851 240 0 FreeSans 400 270 0 0 wb_dat_i[17]
port 583 nsew signal input
flabel metal2 s 265589 -480 265645 240 0 FreeSans 400 270 0 0 wb_dat_i[18]
port 584 nsew signal input
flabel metal2 s 267337 -480 267393 240 0 FreeSans 400 270 0 0 wb_dat_i[19]
port 585 nsew signal input
flabel metal2 s 233665 -480 233721 240 0 FreeSans 400 270 0 0 wb_dat_i[1]
port 586 nsew signal input
flabel metal2 s 269131 -480 269187 240 0 FreeSans 400 270 0 0 wb_dat_i[20]
port 587 nsew signal input
flabel metal2 s 270879 -480 270935 240 0 FreeSans 400 270 0 0 wb_dat_i[21]
port 588 nsew signal input
flabel metal2 s 272673 -480 272729 240 0 FreeSans 400 270 0 0 wb_dat_i[22]
port 589 nsew signal input
flabel metal2 s 274467 -480 274523 240 0 FreeSans 400 270 0 0 wb_dat_i[23]
port 590 nsew signal input
flabel metal2 s 276215 -480 276271 240 0 FreeSans 400 270 0 0 wb_dat_i[24]
port 591 nsew signal input
flabel metal2 s 278009 -480 278065 240 0 FreeSans 400 270 0 0 wb_dat_i[25]
port 592 nsew signal input
flabel metal2 s 279757 -480 279813 240 0 FreeSans 400 270 0 0 wb_dat_i[26]
port 593 nsew signal input
flabel metal2 s 281551 -480 281607 240 0 FreeSans 400 270 0 0 wb_dat_i[27]
port 594 nsew signal input
flabel metal2 s 283299 -480 283355 240 0 FreeSans 400 270 0 0 wb_dat_i[28]
port 595 nsew signal input
flabel metal2 s 285093 -480 285149 240 0 FreeSans 400 270 0 0 wb_dat_i[29]
port 596 nsew signal input
flabel metal2 s 236011 -480 236067 240 0 FreeSans 400 270 0 0 wb_dat_i[2]
port 597 nsew signal input
flabel metal2 s 286841 -480 286897 240 0 FreeSans 400 270 0 0 wb_dat_i[30]
port 598 nsew signal input
flabel metal2 s 288635 -480 288691 240 0 FreeSans 400 270 0 0 wb_dat_i[31]
port 599 nsew signal input
flabel metal2 s 238403 -480 238459 240 0 FreeSans 400 270 0 0 wb_dat_i[3]
port 600 nsew signal input
flabel metal2 s 240749 -480 240805 240 0 FreeSans 400 270 0 0 wb_dat_i[4]
port 601 nsew signal input
flabel metal2 s 242543 -480 242599 240 0 FreeSans 400 270 0 0 wb_dat_i[5]
port 602 nsew signal input
flabel metal2 s 244291 -480 244347 240 0 FreeSans 400 270 0 0 wb_dat_i[6]
port 603 nsew signal input
flabel metal2 s 246085 -480 246141 240 0 FreeSans 400 270 0 0 wb_dat_i[7]
port 604 nsew signal input
flabel metal2 s 247833 -480 247889 240 0 FreeSans 400 270 0 0 wb_dat_i[8]
port 605 nsew signal input
flabel metal2 s 249627 -480 249683 240 0 FreeSans 400 270 0 0 wb_dat_i[9]
port 606 nsew signal input
flabel metal2 s 231871 -480 231927 240 0 FreeSans 400 270 0 0 wb_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 251973 -480 252029 240 0 FreeSans 400 270 0 0 wb_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 253767 -480 253823 240 0 FreeSans 400 270 0 0 wb_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 255515 -480 255571 240 0 FreeSans 400 270 0 0 wb_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 257309 -480 257365 240 0 FreeSans 400 270 0 0 wb_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 259057 -480 259113 240 0 FreeSans 400 270 0 0 wb_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 260851 -480 260907 240 0 FreeSans 400 270 0 0 wb_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 262645 -480 262701 240 0 FreeSans 400 270 0 0 wb_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 264393 -480 264449 240 0 FreeSans 400 270 0 0 wb_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 266187 -480 266243 240 0 FreeSans 400 270 0 0 wb_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 267935 -480 267991 240 0 FreeSans 400 270 0 0 wb_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 234263 -480 234319 240 0 FreeSans 400 270 0 0 wb_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 269729 -480 269785 240 0 FreeSans 400 270 0 0 wb_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 271477 -480 271533 240 0 FreeSans 400 270 0 0 wb_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 273271 -480 273327 240 0 FreeSans 400 270 0 0 wb_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 275019 -480 275075 240 0 FreeSans 400 270 0 0 wb_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 276813 -480 276869 240 0 FreeSans 400 270 0 0 wb_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 278561 -480 278617 240 0 FreeSans 400 270 0 0 wb_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 280355 -480 280411 240 0 FreeSans 400 270 0 0 wb_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 282149 -480 282205 240 0 FreeSans 400 270 0 0 wb_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 283897 -480 283953 240 0 FreeSans 400 270 0 0 wb_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 285691 -480 285747 240 0 FreeSans 400 270 0 0 wb_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 236609 -480 236665 240 0 FreeSans 400 270 0 0 wb_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 287439 -480 287495 240 0 FreeSans 400 270 0 0 wb_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 289233 -480 289289 240 0 FreeSans 400 270 0 0 wb_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 239001 -480 239057 240 0 FreeSans 400 270 0 0 wb_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 241347 -480 241403 240 0 FreeSans 400 270 0 0 wb_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 243095 -480 243151 240 0 FreeSans 400 270 0 0 wb_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 244889 -480 244945 240 0 FreeSans 400 270 0 0 wb_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 246683 -480 246739 240 0 FreeSans 400 270 0 0 wb_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 248431 -480 248487 240 0 FreeSans 400 270 0 0 wb_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 250225 -480 250281 240 0 FreeSans 400 270 0 0 wb_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 232469 -480 232525 240 0 FreeSans 400 270 0 0 wb_sel_i[0]
port 639 nsew signal input
flabel metal2 s 234861 -480 234917 240 0 FreeSans 400 270 0 0 wb_sel_i[1]
port 640 nsew signal input
flabel metal2 s 237207 -480 237263 240 0 FreeSans 400 270 0 0 wb_sel_i[2]
port 641 nsew signal input
flabel metal2 s 239553 -480 239609 240 0 FreeSans 400 270 0 0 wb_sel_i[3]
port 642 nsew signal input
flabel metal2 s 229525 -480 229581 240 0 FreeSans 400 270 0 0 wb_stb_i
port 643 nsew signal input
flabel metal2 s 230123 -480 230179 240 0 FreeSans 400 270 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 292000 352000
string LEFview true
<< end >>
