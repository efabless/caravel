magic
tech sky130A
magscale 1 2
timestamp 1680223961
<< checkpaint >>
rect 6151 8561 12163 9595
rect 6141 6135 12163 8561
rect 6141 5101 12153 6135
<< isosubstrate >>
rect -52 7354 7222 8450
rect -52 -62 11288 7354
<< nwell >>
rect 70 7344 6652 7795
rect 7401 6799 10893 7301
<< pwell >>
rect 463 6569 519 6579
rect 2635 5816 2853 6026
<< psubdiff >>
rect 38 8568 62 8640
rect 11170 8568 11194 8640
<< mvpsubdiff >>
rect 7438 7387 10856 7455
rect 3164 6326 3188 6728
rect 6990 6326 7014 6728
<< mvnsubdiff >>
rect 7467 7201 10827 7235
<< psubdiffcont >>
rect 62 8568 11170 8640
<< mvpsubdiffcont >>
rect 3188 6326 6990 6728
<< locali >>
rect -14 8552 26 8676
rect 11178 8552 11218 8676
rect 41 8275 183 8288
rect 41 8190 57 8275
rect 169 8190 183 8275
rect 41 7451 183 8190
rect 6891 8273 7134 8286
rect 6891 8112 6936 8273
rect 7117 8112 7134 8273
rect 6891 7455 7134 8112
rect 3043 7451 7134 7455
rect 41 7435 7134 7451
rect 41 7305 6927 7435
rect 35 6388 121 7179
rect 3043 7022 6927 7305
rect 7110 7322 7134 7435
rect 7110 7235 10827 7322
rect 7110 7201 7467 7235
rect 7110 7022 7134 7201
rect 3043 7005 7134 7022
rect 2907 6728 7134 6838
rect 2907 6388 3188 6728
rect 35 6326 3188 6388
rect 6990 6387 7134 6728
rect 6990 6326 10860 6387
rect 35 6320 3220 6326
rect 35 6318 505 6320
rect 35 6192 48 6318
rect 286 6192 505 6318
rect 35 6191 505 6192
rect 2951 6253 3220 6320
rect 6116 6253 10860 6326
rect 2951 6191 10860 6253
rect 35 6143 10860 6191
rect 35 5813 689 6143
rect 1006 5813 1393 6029
rect 1778 5813 2165 6029
rect 2550 6015 2937 6029
rect 2550 5829 2648 6015
rect 2840 5829 2937 6015
rect 2550 5813 2937 5829
rect 3322 5813 3709 6029
rect 4094 5813 4481 6029
rect 4866 5813 5253 6029
rect 5638 5813 6025 6029
rect 6410 5813 6797 6029
rect 7182 5813 7569 6029
rect 7954 5813 8341 6029
rect 8726 5813 9113 6029
rect 9498 5813 9885 6029
rect 10656 5813 10837 6029
rect 51 165 234 381
rect 619 165 1006 381
rect 1391 165 1778 381
rect 2163 165 2550 381
rect 2935 165 3322 381
rect 3707 165 4094 381
rect 4479 165 4866 381
rect 5251 165 5638 381
rect 6023 165 6410 381
rect 6795 165 7182 381
rect 7567 165 7954 381
rect 8339 165 8726 381
rect 9111 165 9498 381
rect 9883 165 10270 381
rect 10655 165 10835 381
<< viali >>
rect 26 8640 11178 8676
rect 26 8568 62 8640
rect 62 8568 11170 8640
rect 11170 8568 11178 8640
rect 26 8552 11178 8568
rect 57 8190 169 8275
rect 6936 8112 7117 8273
rect 9224 7854 9270 8060
rect 7604 7754 7807 7801
rect 9459 7754 9796 7801
rect 10785 7683 10819 7879
rect 6927 7022 7110 7435
rect 7870 6775 8128 6834
rect 3220 6326 6116 6693
rect 8439 6684 8506 6878
rect 8650 6720 8853 6767
rect 10270 6735 10316 6896
rect 48 6192 286 6318
rect 505 6191 2951 6320
rect 3220 6253 6116 6326
rect 2648 5829 2840 6015
rect 10202 5598 10340 6030
<< metal1 >>
rect -14 8676 11218 8684
rect -14 8552 26 8676
rect 11178 8552 11218 8676
rect -14 8544 11218 8552
rect 40 8275 7133 8286
rect 40 8190 57 8275
rect 169 8273 7133 8275
rect 169 8269 6936 8273
rect 624 8260 6936 8269
rect 624 8201 1026 8260
rect 169 8193 1026 8201
rect 7117 8209 7133 8273
rect 7284 8252 10841 8278
rect 169 8190 6936 8193
rect 40 8179 6936 8190
rect 218 8110 376 8127
rect 218 8038 436 8110
rect 709 8082 719 8144
rect 801 8129 818 8144
rect 801 8085 2498 8129
rect 2829 8085 2990 8129
rect 801 8082 818 8085
rect 218 8024 282 8038
rect 218 7641 313 8024
rect 375 7641 436 8038
rect 521 7788 567 8040
rect 627 7892 2821 8028
rect 502 7653 2537 7788
rect 218 7568 436 7641
rect 521 7597 567 7653
rect 709 7597 719 7606
rect 218 7554 375 7568
rect 218 7501 282 7554
rect 521 7553 719 7597
rect 709 7544 719 7553
rect 801 7597 818 7606
rect 2866 7597 2944 8085
rect 2993 7658 3300 7804
rect 801 7556 2990 7597
rect 801 7553 2922 7556
rect 801 7544 818 7553
rect 3360 7501 3433 8122
rect 3699 8082 3959 8128
rect 3486 7636 3556 8035
rect 218 7453 3433 7501
rect 218 7248 282 7453
rect 3497 7344 3556 7636
rect 185 7121 282 7248
rect 2382 7274 3556 7344
rect 3699 7642 3781 8082
rect 4283 8081 5747 8125
rect 6083 8081 6237 8125
rect 6910 8112 6936 8179
rect 7117 8112 7134 8209
rect 7284 8153 7318 8252
rect 10802 8153 10841 8252
rect 7284 8125 10841 8153
rect 3988 7805 4025 8041
rect 4109 7872 6071 8033
rect 3966 7645 5802 7805
rect 3699 7600 3773 7642
rect 3699 7554 3958 7600
rect 3988 7597 4025 7645
rect 6126 7597 6188 8081
rect 6249 7884 6537 8029
rect 6249 7690 6262 7884
rect 3699 7501 3773 7554
rect 3988 7553 6239 7597
rect 6612 7501 6674 8112
rect 3699 7453 6674 7501
rect 185 6969 263 7121
rect 2382 7074 2452 7274
rect 3699 7165 3773 7453
rect 2265 7047 2275 7074
rect 185 6573 282 6969
rect 25 6318 301 6326
rect 25 6192 48 6318
rect 286 6192 301 6318
rect 25 6185 301 6192
rect 25 5348 133 6185
rect 345 5944 399 7033
rect 781 7003 2275 7047
rect 2351 7047 2452 7074
rect 2767 7074 3773 7165
rect 2351 7003 2738 7047
rect 463 6745 634 6972
rect 2382 6952 2452 7003
rect 721 6815 2452 6952
rect 463 6579 2560 6745
rect 463 6569 634 6579
rect 505 6326 634 6569
rect 2629 6533 2693 7003
rect 2767 6949 2842 7074
rect 6752 7065 6823 8044
rect 6910 7435 7134 8112
rect 9218 8060 9276 8072
rect 9218 7854 9224 8060
rect 9270 8051 9276 8060
rect 10128 8051 10138 8053
rect 9270 8001 10138 8051
rect 9270 7854 9276 8001
rect 10128 7999 10138 8001
rect 10290 7999 10300 8053
rect 9218 7842 9276 7854
rect 10779 7879 10825 7891
rect 7592 7801 8339 7807
rect 7592 7754 7604 7801
rect 7807 7754 8339 7801
rect 7592 7748 8339 7754
rect 8519 7801 9808 7807
rect 8519 7754 9459 7801
rect 9796 7754 9808 7801
rect 8519 7748 9808 7754
rect 10779 7728 10785 7879
rect 10819 7728 10825 7879
rect 10743 7674 10753 7728
rect 10905 7674 10915 7728
rect 10779 7671 10825 7674
rect 2756 6573 2842 6949
rect 6407 7036 6825 7065
rect 3167 6819 6174 6842
rect 3167 6693 4331 6819
rect 5278 6693 6174 6819
rect 781 6489 2275 6533
rect 2265 6460 2275 6489
rect 2350 6460 2360 6533
rect 2585 6489 2739 6533
rect 3167 6326 3220 6693
rect 493 6320 3220 6326
rect 493 6191 505 6320
rect 2951 6253 3220 6320
rect 6116 6531 6174 6693
rect 6407 6623 6432 7036
rect 6803 6840 6825 7036
rect 6910 7022 6927 7435
rect 7110 7324 7134 7435
rect 7279 7543 10836 7570
rect 7279 7449 7306 7543
rect 8343 7449 8618 7543
rect 10649 7449 10836 7543
rect 7279 7417 10836 7449
rect 7110 7299 10832 7324
rect 7110 7124 7171 7299
rect 8320 7124 8602 7299
rect 10750 7124 10832 7299
rect 7110 7094 10832 7124
rect 7110 7022 7134 7094
rect 10516 7093 10832 7094
rect 6910 6994 7134 7022
rect 10264 6896 10322 6908
rect 8433 6878 8512 6890
rect 6803 6834 8140 6840
rect 6803 6775 7870 6834
rect 8128 6775 8140 6834
rect 6803 6769 8140 6775
rect 6803 6623 6825 6769
rect 8429 6684 8439 6878
rect 8506 6773 8516 6878
rect 8506 6767 8865 6773
rect 8506 6720 8650 6767
rect 8853 6720 8865 6767
rect 10264 6735 10270 6896
rect 10316 6834 10322 6896
rect 10316 6765 10507 6834
rect 10672 6765 10682 6834
rect 10316 6735 10322 6765
rect 10264 6723 10322 6735
rect 8506 6714 8865 6720
rect 8506 6684 8516 6714
rect 8433 6672 8512 6684
rect 6407 6600 6825 6623
rect 6116 6319 10827 6531
rect 6116 6253 6174 6319
rect 2951 6237 6174 6253
rect 10221 6260 10716 6270
rect 2951 6191 6175 6237
rect 493 6185 6175 6191
rect 10221 6187 10233 6260
rect 10700 6187 10716 6260
rect 10221 6176 10716 6187
rect 10221 6045 10315 6176
rect 10187 6030 10353 6045
rect 2635 6015 2853 6026
rect 2635 5944 2648 6015
rect 345 5890 2648 5944
rect 2635 5829 2648 5890
rect 2840 5829 2853 6015
rect 2635 5816 2853 5829
rect 10187 5598 10202 6030
rect 10340 5598 10353 6030
rect 10187 5582 10353 5598
rect 10805 5348 10867 6079
rect 25 4748 10867 5348
rect 25 4348 133 4748
rect 10805 4348 10867 4748
rect 25 3748 10867 4348
rect 25 3348 133 3748
rect 10805 3348 10867 3748
rect 25 2748 10867 3348
rect 25 2348 133 2748
rect 10805 2348 10867 2748
rect 25 1748 10867 2348
rect 25 1348 133 1748
rect 10805 1348 10867 1748
rect 25 748 10867 1348
rect 25 99 133 748
rect 10805 99 10867 748
rect 25 11 10867 99
<< via1 >>
rect 92 8568 11148 8640
rect 60 8201 169 8269
rect 169 8201 624 8269
rect 1026 8193 6936 8260
rect 6936 8193 7093 8260
rect 719 8082 801 8144
rect 719 7544 801 7606
rect 7318 8153 10802 8252
rect 2275 7003 2351 7074
rect 10138 7999 10290 8053
rect 8339 7748 8519 7807
rect 10753 7683 10785 7728
rect 10785 7683 10819 7728
rect 10819 7683 10905 7728
rect 10753 7674 10905 7683
rect 4331 6693 5278 6819
rect 2275 6460 2350 6533
rect 4331 6270 5278 6693
rect 6432 6623 6803 7036
rect 7306 7449 8343 7543
rect 8618 7449 10649 7543
rect 7171 7124 8320 7299
rect 8602 7124 10750 7299
rect 8439 6684 8506 6878
rect 10507 6765 10672 6834
rect 10233 6187 10700 6260
<< metal2 >>
rect -14 8640 11218 8684
rect -14 8568 92 8640
rect 11148 8568 11218 8640
rect -14 8544 11218 8568
rect 985 8286 7132 8287
rect 38 8269 7132 8286
rect 38 8201 60 8269
rect 624 8261 7132 8269
rect 38 8104 77 8201
rect 634 8187 886 8261
rect 7091 8260 7132 8261
rect 7093 8193 7132 8260
rect 634 8104 654 8187
rect 38 8061 654 8104
rect 719 8144 801 8154
rect 719 8072 801 8082
rect 866 8104 886 8187
rect 7091 8104 7132 8193
rect 7284 8252 10841 8278
rect 7284 8153 7318 8252
rect 10802 8153 10841 8252
rect 7284 8125 10841 8153
rect 729 7616 785 8072
rect 866 8060 7132 8104
rect 10138 8056 10290 8066
rect 10138 7986 10290 7996
rect 8339 7807 8519 7817
rect 8339 7738 8519 7748
rect 719 7606 801 7616
rect 719 7534 801 7544
rect 7279 7543 8374 7570
rect 7279 7449 7306 7543
rect 8343 7449 8374 7543
rect 7279 7417 8374 7449
rect 7141 7299 8355 7324
rect 7141 7124 7171 7299
rect 8320 7124 8355 7299
rect 7141 7094 8355 7124
rect 2275 7074 2351 7084
rect 2275 6993 2351 7003
rect 6407 7036 6825 7065
rect 2288 6543 2340 6993
rect 4308 6849 5298 6868
rect 2275 6533 2350 6543
rect 2275 6450 2350 6460
rect 4308 6270 4331 6849
rect 5278 6270 5298 6849
rect 6407 6623 6432 7036
rect 6803 6623 6825 7036
rect 8443 6888 8500 7738
rect 10753 7731 10905 7741
rect 10753 7661 10905 7671
rect 8588 7543 10667 7570
rect 8587 7449 8618 7543
rect 10649 7449 10667 7543
rect 8588 7417 10667 7449
rect 8567 7299 10798 7324
rect 8567 7124 8602 7299
rect 10750 7124 10798 7299
rect 8567 7094 10798 7124
rect 8439 6878 8506 6888
rect 8439 6674 8506 6684
rect 6407 6600 6825 6623
rect 4308 6249 5298 6270
rect 10221 6270 10431 7094
rect 10498 6765 10507 6834
rect 10672 6765 10757 6834
rect 10909 6765 10918 6834
rect 10221 6260 10716 6270
rect 10221 6187 10233 6260
rect 10700 6187 10716 6260
rect 10221 6176 10716 6187
<< via2 >>
rect 92 8568 11148 8640
rect 77 8201 624 8261
rect 624 8201 634 8261
rect 77 8104 634 8201
rect 886 8260 7091 8261
rect 886 8193 1026 8260
rect 1026 8193 7091 8260
rect 886 8104 7091 8193
rect 7318 8153 10802 8252
rect 10138 8053 10290 8056
rect 10138 7999 10290 8053
rect 10138 7996 10290 7999
rect 7306 7449 8343 7543
rect 4331 6819 5278 6849
rect 4331 6522 5278 6819
rect 6432 6623 6803 7036
rect 10753 7728 10905 7731
rect 10753 7674 10905 7728
rect 10753 7671 10905 7674
rect 8618 7449 10649 7543
rect 10757 6765 10909 6834
<< metal3 >>
rect -14 8674 11214 8684
rect -14 8640 7260 8674
rect 7724 8640 11214 8674
rect -14 8568 92 8640
rect 11148 8568 11214 8640
rect -14 8554 7260 8568
rect 7724 8554 11214 8568
rect -14 8438 11214 8554
rect 38 8261 7126 8283
rect 38 8244 77 8261
rect 634 8244 886 8261
rect 38 8000 73 8244
rect 7091 8104 7126 8261
rect 7284 8252 10841 8278
rect 7284 8153 7318 8252
rect 10802 8153 10841 8252
rect 7284 8125 10841 8153
rect 7073 8000 7126 8104
rect 38 7965 7126 8000
rect 10128 8056 10295 8064
rect 10128 7996 10138 8056
rect 10290 7996 10431 8056
rect 10128 7991 10295 7996
rect 10371 7916 10431 7996
rect 10371 7856 11343 7916
rect 10743 7731 10910 7739
rect 10743 7671 10753 7731
rect 10905 7671 10910 7731
rect 10743 7666 10910 7671
rect 7279 7543 10667 7570
rect 7279 7449 7306 7543
rect 10649 7449 10667 7543
rect 10792 7551 10852 7666
rect 10792 7491 11344 7551
rect 7279 7417 10667 7449
rect 4111 7277 5299 7317
rect 4111 6849 4350 7277
rect 5268 6849 5299 7277
rect 4111 6522 4331 6849
rect 5278 6522 5299 6849
rect 6408 7036 6825 7065
rect 6408 6623 6432 7036
rect 6803 6623 6825 7036
rect 10747 6834 10918 6840
rect 10747 6765 10757 6834
rect 10909 6765 11342 6834
rect 10747 6758 10918 6765
rect 6408 6600 6825 6623
rect 4111 6494 5299 6522
rect 4111 6251 4307 6494
<< via3 >>
rect 7260 8640 7724 8674
rect 7260 8568 7724 8640
rect 7260 8554 7724 8568
rect 73 8104 77 8244
rect 77 8104 634 8244
rect 634 8104 886 8244
rect 886 8104 7073 8244
rect 7928 8153 10802 8252
rect 73 8000 7073 8104
rect 7306 7449 8343 7543
rect 8343 7449 8618 7543
rect 8618 7449 10649 7543
rect 4350 6849 5268 7277
rect 4350 6558 5268 6849
rect 6432 6623 6803 7036
<< metal4 >>
rect 7248 8674 7736 8684
rect 7248 8554 7260 8674
rect 7724 8554 7736 8674
rect 38 8244 7126 8283
rect 38 8000 73 8244
rect 7073 8000 7126 8244
rect 38 7965 7126 8000
rect 7248 7655 7736 8554
rect 7918 8252 11180 8291
rect 7918 8153 7928 8252
rect 10802 8153 11180 8252
rect 7918 7962 11180 8153
rect 10843 7755 11178 7774
rect 38 7277 6984 7655
rect 38 7255 4350 7277
rect 3817 6558 4350 7255
rect 5268 7255 6984 7277
rect 7248 7543 10667 7655
rect 7248 7449 7306 7543
rect 10649 7449 10667 7543
rect 7248 7255 10667 7449
rect 5268 6558 5299 7255
rect 10843 7074 10879 7755
rect 6386 7036 10879 7074
rect 6386 6623 6432 7036
rect 6803 6623 10879 7036
rect 6386 6615 10879 6623
rect 11146 6615 11178 7755
rect 6386 6591 11178 6615
rect 3817 6522 5299 6558
rect 3817 51 4011 6522
rect 4101 51 4793 6251
<< via4 >>
rect 4350 6558 5268 7247
rect 10879 6615 11146 7755
<< metal5 >>
rect 10851 7755 11171 7779
rect 4313 7247 5299 7317
rect 4313 6558 4350 7247
rect 5268 6558 5299 7247
rect 4313 6494 5299 6558
rect 4507 6135 5299 6494
rect 10851 6615 10879 7755
rect 11146 6615 11171 7755
rect 10851 6242 11171 6615
use sky130_fd_pr__cap_mim_m3_1_WRT4AW  sky130_fd_pr__cap_mim_m3_1_WRT4AW_0 primitives
timestamp 1606502073
transform -1 0 7027 0 1 3151
box -3136 -3100 3136 3100
use sky130_fd_pr__cap_mim_m3_2_W5U4AW  sky130_fd_pr__cap_mim_m3_2_W5U4AW_0 primitives
timestamp 1606502073
transform 1 0 7970 0 1 3151
box -3179 -3101 3201 3101
use sky130_fd_pr__nfet_g5v0d10v5_PKVMTM  sky130_fd_pr__nfet_g5v0d10v5_PKVMTM_0 primitives
timestamp 1625577137
transform 1 0 2660 0 1 6770
box -308 -458 308 458
use sky130_fd_pr__nfet_g5v0d10v5_TGFUGS  sky130_fd_pr__nfet_g5v0d10v5_TGFUGS_0 primitives
timestamp 1606063140
transform 1 0 1515 0 1 6769
box -962 -458 962 458
use sky130_fd_pr__nfet_g5v0d10v5_ZK8HQC  sky130_fd_pr__nfet_g5v0d10v5_ZK8HQC_1 primitives
timestamp 1605994897
transform -1 0 371 0 1 6769
box -308 -458 308 458
use sky130_fd_pr__pfet_g5v0d10v5_3YBPVB  sky130_fd_pr__pfet_g5v0d10v5_3YBPVB_0 primitives
timestamp 1606063140
transform 1 0 3392 0 1 7841
box -338 -497 338 497
use sky130_fd_pr__pfet_g5v0d10v5_3YBPVB  sky130_fd_pr__pfet_g5v0d10v5_3YBPVB_1
timestamp 1606063140
transform 1 0 3878 0 1 7841
box -338 -497 338 497
use sky130_fd_pr__pfet_g5v0d10v5_3YBPVB  sky130_fd_pr__pfet_g5v0d10v5_3YBPVB_2
timestamp 1606063140
transform 1 0 6644 0 1 7841
box -338 -497 338 497
use sky130_fd_pr__pfet_g5v0d10v5_3YBPVB  sky130_fd_pr__pfet_g5v0d10v5_3YBPVB_3
timestamp 1606063140
transform 1 0 408 0 1 7841
box -338 -497 338 497
use sky130_fd_pr__pfet_g5v0d10v5_YEUEBV  sky130_fd_pr__pfet_g5v0d10v5_YEUEBV_0 primitives
timestamp 1606063140
transform 1 0 5018 0 1 7841
box -992 -497 992 497
use sky130_fd_pr__pfet_g5v0d10v5_YUHPBG  sky130_fd_pr__pfet_g5v0d10v5_YUHPBG_0 primitives
timestamp 1606063140
transform 1 0 2906 0 1 7841
box -338 -497 338 497
use sky130_fd_pr__pfet_g5v0d10v5_YUHPXE  sky130_fd_pr__pfet_g5v0d10v5_YUHPXE_0 primitives
timestamp 1606063140
transform 1 0 6158 0 1 7841
box -338 -497 338 497
use sky130_fd_pr__pfet_g5v0d10v5_ZEUEFZ  sky130_fd_pr__pfet_g5v0d10v5_ZEUEFZ_0 primitives
timestamp 1606063140
transform 1 0 1657 0 1 7841
box -1101 -497 1101 497
use sky130_fd_pr__res_xhigh_po_0p69_S5N9F3  sky130_fd_pr__res_xhigh_po_0p69_S5N9F3_0 primitives
timestamp 1606074388
transform 1 0 5446 0 1 3098
box -5446 -3098 5446 3098
use sky130_fd_sc_hvl__buf_8  sky130_fd_sc_hvl__buf_8_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1692890899
transform 1 0 8523 0 1 6404
box -66 -43 1986 897
use sky130_fd_sc_hvl__buf_8  sky130_fd_sc_hvl__buf_8_1
timestamp 1692890899
transform 1 0 7477 0 1 7438
box -66 -43 1986 897
use sky130_fd_sc_hvl__fill_4  sky130_fd_sc_hvl__fill_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1692890899
transform 1 0 10443 0 1 6404
box -66 -43 450 897
use sky130_fd_sc_hvl__inv_8  sky130_fd_sc_hvl__inv_8_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1692890899
transform 1 0 9397 0 1 7438
box -66 -43 1506 897
use sky130_fd_sc_hvl__schmittbuf_1  sky130_fd_sc_hvl__schmittbuf_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1692890899
transform 1 0 7467 0 1 6404
box -66 -43 1122 897
<< labels >>
flabel metal4 s 38 7965 73 8283 0 FreeSans 320 0 0 0 vdd3v3
port 0 nsew power bidirectional
flabel metal4 s 10974 7962 11180 8291 0 FreeSans 320 0 0 0 vdd1v8
port 1 nsew power bidirectional
flabel metal3 11189 7491 11344 7551 0 FreeSans 320 0 0 0 por_l
port 4 nsew signal output
flabel metal3 11188 7856 11343 7916 0 FreeSans 320 0 0 0 porb_l
port 5 nsew signal output
flabel metal3 10969 6765 11342 6834 0 FreeSans 320 0 0 0 porb_h
port 3 nsew signal output
flabel metal1 -14 8544 58 8684 0 FreeSans 800 0 0 0 vss1v8
port 6 nsew ground bidirectional
flabel metal4 s 38 7255 232 7655 0 FreeSans 320 0 0 0 vss3v3
port 2 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 11344 8338
string GDS_FILE ../gds/simple_por.gds
string GDS_START 0
string LEFclass BLOCK
<< end >>
