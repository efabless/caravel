VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mprj_logic_high
  CLASS BLOCK ;
  FOREIGN mprj_logic_high ;
  ORIGIN 0.000 0.000 ;
  SIZE 350.000 BY 22.000 ;
  PIN HI[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 3.000 19.680 ;
    END
  END HI[0]
  PIN HI[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 3.000 18.320 ;
    END
  END HI[100]
  PIN HI[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 3.000 16.960 ;
    END
  END HI[101]
  PIN HI[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 3.000 15.600 ;
    END
  END HI[102]
  PIN HI[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 3.000 14.240 ;
    END
  END HI[103]
  PIN HI[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 3.000 12.880 ;
    END
  END HI[104]
  PIN HI[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 3.000 11.520 ;
    END
  END HI[105]
  PIN HI[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 3.000 10.160 ;
    END
  END HI[106]
  PIN HI[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 3.000 8.800 ;
    END
  END HI[107]
  PIN HI[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 3.000 7.440 ;
    END
  END HI[108]
  PIN HI[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.480 3.000 6.080 ;
    END
  END HI[109]
  PIN HI[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 3.000 21.040 ;
    END
  END HI[10]
  PIN HI[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 3.000 4.720 ;
    END
  END HI[110]
  PIN HI[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 3.000 2.000 ;
    END
  END HI[111]
  PIN HI[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.040 3.000 0.640 ;
    END
  END HI[112]
  PIN HI[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 3.000 3.360 ;
    END
  END HI[113]
  PIN HI[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 70.470 19.000 70.750 22.000 ;
    END
  END HI[114]
  PIN HI[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 64.950 19.000 65.230 22.000 ;
    END
  END HI[115]
  PIN HI[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 69.090 19.000 69.370 22.000 ;
    END
  END HI[116]
  PIN HI[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 67.710 19.000 67.990 22.000 ;
    END
  END HI[117]
  PIN HI[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 47.010 19.000 47.290 22.000 ;
    END
  END HI[118]
  PIN HI[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 66.330 19.000 66.610 22.000 ;
    END
  END HI[119]
  PIN HI[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 62.190 19.000 62.470 22.000 ;
    END
  END HI[11]
  PIN HI[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 56.670 19.000 56.950 22.000 ;
    END
  END HI[120]
  PIN HI[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 63.570 19.000 63.850 22.000 ;
    END
  END HI[121]
  PIN HI[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 31.830 19.000 32.110 22.000 ;
    END
  END HI[122]
  PIN HI[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 60.810 19.000 61.090 22.000 ;
    END
  END HI[123]
  PIN HI[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 59.430 19.000 59.710 22.000 ;
    END
  END HI[124]
  PIN HI[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 58.050 19.000 58.330 22.000 ;
    END
  END HI[125]
  PIN HI[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 48.390 19.000 48.670 22.000 ;
    END
  END HI[126]
  PIN HI[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 55.290 19.000 55.570 22.000 ;
    END
  END HI[127]
  PIN HI[128]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 53.910 19.000 54.190 22.000 ;
    END
  END HI[128]
  PIN HI[129]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 52.530 19.000 52.810 22.000 ;
    END
  END HI[129]
  PIN HI[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 2.850 19.000 3.130 22.000 ;
    END
  END HI[12]
  PIN HI[130]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 51.150 19.000 51.430 22.000 ;
    END
  END HI[130]
  PIN HI[131]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 49.770 19.000 50.050 22.000 ;
    END
  END HI[131]
  PIN HI[132]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 38.730 19.000 39.010 22.000 ;
    END
  END HI[132]
  PIN HI[133]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 24.930 19.000 25.210 22.000 ;
    END
  END HI[133]
  PIN HI[134]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 45.630 19.000 45.910 22.000 ;
    END
  END HI[134]
  PIN HI[135]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 44.250 19.000 44.530 22.000 ;
    END
  END HI[135]
  PIN HI[136]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 42.870 19.000 43.150 22.000 ;
    END
  END HI[136]
  PIN HI[137]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 41.490 19.000 41.770 22.000 ;
    END
  END HI[137]
  PIN HI[138]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 40.110 19.000 40.390 22.000 ;
    END
  END HI[138]
  PIN HI[139]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 29.070 19.000 29.350 22.000 ;
    END
  END HI[139]
  PIN HI[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 71.850 19.000 72.130 22.000 ;
    END
  END HI[13]
  PIN HI[140]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 37.350 19.000 37.630 22.000 ;
    END
  END HI[140]
  PIN HI[141]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 35.970 19.000 36.250 22.000 ;
    END
  END HI[141]
  PIN HI[142]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 34.590 19.000 34.870 22.000 ;
    END
  END HI[142]
  PIN HI[143]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 33.210 19.000 33.490 22.000 ;
    END
  END HI[143]
  PIN HI[144]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 0.090 19.000 0.370 22.000 ;
    END
  END HI[144]
  PIN HI[145]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 30.450 19.000 30.730 22.000 ;
    END
  END HI[145]
  PIN HI[146]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 18.030 19.000 18.310 22.000 ;
    END
  END HI[146]
  PIN HI[147]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 27.690 19.000 27.970 22.000 ;
    END
  END HI[147]
  PIN HI[148]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 26.310 19.000 26.590 22.000 ;
    END
  END HI[148]
  PIN HI[149]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 1.470 19.000 1.750 22.000 ;
    END
  END HI[149]
  PIN HI[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 22.170 19.000 22.450 22.000 ;
    END
  END HI[14]
  PIN HI[150]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 23.550 19.000 23.830 22.000 ;
    END
  END HI[150]
  PIN HI[151]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 19.410 19.000 19.690 22.000 ;
    END
  END HI[151]
  PIN HI[152]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 20.790 19.000 21.070 22.000 ;
    END
  END HI[152]
  PIN HI[153]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 16.650 19.000 16.930 22.000 ;
    END
  END HI[153]
  PIN HI[154]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 5.610 19.000 5.890 22.000 ;
    END
  END HI[154]
  PIN HI[155]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 15.270 19.000 15.550 22.000 ;
    END
  END HI[155]
  PIN HI[156]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 13.890 19.000 14.170 22.000 ;
    END
  END HI[156]
  PIN HI[157]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 12.510 19.000 12.790 22.000 ;
    END
  END HI[157]
  PIN HI[158]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 11.130 19.000 11.410 22.000 ;
    END
  END HI[158]
  PIN HI[159]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 9.750 19.000 10.030 22.000 ;
    END
  END HI[159]
  PIN HI[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 73.230 19.000 73.510 22.000 ;
    END
  END HI[15]
  PIN HI[160]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 6.990 19.000 7.270 22.000 ;
    END
  END HI[160]
  PIN HI[161]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 8.370 19.000 8.650 22.000 ;
    END
  END HI[161]
  PIN HI[162]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 4.230 19.000 4.510 22.000 ;
    END
  END HI[162]
  PIN HI[163]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 3.000 ;
    END
  END HI[163]
  PIN HI[164]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 3.000 ;
    END
  END HI[164]
  PIN HI[165]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 3.000 ;
    END
  END HI[165]
  PIN HI[166]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 3.000 ;
    END
  END HI[166]
  PIN HI[167]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 3.000 ;
    END
  END HI[167]
  PIN HI[168]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 3.000 ;
    END
  END HI[168]
  PIN HI[169]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 3.000 ;
    END
  END HI[169]
  PIN HI[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 147.750 0.000 148.030 3.000 ;
    END
  END HI[16]
  PIN HI[170]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 227.790 0.000 228.070 3.000 ;
    END
  END HI[170]
  PIN HI[171]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 3.000 ;
    END
  END HI[171]
  PIN HI[172]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 149.130 0.000 149.410 3.000 ;
    END
  END HI[172]
  PIN HI[173]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 256.770 0.000 257.050 3.000 ;
    END
  END HI[173]
  PIN HI[174]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 51.150 0.000 51.430 3.000 ;
    END
  END HI[174]
  PIN HI[175]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 273.330 0.000 273.610 3.000 ;
    END
  END HI[175]
  PIN HI[176]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 95.310 0.000 95.590 3.000 ;
    END
  END HI[176]
  PIN HI[177]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 3.000 ;
    END
  END HI[177]
  PIN HI[178]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 3.000 ;
    END
  END HI[178]
  PIN HI[179]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 3.000 ;
    END
  END HI[179]
  PIN HI[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 3.000 ;
    END
  END HI[17]
  PIN HI[180]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 230.550 0.000 230.830 3.000 ;
    END
  END HI[180]
  PIN HI[181]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 3.000 ;
    END
  END HI[181]
  PIN HI[182]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 70.470 0.000 70.750 3.000 ;
    END
  END HI[182]
  PIN HI[183]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 3.000 ;
    END
  END HI[183]
  PIN HI[184]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 258.150 0.000 258.430 3.000 ;
    END
  END HI[184]
  PIN HI[185]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 3.000 ;
    END
  END HI[185]
  PIN HI[186]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 156.030 0.000 156.310 3.000 ;
    END
  END HI[186]
  PIN HI[187]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 3.000 ;
    END
  END HI[187]
  PIN HI[188]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 3.000 ;
    END
  END HI[188]
  PIN HI[189]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 3.000 ;
    END
  END HI[189]
  PIN HI[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 3.000 ;
    END
  END HI[18]
  PIN HI[190]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 84.270 0.000 84.550 3.000 ;
    END
  END HI[190]
  PIN HI[191]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 233.310 0.000 233.590 3.000 ;
    END
  END HI[191]
  PIN HI[192]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 3.000 ;
    END
  END HI[192]
  PIN HI[193]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 3.000 ;
    END
  END HI[193]
  PIN HI[194]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 259.530 0.000 259.810 3.000 ;
    END
  END HI[194]
  PIN HI[195]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 3.000 ;
    END
  END HI[195]
  PIN HI[196]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 3.000 ;
    END
  END HI[196]
  PIN HI[197]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 161.550 0.000 161.830 3.000 ;
    END
  END HI[197]
  PIN HI[198]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 3.000 ;
    END
  END HI[198]
  PIN HI[199]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 3.000 ;
    END
  END HI[199]
  PIN HI[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 162.930 0.000 163.210 3.000 ;
    END
  END HI[19]
  PIN HI[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 3.000 ;
    END
  END HI[1]
  PIN HI[200]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 3.000 ;
    END
  END HI[200]
  PIN HI[201]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 3.000 ;
    END
  END HI[201]
  PIN HI[202]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 109.110 0.000 109.390 3.000 ;
    END
  END HI[202]
  PIN HI[203]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 236.070 0.000 236.350 3.000 ;
    END
  END HI[203]
  PIN HI[204]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 3.000 ;
    END
  END HI[204]
  PIN HI[205]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 3.000 ;
    END
  END HI[205]
  PIN HI[206]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 3.000 ;
    END
  END HI[206]
  PIN HI[207]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 237.450 0.000 237.730 3.000 ;
    END
  END HI[207]
  PIN HI[208]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 111.870 0.000 112.150 3.000 ;
    END
  END HI[208]
  PIN HI[209]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 4.230 0.000 4.510 3.000 ;
    END
  END HI[209]
  PIN HI[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 3.000 ;
    END
  END HI[20]
  PIN HI[210]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 3.000 ;
    END
  END HI[210]
  PIN HI[211]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 238.830 0.000 239.110 3.000 ;
    END
  END HI[211]
  PIN HI[212]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 169.830 0.000 170.110 3.000 ;
    END
  END HI[212]
  PIN HI[213]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 114.630 0.000 114.910 3.000 ;
    END
  END HI[213]
  PIN HI[214]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 3.000 ;
    END
  END HI[214]
  PIN HI[215]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 171.210 0.000 171.490 3.000 ;
    END
  END HI[215]
  PIN HI[216]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 240.210 0.000 240.490 3.000 ;
    END
  END HI[216]
  PIN HI[217]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 92.550 0.000 92.830 3.000 ;
    END
  END HI[217]
  PIN HI[218]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 172.590 0.000 172.870 3.000 ;
    END
  END HI[218]
  PIN HI[219]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 117.390 0.000 117.670 3.000 ;
    END
  END HI[219]
  PIN HI[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 3.000 ;
    END
  END HI[21]
  PIN HI[220]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 3.000 ;
    END
  END HI[220]
  PIN HI[221]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 3.000 ;
    END
  END HI[221]
  PIN HI[222]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 3.000 ;
    END
  END HI[222]
  PIN HI[223]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 3.000 ;
    END
  END HI[223]
  PIN HI[224]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 120.150 0.000 120.430 3.000 ;
    END
  END HI[224]
  PIN HI[225]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 3.000 ;
    END
  END HI[225]
  PIN HI[226]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 176.730 0.000 177.010 3.000 ;
    END
  END HI[226]
  PIN HI[227]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 3.000 ;
    END
  END HI[227]
  PIN HI[228]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 3.000 ;
    END
  END HI[228]
  PIN HI[229]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 178.110 0.000 178.390 3.000 ;
    END
  END HI[229]
  PIN HI[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 3.000 ;
    END
  END HI[22]
  PIN HI[230]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 3.000 ;
    END
  END HI[230]
  PIN HI[231]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 179.490 0.000 179.770 3.000 ;
    END
  END HI[231]
  PIN HI[232]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 196.050 0.000 196.330 3.000 ;
    END
  END HI[232]
  PIN HI[233]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 3.000 ;
    END
  END HI[233]
  PIN HI[234]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 180.870 0.000 181.150 3.000 ;
    END
  END HI[234]
  PIN HI[235]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 3.000 ;
    END
  END HI[235]
  PIN HI[236]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 100.830 0.000 101.110 3.000 ;
    END
  END HI[236]
  PIN HI[237]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 182.250 0.000 182.530 3.000 ;
    END
  END HI[237]
  PIN HI[238]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 263.670 0.000 263.950 3.000 ;
    END
  END HI[238]
  PIN HI[239]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 274.710 0.000 274.990 3.000 ;
    END
  END HI[239]
  PIN HI[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 3.000 ;
    END
  END HI[23]
  PIN HI[240]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 128.430 0.000 128.710 3.000 ;
    END
  END HI[240]
  PIN HI[241]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 3.000 ;
    END
  END HI[241]
  PIN HI[242]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 3.000 ;
    END
  END HI[242]
  PIN HI[243]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 3.000 ;
    END
  END HI[243]
  PIN HI[244]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 3.000 ;
    END
  END HI[244]
  PIN HI[245]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 186.390 0.000 186.670 3.000 ;
    END
  END HI[245]
  PIN HI[246]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 3.000 ;
    END
  END HI[246]
  PIN HI[247]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 73.230 0.000 73.510 3.000 ;
    END
  END HI[247]
  PIN HI[248]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 3.000 ;
    END
  END HI[248]
  PIN HI[249]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 265.050 0.000 265.330 3.000 ;
    END
  END HI[249]
  PIN HI[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 167.070 0.000 167.350 3.000 ;
    END
  END HI[24]
  PIN HI[250]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 189.150 0.000 189.430 3.000 ;
    END
  END HI[250]
  PIN HI[251]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 133.950 0.000 134.230 3.000 ;
    END
  END HI[251]
  PIN HI[252]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 3.000 ;
    END
  END HI[252]
  PIN HI[253]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 3.000 ;
    END
  END HI[253]
  PIN HI[254]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 3.000 ;
    END
  END HI[254]
  PIN HI[255]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 3.000 ;
    END
  END HI[255]
  PIN HI[256]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 191.910 0.000 192.190 3.000 ;
    END
  END HI[256]
  PIN HI[257]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 136.710 0.000 136.990 3.000 ;
    END
  END HI[257]
  PIN HI[258]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 81.510 0.000 81.790 3.000 ;
    END
  END HI[258]
  PIN HI[259]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 3.000 ;
    END
  END HI[259]
  PIN HI[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 3.000 ;
    END
  END HI[25]
  PIN HI[260]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 3.000 ;
    END
  END HI[260]
  PIN HI[261]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 194.670 0.000 194.950 3.000 ;
    END
  END HI[261]
  PIN HI[262]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 3.000 ;
    END
  END HI[262]
  PIN HI[263]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 3.000 ;
    END
  END HI[263]
  PIN HI[264]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 3.000 ;
    END
  END HI[264]
  PIN HI[265]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 244.350 0.000 244.630 3.000 ;
    END
  END HI[265]
  PIN HI[266]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 140.850 0.000 141.130 3.000 ;
    END
  END HI[266]
  PIN HI[267]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 3.000 ;
    END
  END HI[267]
  PIN HI[268]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 3.000 ;
    END
  END HI[268]
  PIN HI[269]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 197.430 0.000 197.710 3.000 ;
    END
  END HI[269]
  PIN HI[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 3.000 ;
    END
  END HI[26]
  PIN HI[270]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 3.000 ;
    END
  END HI[270]
  PIN HI[271]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 3.000 ;
    END
  END HI[271]
  PIN HI[272]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 198.810 0.000 199.090 3.000 ;
    END
  END HI[272]
  PIN HI[273]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 3.000 ;
    END
  END HI[273]
  PIN HI[274]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 3.000 ;
    END
  END HI[274]
  PIN HI[275]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 245.730 0.000 246.010 3.000 ;
    END
  END HI[275]
  PIN HI[276]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 200.190 0.000 200.470 3.000 ;
    END
  END HI[276]
  PIN HI[277]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 3.000 ;
    END
  END HI[277]
  PIN HI[278]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 3.000 ;
    END
  END HI[278]
  PIN HI[279]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 146.370 0.000 146.650 3.000 ;
    END
  END HI[279]
  PIN HI[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 201.570 0.000 201.850 3.000 ;
    END
  END HI[27]
  PIN HI[280]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 3.000 ;
    END
  END HI[280]
  PIN HI[281]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 247.110 0.000 247.390 3.000 ;
    END
  END HI[281]
  PIN HI[282]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 3.000 ;
    END
  END HI[282]
  PIN HI[283]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 3.000 ;
    END
  END HI[283]
  PIN HI[284]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 3.000 ;
    END
  END HI[284]
  PIN HI[285]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 3.000 ;
    END
  END HI[285]
  PIN HI[286]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 3.000 ;
    END
  END HI[286]
  PIN HI[287]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 204.330 0.000 204.610 3.000 ;
    END
  END HI[287]
  PIN HI[288]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 3.000 ;
    END
  END HI[288]
  PIN HI[289]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 150.510 0.000 150.790 3.000 ;
    END
  END HI[289]
  PIN HI[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 3.000 ;
    END
  END HI[28]
  PIN HI[290]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 3.000 ;
    END
  END HI[290]
  PIN HI[291]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 23.550 0.000 23.830 3.000 ;
    END
  END HI[291]
  PIN HI[292]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 107.730 0.000 108.010 3.000 ;
    END
  END HI[292]
  PIN HI[293]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 3.000 ;
    END
  END HI[293]
  PIN HI[294]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 207.090 0.000 207.370 3.000 ;
    END
  END HI[294]
  PIN HI[295]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 248.490 0.000 248.770 3.000 ;
    END
  END HI[295]
  PIN HI[296]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 153.270 0.000 153.550 3.000 ;
    END
  END HI[296]
  PIN HI[297]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 12.510 0.000 12.790 3.000 ;
    END
  END HI[297]
  PIN HI[298]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 208.470 0.000 208.750 3.000 ;
    END
  END HI[298]
  PIN HI[299]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 3.000 ;
    END
  END HI[299]
  PIN HI[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 3.000 ;
    END
  END HI[29]
  PIN HI[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 3.000 ;
    END
  END HI[2]
  PIN HI[300]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 3.000 ;
    END
  END HI[300]
  PIN HI[301]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 249.870 0.000 250.150 3.000 ;
    END
  END HI[301]
  PIN HI[302]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 3.000 ;
    END
  END HI[302]
  PIN HI[303]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 3.000 ;
    END
  END HI[303]
  PIN HI[304]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 211.230 0.000 211.510 3.000 ;
    END
  END HI[304]
  PIN HI[305]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 3.000 ;
    END
  END HI[305]
  PIN HI[306]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 3.000 ;
    END
  END HI[306]
  PIN HI[307]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 266.430 0.000 266.710 3.000 ;
    END
  END HI[307]
  PIN HI[308]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 271.950 0.000 272.230 3.000 ;
    END
  END HI[308]
  PIN HI[309]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 215.370 0.000 215.650 3.000 ;
    END
  END HI[309]
  PIN HI[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 158.790 0.000 159.070 3.000 ;
    END
  END HI[30]
  PIN HI[310]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 3.000 ;
    END
  END HI[310]
  PIN HI[311]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 213.990 0.000 214.270 3.000 ;
    END
  END HI[311]
  PIN HI[312]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 3.000 ;
    END
  END HI[312]
  PIN HI[313]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 218.130 0.000 218.410 3.000 ;
    END
  END HI[313]
  PIN HI[314]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 252.630 0.000 252.910 3.000 ;
    END
  END HI[314]
  PIN HI[315]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 223.650 0.000 223.930 3.000 ;
    END
  END HI[315]
  PIN HI[316]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 3.000 ;
    END
  END HI[316]
  PIN HI[317]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 3.000 ;
    END
  END HI[317]
  PIN HI[318]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 3.000 ;
    END
  END HI[318]
  PIN HI[319]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 216.750 0.000 217.030 3.000 ;
    END
  END HI[319]
  PIN HI[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 3.000 ;
    END
  END HI[31]
  PIN HI[320]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 3.000 ;
    END
  END HI[320]
  PIN HI[321]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 3.000 ;
    END
  END HI[321]
  PIN HI[322]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 229.170 0.000 229.450 3.000 ;
    END
  END HI[322]
  PIN HI[323]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 254.010 0.000 254.290 3.000 ;
    END
  END HI[323]
  PIN HI[324]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 3.000 ;
    END
  END HI[324]
  PIN HI[325]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 3.000 ;
    END
  END HI[325]
  PIN HI[326]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 219.510 0.000 219.790 3.000 ;
    END
  END HI[326]
  PIN HI[327]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 18.030 0.000 18.310 3.000 ;
    END
  END HI[327]
  PIN HI[328]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 3.000 ;
    END
  END HI[328]
  PIN HI[329]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 40.110 0.000 40.390 3.000 ;
    END
  END HI[329]
  PIN HI[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 220.890 0.000 221.170 3.000 ;
    END
  END HI[32]
  PIN HI[330]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 3.000 ;
    END
  END HI[330]
  PIN HI[331]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 267.810 0.000 268.090 3.000 ;
    END
  END HI[331]
  PIN HI[332]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 3.000 ;
    END
  END HI[332]
  PIN HI[333]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 3.000 ;
    END
  END HI[333]
  PIN HI[334]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 139.470 0.000 139.750 3.000 ;
    END
  END HI[334]
  PIN HI[335]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 3.000 ;
    END
  END HI[335]
  PIN HI[336]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 3.000 ;
    END
  END HI[336]
  PIN HI[337]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 255.390 0.000 255.670 3.000 ;
    END
  END HI[337]
  PIN HI[338]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 3.000 ;
    END
  END HI[338]
  PIN HI[339]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 3.000 ;
    END
  END HI[339]
  PIN HI[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 142.230 0.000 142.510 3.000 ;
    END
  END HI[33]
  PIN HI[340]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 3.000 ;
    END
  END HI[340]
  PIN HI[341]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 269.190 0.000 269.470 3.000 ;
    END
  END HI[341]
  PIN HI[342]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 225.030 0.000 225.310 3.000 ;
    END
  END HI[342]
  PIN HI[343]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 339.570 19.000 339.850 22.000 ;
    END
  END HI[343]
  PIN HI[344]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 74.610 19.000 74.890 22.000 ;
    END
  END HI[344]
  PIN HI[345]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 75.990 19.000 76.270 22.000 ;
    END
  END HI[345]
  PIN HI[346]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 77.370 19.000 77.650 22.000 ;
    END
  END HI[346]
  PIN HI[347]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 78.750 19.000 79.030 22.000 ;
    END
  END HI[347]
  PIN HI[348]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 80.130 19.000 80.410 22.000 ;
    END
  END HI[348]
  PIN HI[349]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 81.510 19.000 81.790 22.000 ;
    END
  END HI[349]
  PIN HI[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 82.890 19.000 83.170 22.000 ;
    END
  END HI[34]
  PIN HI[350]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 84.270 19.000 84.550 22.000 ;
    END
  END HI[350]
  PIN HI[351]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 85.650 19.000 85.930 22.000 ;
    END
  END HI[351]
  PIN HI[352]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 87.030 19.000 87.310 22.000 ;
    END
  END HI[352]
  PIN HI[353]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 88.410 19.000 88.690 22.000 ;
    END
  END HI[353]
  PIN HI[354]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 89.790 19.000 90.070 22.000 ;
    END
  END HI[354]
  PIN HI[355]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 91.170 19.000 91.450 22.000 ;
    END
  END HI[355]
  PIN HI[356]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 92.550 19.000 92.830 22.000 ;
    END
  END HI[356]
  PIN HI[357]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 93.930 19.000 94.210 22.000 ;
    END
  END HI[357]
  PIN HI[358]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 95.310 19.000 95.590 22.000 ;
    END
  END HI[358]
  PIN HI[359]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 96.690 19.000 96.970 22.000 ;
    END
  END HI[359]
  PIN HI[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 98.070 19.000 98.350 22.000 ;
    END
  END HI[35]
  PIN HI[360]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 99.450 19.000 99.730 22.000 ;
    END
  END HI[360]
  PIN HI[361]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 100.830 19.000 101.110 22.000 ;
    END
  END HI[361]
  PIN HI[362]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 102.210 19.000 102.490 22.000 ;
    END
  END HI[362]
  PIN HI[363]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 103.590 19.000 103.870 22.000 ;
    END
  END HI[363]
  PIN HI[364]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 104.970 19.000 105.250 22.000 ;
    END
  END HI[364]
  PIN HI[365]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 106.350 19.000 106.630 22.000 ;
    END
  END HI[365]
  PIN HI[366]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 107.730 19.000 108.010 22.000 ;
    END
  END HI[366]
  PIN HI[367]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 109.110 19.000 109.390 22.000 ;
    END
  END HI[367]
  PIN HI[368]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 110.490 19.000 110.770 22.000 ;
    END
  END HI[368]
  PIN HI[369]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 111.870 19.000 112.150 22.000 ;
    END
  END HI[369]
  PIN HI[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 113.250 19.000 113.530 22.000 ;
    END
  END HI[36]
  PIN HI[370]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 114.630 19.000 114.910 22.000 ;
    END
  END HI[370]
  PIN HI[371]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 116.010 19.000 116.290 22.000 ;
    END
  END HI[371]
  PIN HI[372]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 117.390 19.000 117.670 22.000 ;
    END
  END HI[372]
  PIN HI[373]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 118.770 19.000 119.050 22.000 ;
    END
  END HI[373]
  PIN HI[374]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 120.150 19.000 120.430 22.000 ;
    END
  END HI[374]
  PIN HI[375]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 121.530 19.000 121.810 22.000 ;
    END
  END HI[375]
  PIN HI[376]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 122.910 19.000 123.190 22.000 ;
    END
  END HI[376]
  PIN HI[377]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 124.290 19.000 124.570 22.000 ;
    END
  END HI[377]
  PIN HI[378]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 125.670 19.000 125.950 22.000 ;
    END
  END HI[378]
  PIN HI[379]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 127.050 19.000 127.330 22.000 ;
    END
  END HI[379]
  PIN HI[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 128.430 19.000 128.710 22.000 ;
    END
  END HI[37]
  PIN HI[380]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 129.810 19.000 130.090 22.000 ;
    END
  END HI[380]
  PIN HI[381]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 131.190 19.000 131.470 22.000 ;
    END
  END HI[381]
  PIN HI[382]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 132.570 19.000 132.850 22.000 ;
    END
  END HI[382]
  PIN HI[383]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 133.950 19.000 134.230 22.000 ;
    END
  END HI[383]
  PIN HI[384]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 135.330 19.000 135.610 22.000 ;
    END
  END HI[384]
  PIN HI[385]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 136.710 19.000 136.990 22.000 ;
    END
  END HI[385]
  PIN HI[386]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 138.090 19.000 138.370 22.000 ;
    END
  END HI[386]
  PIN HI[387]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 139.470 19.000 139.750 22.000 ;
    END
  END HI[387]
  PIN HI[388]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 140.850 19.000 141.130 22.000 ;
    END
  END HI[388]
  PIN HI[389]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 142.230 19.000 142.510 22.000 ;
    END
  END HI[389]
  PIN HI[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 143.610 19.000 143.890 22.000 ;
    END
  END HI[38]
  PIN HI[390]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 144.990 19.000 145.270 22.000 ;
    END
  END HI[390]
  PIN HI[391]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 146.370 19.000 146.650 22.000 ;
    END
  END HI[391]
  PIN HI[392]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 147.750 19.000 148.030 22.000 ;
    END
  END HI[392]
  PIN HI[393]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 149.130 19.000 149.410 22.000 ;
    END
  END HI[393]
  PIN HI[394]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 150.510 19.000 150.790 22.000 ;
    END
  END HI[394]
  PIN HI[395]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 151.890 19.000 152.170 22.000 ;
    END
  END HI[395]
  PIN HI[396]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 153.270 19.000 153.550 22.000 ;
    END
  END HI[396]
  PIN HI[397]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 154.650 19.000 154.930 22.000 ;
    END
  END HI[397]
  PIN HI[398]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 156.030 19.000 156.310 22.000 ;
    END
  END HI[398]
  PIN HI[399]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 157.410 19.000 157.690 22.000 ;
    END
  END HI[399]
  PIN HI[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 158.790 19.000 159.070 22.000 ;
    END
  END HI[39]
  PIN HI[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 160.170 19.000 160.450 22.000 ;
    END
  END HI[3]
  PIN HI[400]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 161.550 19.000 161.830 22.000 ;
    END
  END HI[400]
  PIN HI[401]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 162.930 19.000 163.210 22.000 ;
    END
  END HI[401]
  PIN HI[402]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 164.310 19.000 164.590 22.000 ;
    END
  END HI[402]
  PIN HI[403]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 165.690 19.000 165.970 22.000 ;
    END
  END HI[403]
  PIN HI[404]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 167.070 19.000 167.350 22.000 ;
    END
  END HI[404]
  PIN HI[405]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 168.450 19.000 168.730 22.000 ;
    END
  END HI[405]
  PIN HI[406]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 169.830 19.000 170.110 22.000 ;
    END
  END HI[406]
  PIN HI[407]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 171.210 19.000 171.490 22.000 ;
    END
  END HI[407]
  PIN HI[408]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 172.590 19.000 172.870 22.000 ;
    END
  END HI[408]
  PIN HI[409]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 173.970 19.000 174.250 22.000 ;
    END
  END HI[409]
  PIN HI[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 175.350 19.000 175.630 22.000 ;
    END
  END HI[40]
  PIN HI[410]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 176.730 19.000 177.010 22.000 ;
    END
  END HI[410]
  PIN HI[411]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 178.110 19.000 178.390 22.000 ;
    END
  END HI[411]
  PIN HI[412]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 179.490 19.000 179.770 22.000 ;
    END
  END HI[412]
  PIN HI[413]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 180.870 19.000 181.150 22.000 ;
    END
  END HI[413]
  PIN HI[414]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 182.250 19.000 182.530 22.000 ;
    END
  END HI[414]
  PIN HI[415]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 183.630 19.000 183.910 22.000 ;
    END
  END HI[415]
  PIN HI[416]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 185.010 19.000 185.290 22.000 ;
    END
  END HI[416]
  PIN HI[417]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 186.390 19.000 186.670 22.000 ;
    END
  END HI[417]
  PIN HI[418]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 187.770 19.000 188.050 22.000 ;
    END
  END HI[418]
  PIN HI[419]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 189.150 19.000 189.430 22.000 ;
    END
  END HI[419]
  PIN HI[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 190.530 19.000 190.810 22.000 ;
    END
  END HI[41]
  PIN HI[420]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 191.910 19.000 192.190 22.000 ;
    END
  END HI[420]
  PIN HI[421]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 193.290 19.000 193.570 22.000 ;
    END
  END HI[421]
  PIN HI[422]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 194.670 19.000 194.950 22.000 ;
    END
  END HI[422]
  PIN HI[423]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 196.050 19.000 196.330 22.000 ;
    END
  END HI[423]
  PIN HI[424]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 197.430 19.000 197.710 22.000 ;
    END
  END HI[424]
  PIN HI[425]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 198.810 19.000 199.090 22.000 ;
    END
  END HI[425]
  PIN HI[426]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 200.190 19.000 200.470 22.000 ;
    END
  END HI[426]
  PIN HI[427]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 201.570 19.000 201.850 22.000 ;
    END
  END HI[427]
  PIN HI[428]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 202.950 19.000 203.230 22.000 ;
    END
  END HI[428]
  PIN HI[429]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 204.330 19.000 204.610 22.000 ;
    END
  END HI[429]
  PIN HI[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 205.710 19.000 205.990 22.000 ;
    END
  END HI[42]
  PIN HI[430]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 207.090 19.000 207.370 22.000 ;
    END
  END HI[430]
  PIN HI[431]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 208.470 19.000 208.750 22.000 ;
    END
  END HI[431]
  PIN HI[432]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 209.850 19.000 210.130 22.000 ;
    END
  END HI[432]
  PIN HI[433]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 211.230 19.000 211.510 22.000 ;
    END
  END HI[433]
  PIN HI[434]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 212.610 19.000 212.890 22.000 ;
    END
  END HI[434]
  PIN HI[435]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 213.990 19.000 214.270 22.000 ;
    END
  END HI[435]
  PIN HI[436]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 215.370 19.000 215.650 22.000 ;
    END
  END HI[436]
  PIN HI[437]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 216.750 19.000 217.030 22.000 ;
    END
  END HI[437]
  PIN HI[438]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 218.130 19.000 218.410 22.000 ;
    END
  END HI[438]
  PIN HI[439]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 219.510 19.000 219.790 22.000 ;
    END
  END HI[439]
  PIN HI[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 220.890 19.000 221.170 22.000 ;
    END
  END HI[43]
  PIN HI[440]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 222.270 19.000 222.550 22.000 ;
    END
  END HI[440]
  PIN HI[441]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 223.650 19.000 223.930 22.000 ;
    END
  END HI[441]
  PIN HI[442]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 225.030 19.000 225.310 22.000 ;
    END
  END HI[442]
  PIN HI[443]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 226.410 19.000 226.690 22.000 ;
    END
  END HI[443]
  PIN HI[444]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 227.790 19.000 228.070 22.000 ;
    END
  END HI[444]
  PIN HI[445]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 229.170 19.000 229.450 22.000 ;
    END
  END HI[445]
  PIN HI[446]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 230.550 19.000 230.830 22.000 ;
    END
  END HI[446]
  PIN HI[447]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 231.930 19.000 232.210 22.000 ;
    END
  END HI[447]
  PIN HI[448]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 233.310 19.000 233.590 22.000 ;
    END
  END HI[448]
  PIN HI[449]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 234.690 19.000 234.970 22.000 ;
    END
  END HI[449]
  PIN HI[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 236.070 19.000 236.350 22.000 ;
    END
  END HI[44]
  PIN HI[450]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 237.450 19.000 237.730 22.000 ;
    END
  END HI[450]
  PIN HI[451]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 238.830 19.000 239.110 22.000 ;
    END
  END HI[451]
  PIN HI[452]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 240.210 19.000 240.490 22.000 ;
    END
  END HI[452]
  PIN HI[453]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 241.590 19.000 241.870 22.000 ;
    END
  END HI[453]
  PIN HI[454]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 242.970 19.000 243.250 22.000 ;
    END
  END HI[454]
  PIN HI[455]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 244.350 19.000 244.630 22.000 ;
    END
  END HI[455]
  PIN HI[456]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 245.730 19.000 246.010 22.000 ;
    END
  END HI[456]
  PIN HI[457]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 247.110 19.000 247.390 22.000 ;
    END
  END HI[457]
  PIN HI[458]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 248.490 19.000 248.770 22.000 ;
    END
  END HI[458]
  PIN HI[459]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 249.870 19.000 250.150 22.000 ;
    END
  END HI[459]
  PIN HI[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 251.250 19.000 251.530 22.000 ;
    END
  END HI[45]
  PIN HI[460]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 252.630 19.000 252.910 22.000 ;
    END
  END HI[460]
  PIN HI[461]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 254.010 19.000 254.290 22.000 ;
    END
  END HI[461]
  PIN HI[462]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 255.390 19.000 255.670 22.000 ;
    END
  END HI[462]
  PIN HI[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 256.770 19.000 257.050 22.000 ;
    END
  END HI[46]
  PIN HI[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 258.150 19.000 258.430 22.000 ;
    END
  END HI[47]
  PIN HI[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 259.530 19.000 259.810 22.000 ;
    END
  END HI[48]
  PIN HI[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 260.910 19.000 261.190 22.000 ;
    END
  END HI[49]
  PIN HI[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 262.290 19.000 262.570 22.000 ;
    END
  END HI[4]
  PIN HI[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 263.670 19.000 263.950 22.000 ;
    END
  END HI[50]
  PIN HI[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 265.050 19.000 265.330 22.000 ;
    END
  END HI[51]
  PIN HI[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 266.430 19.000 266.710 22.000 ;
    END
  END HI[52]
  PIN HI[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 267.810 19.000 268.090 22.000 ;
    END
  END HI[53]
  PIN HI[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 269.190 19.000 269.470 22.000 ;
    END
  END HI[54]
  PIN HI[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 270.570 19.000 270.850 22.000 ;
    END
  END HI[55]
  PIN HI[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 271.950 19.000 272.230 22.000 ;
    END
  END HI[56]
  PIN HI[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 273.330 19.000 273.610 22.000 ;
    END
  END HI[57]
  PIN HI[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 274.710 19.000 274.990 22.000 ;
    END
  END HI[58]
  PIN HI[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 276.090 19.000 276.370 22.000 ;
    END
  END HI[59]
  PIN HI[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 277.470 19.000 277.750 22.000 ;
    END
  END HI[5]
  PIN HI[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 278.850 19.000 279.130 22.000 ;
    END
  END HI[60]
  PIN HI[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 280.230 19.000 280.510 22.000 ;
    END
  END HI[61]
  PIN HI[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 281.610 19.000 281.890 22.000 ;
    END
  END HI[62]
  PIN HI[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 282.990 19.000 283.270 22.000 ;
    END
  END HI[63]
  PIN HI[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 284.370 19.000 284.650 22.000 ;
    END
  END HI[64]
  PIN HI[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 285.750 19.000 286.030 22.000 ;
    END
  END HI[65]
  PIN HI[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 287.130 19.000 287.410 22.000 ;
    END
  END HI[66]
  PIN HI[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 288.510 19.000 288.790 22.000 ;
    END
  END HI[67]
  PIN HI[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 289.890 19.000 290.170 22.000 ;
    END
  END HI[68]
  PIN HI[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 291.270 19.000 291.550 22.000 ;
    END
  END HI[69]
  PIN HI[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 292.650 19.000 292.930 22.000 ;
    END
  END HI[6]
  PIN HI[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 294.030 19.000 294.310 22.000 ;
    END
  END HI[70]
  PIN HI[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 295.410 19.000 295.690 22.000 ;
    END
  END HI[71]
  PIN HI[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 296.790 19.000 297.070 22.000 ;
    END
  END HI[72]
  PIN HI[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 298.170 19.000 298.450 22.000 ;
    END
  END HI[73]
  PIN HI[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 299.550 19.000 299.830 22.000 ;
    END
  END HI[74]
  PIN HI[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 300.930 19.000 301.210 22.000 ;
    END
  END HI[75]
  PIN HI[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 302.310 19.000 302.590 22.000 ;
    END
  END HI[76]
  PIN HI[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 303.690 19.000 303.970 22.000 ;
    END
  END HI[77]
  PIN HI[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 305.070 19.000 305.350 22.000 ;
    END
  END HI[78]
  PIN HI[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 306.450 19.000 306.730 22.000 ;
    END
  END HI[79]
  PIN HI[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 307.830 19.000 308.110 22.000 ;
    END
  END HI[7]
  PIN HI[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 309.210 19.000 309.490 22.000 ;
    END
  END HI[80]
  PIN HI[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 310.590 19.000 310.870 22.000 ;
    END
  END HI[81]
  PIN HI[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 311.970 19.000 312.250 22.000 ;
    END
  END HI[82]
  PIN HI[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 313.350 19.000 313.630 22.000 ;
    END
  END HI[83]
  PIN HI[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 314.730 19.000 315.010 22.000 ;
    END
  END HI[84]
  PIN HI[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 316.110 19.000 316.390 22.000 ;
    END
  END HI[85]
  PIN HI[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 317.490 19.000 317.770 22.000 ;
    END
  END HI[86]
  PIN HI[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 318.870 19.000 319.150 22.000 ;
    END
  END HI[87]
  PIN HI[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 320.250 19.000 320.530 22.000 ;
    END
  END HI[88]
  PIN HI[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 321.630 19.000 321.910 22.000 ;
    END
  END HI[89]
  PIN HI[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 323.010 19.000 323.290 22.000 ;
    END
  END HI[8]
  PIN HI[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 324.390 19.000 324.670 22.000 ;
    END
  END HI[90]
  PIN HI[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 325.770 19.000 326.050 22.000 ;
    END
  END HI[91]
  PIN HI[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 327.150 19.000 327.430 22.000 ;
    END
  END HI[92]
  PIN HI[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 328.530 19.000 328.810 22.000 ;
    END
  END HI[93]
  PIN HI[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 329.910 19.000 330.190 22.000 ;
    END
  END HI[94]
  PIN HI[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 331.290 19.000 331.570 22.000 ;
    END
  END HI[95]
  PIN HI[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 332.670 19.000 332.950 22.000 ;
    END
  END HI[96]
  PIN HI[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 334.050 19.000 334.330 22.000 ;
    END
  END HI[97]
  PIN HI[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 335.430 19.000 335.710 22.000 ;
    END
  END HI[98]
  PIN HI[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 336.810 19.000 337.090 22.000 ;
    END
  END HI[99]
  PIN HI[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 338.190 19.000 338.470 22.000 ;
    END
  END HI[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 6.440 5.950 344.080 6.450 ;
    END
    PORT
      LAYER met2 ;
        RECT 36.190 5.200 36.690 16.560 ;
    END
    PORT
      LAYER met2 ;
        RECT 96.190 5.200 96.690 16.560 ;
    END
    PORT
      LAYER met2 ;
        RECT 156.190 5.200 156.690 16.560 ;
    END
    PORT
      LAYER met2 ;
        RECT 216.190 5.200 216.690 16.560 ;
    END
    PORT
      LAYER met2 ;
        RECT 276.190 5.200 276.690 16.560 ;
    END
    PORT
      LAYER met2 ;
        RECT 336.190 5.200 336.690 16.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 6.440 11.350 344.080 11.850 ;
    END
    PORT
      LAYER met2 ;
        RECT 66.190 5.200 66.690 16.560 ;
    END
    PORT
      LAYER met2 ;
        RECT 126.190 5.200 126.690 16.560 ;
    END
    PORT
      LAYER met2 ;
        RECT 186.190 5.200 186.690 16.560 ;
    END
    PORT
      LAYER met2 ;
        RECT 246.190 5.200 246.690 16.560 ;
    END
    PORT
      LAYER met2 ;
        RECT 306.190 5.200 306.690 16.560 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 6.440 5.355 344.080 16.405 ;
      LAYER met1 ;
        RECT 0.070 2.760 344.080 17.300 ;
      LAYER met2 ;
        RECT 0.650 18.720 1.190 19.000 ;
        RECT 2.030 18.720 2.570 19.000 ;
        RECT 3.410 18.720 3.950 19.000 ;
        RECT 4.790 18.720 5.330 19.000 ;
        RECT 6.170 18.720 6.710 19.000 ;
        RECT 7.550 18.720 8.090 19.000 ;
        RECT 8.930 18.720 9.470 19.000 ;
        RECT 10.310 18.720 10.850 19.000 ;
        RECT 11.690 18.720 12.230 19.000 ;
        RECT 13.070 18.720 13.610 19.000 ;
        RECT 14.450 18.720 14.990 19.000 ;
        RECT 15.830 18.720 16.370 19.000 ;
        RECT 17.210 18.720 17.750 19.000 ;
        RECT 18.590 18.720 19.130 19.000 ;
        RECT 19.970 18.720 20.510 19.000 ;
        RECT 21.350 18.720 21.890 19.000 ;
        RECT 22.730 18.720 23.270 19.000 ;
        RECT 24.110 18.720 24.650 19.000 ;
        RECT 25.490 18.720 26.030 19.000 ;
        RECT 26.870 18.720 27.410 19.000 ;
        RECT 28.250 18.720 28.790 19.000 ;
        RECT 29.630 18.720 30.170 19.000 ;
        RECT 31.010 18.720 31.550 19.000 ;
        RECT 32.390 18.720 32.930 19.000 ;
        RECT 33.770 18.720 34.310 19.000 ;
        RECT 35.150 18.720 35.690 19.000 ;
        RECT 36.530 18.720 37.070 19.000 ;
        RECT 37.910 18.720 38.450 19.000 ;
        RECT 39.290 18.720 39.830 19.000 ;
        RECT 40.670 18.720 41.210 19.000 ;
        RECT 42.050 18.720 42.590 19.000 ;
        RECT 43.430 18.720 43.970 19.000 ;
        RECT 44.810 18.720 45.350 19.000 ;
        RECT 46.190 18.720 46.730 19.000 ;
        RECT 47.570 18.720 48.110 19.000 ;
        RECT 48.950 18.720 49.490 19.000 ;
        RECT 50.330 18.720 50.870 19.000 ;
        RECT 51.710 18.720 52.250 19.000 ;
        RECT 53.090 18.720 53.630 19.000 ;
        RECT 54.470 18.720 55.010 19.000 ;
        RECT 55.850 18.720 56.390 19.000 ;
        RECT 57.230 18.720 57.770 19.000 ;
        RECT 58.610 18.720 59.150 19.000 ;
        RECT 59.990 18.720 60.530 19.000 ;
        RECT 61.370 18.720 61.910 19.000 ;
        RECT 62.750 18.720 63.290 19.000 ;
        RECT 64.130 18.720 64.670 19.000 ;
        RECT 65.510 18.720 66.050 19.000 ;
        RECT 66.890 18.720 67.430 19.000 ;
        RECT 68.270 18.720 68.810 19.000 ;
        RECT 69.650 18.720 70.190 19.000 ;
        RECT 71.030 18.720 71.570 19.000 ;
        RECT 72.410 18.720 72.950 19.000 ;
        RECT 73.790 18.720 74.330 19.000 ;
        RECT 75.170 18.720 75.710 19.000 ;
        RECT 76.550 18.720 77.090 19.000 ;
        RECT 77.930 18.720 78.470 19.000 ;
        RECT 79.310 18.720 79.850 19.000 ;
        RECT 80.690 18.720 81.230 19.000 ;
        RECT 82.070 18.720 82.610 19.000 ;
        RECT 83.450 18.720 83.990 19.000 ;
        RECT 84.830 18.720 85.370 19.000 ;
        RECT 86.210 18.720 86.750 19.000 ;
        RECT 87.590 18.720 88.130 19.000 ;
        RECT 88.970 18.720 89.510 19.000 ;
        RECT 90.350 18.720 90.890 19.000 ;
        RECT 91.730 18.720 92.270 19.000 ;
        RECT 93.110 18.720 93.650 19.000 ;
        RECT 94.490 18.720 95.030 19.000 ;
        RECT 95.870 18.720 96.410 19.000 ;
        RECT 97.250 18.720 97.790 19.000 ;
        RECT 98.630 18.720 99.170 19.000 ;
        RECT 100.010 18.720 100.550 19.000 ;
        RECT 101.390 18.720 101.930 19.000 ;
        RECT 102.770 18.720 103.310 19.000 ;
        RECT 104.150 18.720 104.690 19.000 ;
        RECT 105.530 18.720 106.070 19.000 ;
        RECT 106.910 18.720 107.450 19.000 ;
        RECT 108.290 18.720 108.830 19.000 ;
        RECT 109.670 18.720 110.210 19.000 ;
        RECT 111.050 18.720 111.590 19.000 ;
        RECT 112.430 18.720 112.970 19.000 ;
        RECT 113.810 18.720 114.350 19.000 ;
        RECT 115.190 18.720 115.730 19.000 ;
        RECT 116.570 18.720 117.110 19.000 ;
        RECT 117.950 18.720 118.490 19.000 ;
        RECT 119.330 18.720 119.870 19.000 ;
        RECT 120.710 18.720 121.250 19.000 ;
        RECT 122.090 18.720 122.630 19.000 ;
        RECT 123.470 18.720 124.010 19.000 ;
        RECT 124.850 18.720 125.390 19.000 ;
        RECT 126.230 18.720 126.770 19.000 ;
        RECT 127.610 18.720 128.150 19.000 ;
        RECT 128.990 18.720 129.530 19.000 ;
        RECT 130.370 18.720 130.910 19.000 ;
        RECT 131.750 18.720 132.290 19.000 ;
        RECT 133.130 18.720 133.670 19.000 ;
        RECT 134.510 18.720 135.050 19.000 ;
        RECT 135.890 18.720 136.430 19.000 ;
        RECT 137.270 18.720 137.810 19.000 ;
        RECT 138.650 18.720 139.190 19.000 ;
        RECT 140.030 18.720 140.570 19.000 ;
        RECT 141.410 18.720 141.950 19.000 ;
        RECT 142.790 18.720 143.330 19.000 ;
        RECT 144.170 18.720 144.710 19.000 ;
        RECT 145.550 18.720 146.090 19.000 ;
        RECT 146.930 18.720 147.470 19.000 ;
        RECT 148.310 18.720 148.850 19.000 ;
        RECT 149.690 18.720 150.230 19.000 ;
        RECT 151.070 18.720 151.610 19.000 ;
        RECT 152.450 18.720 152.990 19.000 ;
        RECT 153.830 18.720 154.370 19.000 ;
        RECT 155.210 18.720 155.750 19.000 ;
        RECT 156.590 18.720 157.130 19.000 ;
        RECT 157.970 18.720 158.510 19.000 ;
        RECT 159.350 18.720 159.890 19.000 ;
        RECT 160.730 18.720 161.270 19.000 ;
        RECT 162.110 18.720 162.650 19.000 ;
        RECT 163.490 18.720 164.030 19.000 ;
        RECT 164.870 18.720 165.410 19.000 ;
        RECT 166.250 18.720 166.790 19.000 ;
        RECT 167.630 18.720 168.170 19.000 ;
        RECT 169.010 18.720 169.550 19.000 ;
        RECT 170.390 18.720 170.930 19.000 ;
        RECT 171.770 18.720 172.310 19.000 ;
        RECT 173.150 18.720 173.690 19.000 ;
        RECT 174.530 18.720 175.070 19.000 ;
        RECT 175.910 18.720 176.450 19.000 ;
        RECT 177.290 18.720 177.830 19.000 ;
        RECT 178.670 18.720 179.210 19.000 ;
        RECT 180.050 18.720 180.590 19.000 ;
        RECT 181.430 18.720 181.970 19.000 ;
        RECT 182.810 18.720 183.350 19.000 ;
        RECT 184.190 18.720 184.730 19.000 ;
        RECT 185.570 18.720 186.110 19.000 ;
        RECT 186.950 18.720 187.490 19.000 ;
        RECT 188.330 18.720 188.870 19.000 ;
        RECT 189.710 18.720 190.250 19.000 ;
        RECT 191.090 18.720 191.630 19.000 ;
        RECT 192.470 18.720 193.010 19.000 ;
        RECT 193.850 18.720 194.390 19.000 ;
        RECT 195.230 18.720 195.770 19.000 ;
        RECT 196.610 18.720 197.150 19.000 ;
        RECT 197.990 18.720 198.530 19.000 ;
        RECT 199.370 18.720 199.910 19.000 ;
        RECT 200.750 18.720 201.290 19.000 ;
        RECT 202.130 18.720 202.670 19.000 ;
        RECT 203.510 18.720 204.050 19.000 ;
        RECT 204.890 18.720 205.430 19.000 ;
        RECT 206.270 18.720 206.810 19.000 ;
        RECT 207.650 18.720 208.190 19.000 ;
        RECT 209.030 18.720 209.570 19.000 ;
        RECT 210.410 18.720 210.950 19.000 ;
        RECT 211.790 18.720 212.330 19.000 ;
        RECT 213.170 18.720 213.710 19.000 ;
        RECT 214.550 18.720 215.090 19.000 ;
        RECT 215.930 18.720 216.470 19.000 ;
        RECT 217.310 18.720 217.850 19.000 ;
        RECT 218.690 18.720 219.230 19.000 ;
        RECT 220.070 18.720 220.610 19.000 ;
        RECT 221.450 18.720 221.990 19.000 ;
        RECT 222.830 18.720 223.370 19.000 ;
        RECT 224.210 18.720 224.750 19.000 ;
        RECT 225.590 18.720 226.130 19.000 ;
        RECT 226.970 18.720 227.510 19.000 ;
        RECT 228.350 18.720 228.890 19.000 ;
        RECT 229.730 18.720 230.270 19.000 ;
        RECT 231.110 18.720 231.650 19.000 ;
        RECT 232.490 18.720 233.030 19.000 ;
        RECT 233.870 18.720 234.410 19.000 ;
        RECT 235.250 18.720 235.790 19.000 ;
        RECT 236.630 18.720 237.170 19.000 ;
        RECT 238.010 18.720 238.550 19.000 ;
        RECT 239.390 18.720 239.930 19.000 ;
        RECT 240.770 18.720 241.310 19.000 ;
        RECT 242.150 18.720 242.690 19.000 ;
        RECT 243.530 18.720 244.070 19.000 ;
        RECT 244.910 18.720 245.450 19.000 ;
        RECT 246.290 18.720 246.830 19.000 ;
        RECT 247.670 18.720 248.210 19.000 ;
        RECT 249.050 18.720 249.590 19.000 ;
        RECT 250.430 18.720 250.970 19.000 ;
        RECT 251.810 18.720 252.350 19.000 ;
        RECT 253.190 18.720 253.730 19.000 ;
        RECT 254.570 18.720 255.110 19.000 ;
        RECT 255.950 18.720 256.490 19.000 ;
        RECT 257.330 18.720 257.870 19.000 ;
        RECT 258.710 18.720 259.250 19.000 ;
        RECT 260.090 18.720 260.630 19.000 ;
        RECT 261.470 18.720 262.010 19.000 ;
        RECT 262.850 18.720 263.390 19.000 ;
        RECT 264.230 18.720 264.770 19.000 ;
        RECT 265.610 18.720 266.150 19.000 ;
        RECT 266.990 18.720 267.530 19.000 ;
        RECT 268.370 18.720 268.910 19.000 ;
        RECT 269.750 18.720 270.290 19.000 ;
        RECT 271.130 18.720 271.670 19.000 ;
        RECT 272.510 18.720 273.050 19.000 ;
        RECT 273.890 18.720 274.430 19.000 ;
        RECT 275.270 18.720 275.810 19.000 ;
        RECT 276.650 18.720 277.190 19.000 ;
        RECT 278.030 18.720 278.570 19.000 ;
        RECT 279.410 18.720 279.950 19.000 ;
        RECT 280.790 18.720 281.330 19.000 ;
        RECT 282.170 18.720 282.710 19.000 ;
        RECT 283.550 18.720 284.090 19.000 ;
        RECT 284.930 18.720 285.470 19.000 ;
        RECT 286.310 18.720 286.850 19.000 ;
        RECT 287.690 18.720 288.230 19.000 ;
        RECT 289.070 18.720 289.610 19.000 ;
        RECT 290.450 18.720 290.990 19.000 ;
        RECT 291.830 18.720 292.370 19.000 ;
        RECT 293.210 18.720 293.750 19.000 ;
        RECT 294.590 18.720 295.130 19.000 ;
        RECT 295.970 18.720 296.510 19.000 ;
        RECT 297.350 18.720 297.890 19.000 ;
        RECT 298.730 18.720 299.270 19.000 ;
        RECT 300.110 18.720 300.650 19.000 ;
        RECT 301.490 18.720 302.030 19.000 ;
        RECT 302.870 18.720 303.410 19.000 ;
        RECT 304.250 18.720 304.790 19.000 ;
        RECT 305.630 18.720 306.170 19.000 ;
        RECT 307.010 18.720 307.550 19.000 ;
        RECT 308.390 18.720 308.930 19.000 ;
        RECT 309.770 18.720 310.310 19.000 ;
        RECT 311.150 18.720 311.690 19.000 ;
        RECT 312.530 18.720 313.070 19.000 ;
        RECT 313.910 18.720 314.450 19.000 ;
        RECT 315.290 18.720 315.830 19.000 ;
        RECT 316.670 18.720 317.210 19.000 ;
        RECT 318.050 18.720 318.590 19.000 ;
        RECT 319.430 18.720 319.970 19.000 ;
        RECT 320.810 18.720 321.350 19.000 ;
        RECT 322.190 18.720 322.730 19.000 ;
        RECT 323.570 18.720 324.110 19.000 ;
        RECT 324.950 18.720 325.490 19.000 ;
        RECT 326.330 18.720 326.870 19.000 ;
        RECT 327.710 18.720 328.250 19.000 ;
        RECT 329.090 18.720 329.630 19.000 ;
        RECT 330.470 18.720 331.010 19.000 ;
        RECT 331.850 18.720 332.390 19.000 ;
        RECT 333.230 18.720 333.770 19.000 ;
        RECT 334.610 18.720 335.150 19.000 ;
        RECT 335.990 18.720 336.530 19.000 ;
        RECT 337.370 18.720 337.910 19.000 ;
        RECT 338.750 18.720 339.290 19.000 ;
        RECT 0.100 16.840 339.840 18.720 ;
        RECT 0.100 4.920 35.910 16.840 ;
        RECT 36.970 4.920 65.910 16.840 ;
        RECT 66.970 4.920 95.910 16.840 ;
        RECT 96.970 4.920 125.910 16.840 ;
        RECT 126.970 4.920 155.910 16.840 ;
        RECT 156.970 4.920 185.910 16.840 ;
        RECT 186.970 4.920 215.910 16.840 ;
        RECT 216.970 4.920 245.910 16.840 ;
        RECT 246.970 4.920 275.910 16.840 ;
        RECT 276.970 4.920 305.910 16.840 ;
        RECT 306.970 4.920 335.910 16.840 ;
        RECT 336.970 4.920 339.840 16.840 ;
        RECT 0.100 3.280 339.840 4.920 ;
        RECT 0.650 2.730 1.190 3.280 ;
        RECT 2.030 2.730 2.570 3.280 ;
        RECT 3.410 2.730 3.950 3.280 ;
        RECT 4.790 2.730 5.330 3.280 ;
        RECT 6.170 2.730 6.710 3.280 ;
        RECT 7.550 2.730 8.090 3.280 ;
        RECT 8.930 2.730 9.470 3.280 ;
        RECT 10.310 2.730 10.850 3.280 ;
        RECT 11.690 2.730 12.230 3.280 ;
        RECT 13.070 2.730 13.610 3.280 ;
        RECT 14.450 2.730 14.990 3.280 ;
        RECT 15.830 2.730 16.370 3.280 ;
        RECT 17.210 2.730 17.750 3.280 ;
        RECT 18.590 2.730 19.130 3.280 ;
        RECT 19.970 2.730 20.510 3.280 ;
        RECT 21.350 2.730 21.890 3.280 ;
        RECT 22.730 2.730 23.270 3.280 ;
        RECT 24.110 2.730 24.650 3.280 ;
        RECT 25.490 2.730 26.030 3.280 ;
        RECT 26.870 2.730 27.410 3.280 ;
        RECT 28.250 2.730 28.790 3.280 ;
        RECT 29.630 2.730 30.170 3.280 ;
        RECT 31.010 2.730 31.550 3.280 ;
        RECT 32.390 2.730 32.930 3.280 ;
        RECT 33.770 2.730 34.310 3.280 ;
        RECT 35.150 2.730 35.690 3.280 ;
        RECT 36.530 2.730 37.070 3.280 ;
        RECT 37.910 2.730 38.450 3.280 ;
        RECT 39.290 2.730 39.830 3.280 ;
        RECT 40.670 2.730 41.210 3.280 ;
        RECT 42.050 2.730 42.590 3.280 ;
        RECT 43.430 2.730 43.970 3.280 ;
        RECT 44.810 2.730 45.350 3.280 ;
        RECT 46.190 2.730 46.730 3.280 ;
        RECT 47.570 2.730 48.110 3.280 ;
        RECT 48.950 2.730 49.490 3.280 ;
        RECT 50.330 2.730 50.870 3.280 ;
        RECT 51.710 2.730 52.250 3.280 ;
        RECT 53.090 2.730 53.630 3.280 ;
        RECT 54.470 2.730 55.010 3.280 ;
        RECT 55.850 2.730 56.390 3.280 ;
        RECT 57.230 2.730 57.770 3.280 ;
        RECT 58.610 2.730 59.150 3.280 ;
        RECT 59.990 2.730 60.530 3.280 ;
        RECT 61.370 2.730 61.910 3.280 ;
        RECT 62.750 2.730 63.290 3.280 ;
        RECT 64.130 2.730 64.670 3.280 ;
        RECT 65.510 2.730 66.050 3.280 ;
        RECT 66.890 2.730 67.430 3.280 ;
        RECT 68.270 2.730 68.810 3.280 ;
        RECT 69.650 2.730 70.190 3.280 ;
        RECT 71.030 2.730 71.570 3.280 ;
        RECT 72.410 2.730 72.950 3.280 ;
        RECT 73.790 2.730 74.330 3.280 ;
        RECT 75.170 2.730 75.710 3.280 ;
        RECT 76.550 2.730 77.090 3.280 ;
        RECT 77.930 2.730 78.470 3.280 ;
        RECT 79.310 2.730 79.850 3.280 ;
        RECT 80.690 2.730 81.230 3.280 ;
        RECT 82.070 2.730 82.610 3.280 ;
        RECT 83.450 2.730 83.990 3.280 ;
        RECT 84.830 2.730 85.370 3.280 ;
        RECT 86.210 2.730 86.750 3.280 ;
        RECT 87.590 2.730 88.130 3.280 ;
        RECT 88.970 2.730 89.510 3.280 ;
        RECT 90.350 2.730 90.890 3.280 ;
        RECT 91.730 2.730 92.270 3.280 ;
        RECT 93.110 2.730 93.650 3.280 ;
        RECT 94.490 2.730 95.030 3.280 ;
        RECT 95.870 2.730 96.410 3.280 ;
        RECT 97.250 2.730 97.790 3.280 ;
        RECT 98.630 2.730 99.170 3.280 ;
        RECT 100.010 2.730 100.550 3.280 ;
        RECT 101.390 2.730 101.930 3.280 ;
        RECT 102.770 2.730 103.310 3.280 ;
        RECT 104.150 2.730 104.690 3.280 ;
        RECT 105.530 2.730 106.070 3.280 ;
        RECT 106.910 2.730 107.450 3.280 ;
        RECT 108.290 2.730 108.830 3.280 ;
        RECT 109.670 2.730 110.210 3.280 ;
        RECT 111.050 2.730 111.590 3.280 ;
        RECT 112.430 2.730 112.970 3.280 ;
        RECT 113.810 2.730 114.350 3.280 ;
        RECT 115.190 2.730 115.730 3.280 ;
        RECT 116.570 2.730 117.110 3.280 ;
        RECT 117.950 2.730 118.490 3.280 ;
        RECT 119.330 2.730 119.870 3.280 ;
        RECT 120.710 2.730 121.250 3.280 ;
        RECT 122.090 2.730 122.630 3.280 ;
        RECT 123.470 2.730 124.010 3.280 ;
        RECT 124.850 2.730 125.390 3.280 ;
        RECT 126.230 2.730 126.770 3.280 ;
        RECT 127.610 2.730 128.150 3.280 ;
        RECT 128.990 2.730 129.530 3.280 ;
        RECT 130.370 2.730 130.910 3.280 ;
        RECT 131.750 2.730 132.290 3.280 ;
        RECT 133.130 2.730 133.670 3.280 ;
        RECT 134.510 2.730 135.050 3.280 ;
        RECT 135.890 2.730 136.430 3.280 ;
        RECT 137.270 2.730 137.810 3.280 ;
        RECT 138.650 2.730 139.190 3.280 ;
        RECT 140.030 2.730 140.570 3.280 ;
        RECT 141.410 2.730 141.950 3.280 ;
        RECT 142.790 2.730 143.330 3.280 ;
        RECT 144.170 2.730 144.710 3.280 ;
        RECT 145.550 2.730 146.090 3.280 ;
        RECT 146.930 2.730 147.470 3.280 ;
        RECT 148.310 2.730 148.850 3.280 ;
        RECT 149.690 2.730 150.230 3.280 ;
        RECT 151.070 2.730 151.610 3.280 ;
        RECT 152.450 2.730 152.990 3.280 ;
        RECT 153.830 2.730 154.370 3.280 ;
        RECT 155.210 2.730 155.750 3.280 ;
        RECT 156.590 2.730 157.130 3.280 ;
        RECT 157.970 2.730 158.510 3.280 ;
        RECT 159.350 2.730 159.890 3.280 ;
        RECT 160.730 2.730 161.270 3.280 ;
        RECT 162.110 2.730 162.650 3.280 ;
        RECT 163.490 2.730 164.030 3.280 ;
        RECT 164.870 2.730 165.410 3.280 ;
        RECT 166.250 2.730 166.790 3.280 ;
        RECT 167.630 2.730 168.170 3.280 ;
        RECT 169.010 2.730 169.550 3.280 ;
        RECT 170.390 2.730 170.930 3.280 ;
        RECT 171.770 2.730 172.310 3.280 ;
        RECT 173.150 2.730 173.690 3.280 ;
        RECT 174.530 2.730 175.070 3.280 ;
        RECT 175.910 2.730 176.450 3.280 ;
        RECT 177.290 2.730 177.830 3.280 ;
        RECT 178.670 2.730 179.210 3.280 ;
        RECT 180.050 2.730 180.590 3.280 ;
        RECT 181.430 2.730 181.970 3.280 ;
        RECT 182.810 2.730 183.350 3.280 ;
        RECT 184.190 2.730 184.730 3.280 ;
        RECT 185.570 2.730 186.110 3.280 ;
        RECT 186.950 2.730 187.490 3.280 ;
        RECT 188.330 2.730 188.870 3.280 ;
        RECT 189.710 2.730 190.250 3.280 ;
        RECT 191.090 2.730 191.630 3.280 ;
        RECT 192.470 2.730 193.010 3.280 ;
        RECT 193.850 2.730 194.390 3.280 ;
        RECT 195.230 2.730 195.770 3.280 ;
        RECT 196.610 2.730 197.150 3.280 ;
        RECT 197.990 2.730 198.530 3.280 ;
        RECT 199.370 2.730 199.910 3.280 ;
        RECT 200.750 2.730 201.290 3.280 ;
        RECT 202.130 2.730 202.670 3.280 ;
        RECT 203.510 2.730 204.050 3.280 ;
        RECT 204.890 2.730 205.430 3.280 ;
        RECT 206.270 2.730 206.810 3.280 ;
        RECT 207.650 2.730 208.190 3.280 ;
        RECT 209.030 2.730 209.570 3.280 ;
        RECT 210.410 2.730 210.950 3.280 ;
        RECT 211.790 2.730 212.330 3.280 ;
        RECT 213.170 2.730 213.710 3.280 ;
        RECT 214.550 2.730 215.090 3.280 ;
        RECT 215.930 2.730 216.470 3.280 ;
        RECT 217.310 2.730 217.850 3.280 ;
        RECT 218.690 2.730 219.230 3.280 ;
        RECT 220.070 2.730 220.610 3.280 ;
        RECT 221.450 2.730 221.990 3.280 ;
        RECT 222.830 2.730 223.370 3.280 ;
        RECT 224.210 2.730 224.750 3.280 ;
        RECT 225.590 2.730 226.130 3.280 ;
        RECT 226.970 2.730 227.510 3.280 ;
        RECT 228.350 2.730 228.890 3.280 ;
        RECT 229.730 2.730 230.270 3.280 ;
        RECT 231.110 2.730 231.650 3.280 ;
        RECT 232.490 2.730 233.030 3.280 ;
        RECT 233.870 2.730 234.410 3.280 ;
        RECT 235.250 2.730 235.790 3.280 ;
        RECT 236.630 2.730 237.170 3.280 ;
        RECT 238.010 2.730 238.550 3.280 ;
        RECT 239.390 2.730 239.930 3.280 ;
        RECT 240.770 2.730 241.310 3.280 ;
        RECT 242.150 2.730 242.690 3.280 ;
        RECT 243.530 2.730 244.070 3.280 ;
        RECT 244.910 2.730 245.450 3.280 ;
        RECT 246.290 2.730 246.830 3.280 ;
        RECT 247.670 2.730 248.210 3.280 ;
        RECT 249.050 2.730 249.590 3.280 ;
        RECT 250.430 2.730 250.970 3.280 ;
        RECT 251.810 2.730 252.350 3.280 ;
        RECT 253.190 2.730 253.730 3.280 ;
        RECT 254.570 2.730 255.110 3.280 ;
        RECT 255.950 2.730 256.490 3.280 ;
        RECT 257.330 2.730 257.870 3.280 ;
        RECT 258.710 2.730 259.250 3.280 ;
        RECT 260.090 2.730 260.630 3.280 ;
        RECT 261.470 2.730 262.010 3.280 ;
        RECT 262.850 2.730 263.390 3.280 ;
        RECT 264.230 2.730 264.770 3.280 ;
        RECT 265.610 2.730 266.150 3.280 ;
        RECT 266.990 2.730 267.530 3.280 ;
        RECT 268.370 2.730 268.910 3.280 ;
        RECT 269.750 2.730 270.290 3.280 ;
        RECT 271.130 2.730 271.670 3.280 ;
        RECT 272.510 2.730 273.050 3.280 ;
        RECT 273.890 2.730 274.430 3.280 ;
        RECT 275.270 2.730 339.840 3.280 ;
      LAYER met3 ;
        RECT 3.400 12.250 21.555 20.890 ;
        RECT 3.400 10.950 6.040 12.250 ;
        RECT 3.400 6.850 21.555 10.950 ;
        RECT 3.400 5.550 6.040 6.850 ;
        RECT 3.400 0.190 21.555 5.550 ;
  END
END mprj_logic_high
END LIBRARY

