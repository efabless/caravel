module chip_io (clock,
    clock_core,
    por,
    flash_clk,
    flash_clk_core,
    flash_clk_oeb_core,
    flash_csb,
    flash_csb_core,
    flash_csb_oeb_core,
    flash_io0,
    flash_io0_di_core,
    flash_io0_do_core,
    flash_io0_ieb_core,
    flash_io0_oeb_core,
    flash_io1,
    flash_io1_di_core,
    flash_io1_do_core,
    flash_io1_oeb_core,
    gpio,
    gpio_in_core,
    gpio_inenb_core,
    gpio_mode0_core,
    gpio_mode1_core,
    gpio_out_core,
    gpio_outenb_core,
    vccd_pad,
    vdda_pad,
    vddio_pad,
    vddio_pad2,
    vssa_pad,
    vssd_pad,
    vssio_pad,
    vssio_pad2,
    resetb,
    vdda,
    vccd1_pad,
    vdda1_pad,
    vdda1_pad2,
    vssa1_pad,
    vssa1_pad2,
    vssd1_pad,
    vccd2_pad,
    vdda2_pad,
    vssa2_pad,
    vdda2,
    vssa2,
    vssd2_pad,
    resetb_core_h,
    vssd2,
    vccd2,
    vssd1,
    vccd1,
    flash_io1_ieb_core,
    porb_h,
    vccd,
    vdda1,
    vddio,
    vssa,
    vssa1,
    vssd,
    vssio,
    mprj_analog_io,
    mprj_io,
    mprj_io_analog_en,
    mprj_io_analog_pol,
    mprj_io_analog_sel,
    mprj_io_dm,
    mprj_io_holdover,
    mprj_io_ib_mode_sel,
    mprj_io_in,
    mprj_io_inp_dis,
    mprj_io_oeb,
    mprj_io_one,
    mprj_io_out,
    mprj_io_slow_sel,
    mprj_io_vtrip_sel);
 input clock;
 inout clock_core;
 input por;
 inout flash_clk;
 input flash_clk_core;
 input flash_clk_oeb_core;
 inout flash_csb;
 input flash_csb_core;
 input flash_csb_oeb_core;
 inout flash_io0;
 inout flash_io0_di_core;
 input flash_io0_do_core;
 input flash_io0_ieb_core;
 input flash_io0_oeb_core;
 inout flash_io1;
 inout flash_io1_di_core;
 input flash_io1_do_core;
 input flash_io1_oeb_core;
 inout gpio;
 inout gpio_in_core;
 input gpio_inenb_core;
 input gpio_mode0_core;
 input gpio_mode1_core;
 input gpio_out_core;
 input gpio_outenb_core;
 inout vccd_pad;
 inout vdda_pad;
 inout vddio_pad;
 inout vddio_pad2;
 inout vssa_pad;
 inout vssd_pad;
 inout vssio_pad;
 inout vssio_pad2;
 input resetb;
 inout vdda;
 inout vccd1_pad;
 inout vdda1_pad;
 inout vdda1_pad2;
 inout vssa1_pad;
 inout vssa1_pad2;
 inout vssd1_pad;
 inout vccd2_pad;
 inout vdda2_pad;
 inout vssa2_pad;
 inout vdda2;
 inout vssa2;
 inout vssd2_pad;
 inout resetb_core_h;
 inout vssd2;
 inout vccd2;
 inout vssd1;
 inout vccd1;
 input flash_io1_ieb_core;
 input porb_h;
 input vccd;
 input vdda1;
 input vddio;
 input vssa;
 input vssa1;
 input vssd;
 input vssio;
 inout [28:0] mprj_analog_io;
 inout [37:0] mprj_io;
 input [37:0] mprj_io_analog_en;
 input [37:0] mprj_io_analog_pol;
 input [37:0] mprj_io_analog_sel;
 input [113:0] mprj_io_dm;
 input [37:0] mprj_io_holdover;
 input [37:0] mprj_io_ib_mode_sel;
 inout [37:0] mprj_io_in;
 input [37:0] mprj_io_inp_dis;
 input [37:0] mprj_io_oeb;
 input [37:0] mprj_io_one;
 input [37:0] mprj_io_out;
 input [37:0] mprj_io_slow_sel;
 input [37:0] mprj_io_vtrip_sel;

 wire clock_pad__OE_N;
 wire \mprj_pads.area1_io_pad[13]__TIE_LO_ESD ;
 wire \mprj_pads.area1_io_pad[13]__HLD_H_N ;
 wire \mprj_pads.area1_io_pad[13]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area1_io_pad[13]__PAD_A_NOESD_H ;
 wire \mprj_pads.area1_io_pad[13]__IN_H ;
 wire flash_clk_pad__TIE_LO_ESD;
 wire flash_clk_pad__IN;
 wire flash_clk_pad__HLD_H_N;
 wire flash_clk_pad__SLOW;
 wire flash_clk_pad__PAD_A_ESD_0_H;
 wire flash_clk_pad__PAD_A_ESD_1_H;
 wire flash_clk_pad__PAD_A_NOESD_H;
 wire flash_clk_pad__IN_H;
 wire constant_block_0__zero;
 wire \mprj_pads.area1_io_pad[9]__TIE_LO_ESD ;
 wire \mprj_pads.area1_io_pad[9]__HLD_H_N ;
 wire \mprj_pads.area1_io_pad[9]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area1_io_pad[9]__PAD_A_NOESD_H ;
 wire \mprj_pads.area1_io_pad[9]__IN_H ;
 wire gpio_pad__VDDIO_Q;
 wire gpio_pad__VSSIO_Q;
 wire gpio_pad__AMUXBUS_A;
 wire gpio_pad__AMUXBUS_B;
 wire flash_io0_pad__TIE_LO_ESD;
 wire flash_io0_pad__HLD_H_N;
 wire flash_io0_pad__SLOW;
 wire flash_io0_pad__PAD_A_ESD_0_H;
 wire flash_io0_pad__PAD_A_ESD_1_H;
 wire flash_io0_pad__PAD_A_NOESD_H;
 wire flash_io0_pad__IN_H;
 wire \mprj_pads.area2_io_pad[9]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area2_io_pad[9]__PAD_A_NOESD_H ;
 wire \mprj_pads.area2_io_pad[9]__HLD_H_N ;
 wire \mprj_pads.area2_io_pad[9]__TIE_LO_ESD ;
 wire \mprj_pads.area2_io_pad[9]__IN_H ;
 wire \mprj_pads.area1_io_pad[15]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area1_io_pad[15]__PAD_A_NOESD_H ;
 wire \mprj_pads.area1_io_pad[15]__HLD_H_N ;
 wire \mprj_pads.area1_io_pad[15]__TIE_LO_ESD ;
 wire \mprj_pads.area1_io_pad[15]__IN_H ;
 wire \mprj_pads.area1_io_pad[0]__TIE_LO_ESD ;
 wire \mprj_pads.area1_io_pad[0]__HLD_H_N ;
 wire \mprj_pads.area1_io_pad[0]__PAD_A_ESD_0_H ;
 wire \mprj_pads.area1_io_pad[0]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area1_io_pad[0]__PAD_A_NOESD_H ;
 wire \mprj_pads.area1_io_pad[0]__IN_H ;
 wire \mprj_pads.area2_io_pad[0]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area2_io_pad[0]__PAD_A_NOESD_H ;
 wire \mprj_pads.area2_io_pad[0]__HLD_H_N ;
 wire \mprj_pads.area2_io_pad[0]__TIE_LO_ESD ;
 wire \mprj_pads.area2_io_pad[0]__IN_H ;
 wire \mprj_pads.area2_io_pad[10]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area2_io_pad[10]__PAD_A_NOESD_H ;
 wire \mprj_pads.area2_io_pad[10]__HLD_H_N ;
 wire \mprj_pads.area2_io_pad[10]__TIE_LO_ESD ;
 wire \mprj_pads.area2_io_pad[10]__IN_H ;
 wire \mprj_pads.area1_io_pad[17]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area1_io_pad[17]__PAD_A_NOESD_H ;
 wire \mprj_pads.area1_io_pad[17]__HLD_H_N ;
 wire \mprj_pads.area1_io_pad[17]__TIE_LO_ESD ;
 wire \mprj_pads.area1_io_pad[17]__IN_H ;
 wire \mprj_pads.area1_io_pad[2]__TIE_LO_ESD ;
 wire \mprj_pads.area1_io_pad[2]__HLD_H_N ;
 wire \mprj_pads.area1_io_pad[2]__PAD_A_ESD_0_H ;
 wire \mprj_pads.area1_io_pad[2]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area1_io_pad[2]__PAD_A_NOESD_H ;
 wire \mprj_pads.area1_io_pad[2]__IN_H ;
 wire \mprj_pads.area2_io_pad[2]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area2_io_pad[2]__PAD_A_NOESD_H ;
 wire \mprj_pads.area2_io_pad[2]__HLD_H_N ;
 wire \mprj_pads.area2_io_pad[2]__TIE_LO_ESD ;
 wire \mprj_pads.area2_io_pad[2]__IN_H ;
 wire \mprj_pads.area2_io_pad[12]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area2_io_pad[12]__PAD_A_NOESD_H ;
 wire \mprj_pads.area2_io_pad[12]__HLD_H_N ;
 wire \mprj_pads.area2_io_pad[12]__TIE_LO_ESD ;
 wire \mprj_pads.area2_io_pad[12]__IN_H ;
 wire \mprj_pads.area1_io_pad[4]__TIE_LO_ESD ;
 wire \mprj_pads.area1_io_pad[4]__HLD_H_N ;
 wire \mprj_pads.area1_io_pad[4]__PAD_A_ESD_0_H ;
 wire \mprj_pads.area1_io_pad[4]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area1_io_pad[4]__PAD_A_NOESD_H ;
 wire \mprj_pads.area1_io_pad[4]__IN_H ;
 wire \mprj_pads.area2_io_pad[4]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area2_io_pad[4]__PAD_A_NOESD_H ;
 wire \mprj_pads.area2_io_pad[4]__HLD_H_N ;
 wire \mprj_pads.area2_io_pad[4]__TIE_LO_ESD ;
 wire \mprj_pads.area2_io_pad[4]__IN_H ;
 wire \mprj_pads.area2_io_pad[14]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area2_io_pad[14]__PAD_A_NOESD_H ;
 wire \mprj_pads.area2_io_pad[14]__HLD_H_N ;
 wire \mprj_pads.area2_io_pad[14]__TIE_LO_ESD ;
 wire \mprj_pads.area2_io_pad[14]__IN_H ;
 wire flash_io1_pad__TIE_LO_ESD;
 wire flash_io1_pad__HLD_H_N;
 wire flash_io1_pad__SLOW;
 wire flash_io1_pad__PAD_A_ESD_0_H;
 wire flash_io1_pad__PAD_A_ESD_1_H;
 wire flash_io1_pad__PAD_A_NOESD_H;
 wire flash_io1_pad__IN_H;
 wire \mprj_pads.area1_io_pad[10]__TIE_LO_ESD ;
 wire \mprj_pads.area1_io_pad[10]__HLD_H_N ;
 wire \mprj_pads.area1_io_pad[10]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area1_io_pad[10]__PAD_A_NOESD_H ;
 wire \mprj_pads.area1_io_pad[10]__IN_H ;
 wire \mprj_pads.area1_io_pad[6]__TIE_LO_ESD ;
 wire \mprj_pads.area1_io_pad[6]__HLD_H_N ;
 wire \mprj_pads.area1_io_pad[6]__PAD_A_ESD_0_H ;
 wire \mprj_pads.area1_io_pad[6]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area1_io_pad[6]__PAD_A_NOESD_H ;
 wire \mprj_pads.area1_io_pad[6]__IN_H ;
 wire flash_csb_pad__TIE_LO_ESD;
 wire flash_csb_pad__IN;
 wire flash_csb_pad__HLD_H_N;
 wire flash_csb_pad__SLOW;
 wire flash_csb_pad__PAD_A_ESD_0_H;
 wire flash_csb_pad__PAD_A_ESD_1_H;
 wire flash_csb_pad__PAD_A_NOESD_H;
 wire flash_csb_pad__IN_H;
 wire \mprj_pads.area2_io_pad[6]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area2_io_pad[6]__PAD_A_NOESD_H ;
 wire \mprj_pads.area2_io_pad[6]__HLD_H_N ;
 wire \mprj_pads.area2_io_pad[6]__TIE_LO_ESD ;
 wire \mprj_pads.area2_io_pad[6]__IN_H ;
 wire \mprj_pads.area2_io_pad[16]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area2_io_pad[16]__PAD_A_NOESD_H ;
 wire \mprj_pads.area2_io_pad[16]__HLD_H_N ;
 wire \mprj_pads.area2_io_pad[16]__TIE_LO_ESD ;
 wire \mprj_pads.area2_io_pad[16]__IN_H ;
 wire \mprj_pads.area1_io_pad[12]__TIE_LO_ESD ;
 wire \mprj_pads.area1_io_pad[12]__HLD_H_N ;
 wire \mprj_pads.area1_io_pad[12]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area1_io_pad[12]__PAD_A_NOESD_H ;
 wire \mprj_pads.area1_io_pad[12]__IN_H ;
 wire xresloop;
 wire constant_block_0__one;
 wire xres_vss_loop;
 wire resetb_pad__TIE_HI_ESD;
 wire \mprj_pads.area1_io_pad[8]__TIE_LO_ESD ;
 wire \mprj_pads.area1_io_pad[8]__HLD_H_N ;
 wire \mprj_pads.area1_io_pad[8]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area1_io_pad[8]__PAD_A_NOESD_H ;
 wire \mprj_pads.area1_io_pad[8]__IN_H ;
 wire \mprj_pads.area2_io_pad[8]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area2_io_pad[8]__PAD_A_NOESD_H ;
 wire \mprj_pads.area2_io_pad[8]__HLD_H_N ;
 wire \mprj_pads.area2_io_pad[8]__TIE_LO_ESD ;
 wire \mprj_pads.area2_io_pad[8]__IN_H ;
 wire \mprj_pads.area2_io_pad[18]__PAD_A_ESD_0_H ;
 wire \mprj_pads.area2_io_pad[18]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area2_io_pad[18]__PAD_A_NOESD_H ;
 wire \mprj_pads.area2_io_pad[18]__HLD_H_N ;
 wire \mprj_pads.area2_io_pad[18]__TIE_LO_ESD ;
 wire \mprj_pads.area2_io_pad[18]__IN_H ;
 wire \mprj_pads.area1_io_pad[14]__TIE_LO_ESD ;
 wire \mprj_pads.area1_io_pad[14]__HLD_H_N ;
 wire \mprj_pads.area1_io_pad[14]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area1_io_pad[14]__PAD_A_NOESD_H ;
 wire \mprj_pads.area1_io_pad[14]__IN_H ;
 wire \mprj_pads.area1_io_pad[16]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area1_io_pad[16]__PAD_A_NOESD_H ;
 wire \mprj_pads.area1_io_pad[16]__HLD_H_N ;
 wire \mprj_pads.area1_io_pad[16]__TIE_LO_ESD ;
 wire \mprj_pads.area1_io_pad[16]__IN_H ;
 wire gpio_pad__TIE_LO_ESD;
 wire gpio_pad__HLD_H_N;
 wire gpio_pad__SLOW;
 wire gpio_pad__PAD_A_ESD_0_H;
 wire gpio_pad__PAD_A_ESD_1_H;
 wire gpio_pad__PAD_A_NOESD_H;
 wire gpio_pad__IN_H;
 wire \mprj_pads.area1_io_pad[1]__TIE_LO_ESD ;
 wire \mprj_pads.area1_io_pad[1]__HLD_H_N ;
 wire \mprj_pads.area1_io_pad[1]__PAD_A_ESD_0_H ;
 wire \mprj_pads.area1_io_pad[1]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area1_io_pad[1]__PAD_A_NOESD_H ;
 wire \mprj_pads.area1_io_pad[1]__IN_H ;
 wire \mprj_pads.area2_io_pad[1]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area2_io_pad[1]__PAD_A_NOESD_H ;
 wire \mprj_pads.area2_io_pad[1]__HLD_H_N ;
 wire \mprj_pads.area2_io_pad[1]__TIE_LO_ESD ;
 wire \mprj_pads.area2_io_pad[1]__IN_H ;
 wire \mprj_pads.area2_io_pad[11]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area2_io_pad[11]__PAD_A_NOESD_H ;
 wire \mprj_pads.area2_io_pad[11]__HLD_H_N ;
 wire \mprj_pads.area2_io_pad[11]__TIE_LO_ESD ;
 wire \mprj_pads.area2_io_pad[11]__IN_H ;
 wire \mprj_pads.area1_io_pad[18]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area1_io_pad[18]__PAD_A_NOESD_H ;
 wire \mprj_pads.area1_io_pad[18]__HLD_H_N ;
 wire \mprj_pads.area1_io_pad[18]__TIE_LO_ESD ;
 wire \mprj_pads.area1_io_pad[18]__IN_H ;
 wire \mprj_pads.area1_io_pad[3]__TIE_LO_ESD ;
 wire \mprj_pads.area1_io_pad[3]__HLD_H_N ;
 wire \mprj_pads.area1_io_pad[3]__PAD_A_ESD_0_H ;
 wire \mprj_pads.area1_io_pad[3]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area1_io_pad[3]__PAD_A_NOESD_H ;
 wire \mprj_pads.area1_io_pad[3]__IN_H ;
 wire \mprj_pads.area2_io_pad[3]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area2_io_pad[3]__PAD_A_NOESD_H ;
 wire \mprj_pads.area2_io_pad[3]__HLD_H_N ;
 wire \mprj_pads.area2_io_pad[3]__TIE_LO_ESD ;
 wire \mprj_pads.area2_io_pad[3]__IN_H ;
 wire \mprj_pads.area2_io_pad[13]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area2_io_pad[13]__PAD_A_NOESD_H ;
 wire \mprj_pads.area2_io_pad[13]__HLD_H_N ;
 wire \mprj_pads.area2_io_pad[13]__TIE_LO_ESD ;
 wire \mprj_pads.area2_io_pad[13]__IN_H ;
 wire constant_block_6__one;
 wire \mprj_pads.area1_io_pad[5]__TIE_LO_ESD ;
 wire \mprj_pads.area1_io_pad[5]__HLD_H_N ;
 wire \mprj_pads.area1_io_pad[5]__PAD_A_ESD_0_H ;
 wire \mprj_pads.area1_io_pad[5]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area1_io_pad[5]__PAD_A_NOESD_H ;
 wire \mprj_pads.area1_io_pad[5]__IN_H ;
 wire \mprj_pads.area2_io_pad[5]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area2_io_pad[5]__PAD_A_NOESD_H ;
 wire \mprj_pads.area2_io_pad[5]__HLD_H_N ;
 wire \mprj_pads.area2_io_pad[5]__TIE_LO_ESD ;
 wire \mprj_pads.area2_io_pad[5]__IN_H ;
 wire constant_block_5__one;
 wire \mprj_pads.area2_io_pad[15]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area2_io_pad[15]__PAD_A_NOESD_H ;
 wire \mprj_pads.area2_io_pad[15]__HLD_H_N ;
 wire \mprj_pads.area2_io_pad[15]__TIE_LO_ESD ;
 wire \mprj_pads.area2_io_pad[15]__IN_H ;
 wire constant_block_4__one;
 wire \mprj_pads.area1_io_pad[11]__TIE_LO_ESD ;
 wire \mprj_pads.area1_io_pad[11]__HLD_H_N ;
 wire \mprj_pads.area1_io_pad[11]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area1_io_pad[11]__PAD_A_NOESD_H ;
 wire \mprj_pads.area1_io_pad[11]__IN_H ;
 wire \mprj_pads.area1_io_pad[7]__TIE_LO_ESD ;
 wire \mprj_pads.area1_io_pad[7]__HLD_H_N ;
 wire \mprj_pads.area1_io_pad[7]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area1_io_pad[7]__PAD_A_NOESD_H ;
 wire \mprj_pads.area1_io_pad[7]__IN_H ;
 wire \mprj_pads.area2_io_pad[7]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area2_io_pad[7]__PAD_A_NOESD_H ;
 wire \mprj_pads.area2_io_pad[7]__HLD_H_N ;
 wire \mprj_pads.area2_io_pad[7]__TIE_LO_ESD ;
 wire \mprj_pads.area2_io_pad[7]__IN_H ;
 wire \mprj_pads.area2_io_pad[17]__PAD_A_ESD_0_H ;
 wire \mprj_pads.area2_io_pad[17]__PAD_A_ESD_1_H ;
 wire \mprj_pads.area2_io_pad[17]__PAD_A_NOESD_H ;
 wire \mprj_pads.area2_io_pad[17]__HLD_H_N ;
 wire \mprj_pads.area2_io_pad[17]__TIE_LO_ESD ;
 wire \mprj_pads.area2_io_pad[17]__IN_H ;
 wire clock_pad__TIE_LO_ESD;
 wire clock_pad__HLD_H_N;
 wire clock_pad__OUT;
 wire clock_pad__PAD_A_ESD_0_H;
 wire clock_pad__PAD_A_ESD_1_H;
 wire clock_pad__PAD_A_NOESD_H;
 wire clock_pad__IN_H;
 wire [2:0] flash_clk_pad__DM;
 wire [2:0] flash_csb_pad__DM;

 sky130_ef_io__com_bus_slice_20um FILLER_170 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_374 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__corner_pad \mgmt_corner[0]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_10um FILLER_171 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_172 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_174 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_173 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_3 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_2 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_1 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_6 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_5 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_4 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_181 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__vssa_hvc_clamped_pad mgmt_vssa_hvclamp_pad (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA_PAD(vssa_pad),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_10um FILLER_182 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_183 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_185 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_184 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_187 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_10um FILLER_188 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_189 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_191 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_190 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_7 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_8 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_9 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_10 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_11 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_12 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_198 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_fd_io__top_xres4v2 resetb_pad (.PAD_A_ESD_H(xresloop),
    .XRES_H_N(resetb_core_h),
    .FILT_IN_H(xres_vss_loop),
    .ENABLE_VDDIO(constant_block_0__one),
    .TIE_WEAK_HI_H(xresloop),
    .ENABLE_H(porb_h),
    .PULLUP_H(xres_vss_loop),
    .EN_VDDIO_SIG_H(xres_vss_loop),
    .TIE_LO_ESD(xres_vss_loop),
    .TIE_HI_ESD(resetb_pad__TIE_HI_ESD),
    .DISABLE_PULLUP_H(xres_vss_loop),
    .INP_SEL_H(xres_vss_loop),
    .VSSIO(vssio),
    .VSSA(vssa),
    .VSSD(vssd),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VDDIO(vddio),
    .VSWITCH(vddio),
    .VDDA(vdda),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .PAD(resetb));
 sky130_ef_io__com_bus_slice_10um FILLER_199 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_200 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_202 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_201 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 constant_block constant_block_0 (.one(constant_block_0__one),
    .vccd(vccd),
    .vssd(vssd),
    .zero(constant_block_0__zero));
 sky130_ef_io__com_bus_slice_10um FILLER_205 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_206 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_208 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_207 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_13 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_204 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_16 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_15 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_14 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_10um FILLER_216 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_18 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_17 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_215 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped clock_pad (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(clock_pad__OUT),
    .ANALOG_POL(clock_pad__OUT),
    .ANALOG_SEL(clock_pad__OUT),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(clock_pad__TIE_LO_ESD),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(clock_pad__OE_N),
    .ENABLE_VSWITCH_H(clock_pad__TIE_LO_ESD),
    .HLD_H_N(clock_pad__HLD_H_N),
    .HLD_OVR(clock_pad__OUT),
    .IB_MODE_SEL(clock_pad__OUT),
    .IN(clock_core),
    .IN_H(clock_pad__IN_H),
    .INP_DIS(por),
    .OE_N(clock_pad__OE_N),
    .OUT(clock_pad__OUT),
    .PAD(clock),
    .PAD_A_ESD_0_H(clock_pad__PAD_A_ESD_0_H),
    .PAD_A_ESD_1_H(clock_pad__PAD_A_ESD_1_H),
    .PAD_A_NOESD_H(clock_pad__PAD_A_NOESD_H),
    .SLOW(clock_pad__OUT),
    .TIE_HI_ESD(clock_pad__HLD_H_N),
    .TIE_LO_ESD(clock_pad__TIE_LO_ESD),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(clock_pad__OUT),
    .DM({clock_pad__OUT,
    clock_pad__OUT,
    clock_pad__OE_N}));
 sky130_ef_io__com_bus_slice_5um FILLER_217 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_219 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_218 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 constant_block constant_block_1 (.one(clock_pad__OE_N),
    .vccd(vccd),
    .vssd(vssd),
    .zero(clock_pad__OUT));
 sky130_ef_io__com_bus_slice_10um FILLER_222 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_223 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_225 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_224 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_19 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_221 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_23 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_22 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_21 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_20 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__vssd_lvc_clamped_pad mgmt_vssd_lvclamp_pad (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSD_PAD(vssd_pad),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_10um FILLER_233 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_234 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_236 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_235 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_24 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_232 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_10um FILLER_239 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_240 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_242 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_241 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_26 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_25 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_238 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_30 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_29 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_28 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_27 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped flash_csb_pad (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(flash_csb_pad__SLOW),
    .ANALOG_POL(flash_csb_pad__SLOW),
    .ANALOG_SEL(flash_csb_pad__SLOW),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(flash_csb_pad__TIE_LO_ESD),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(flash_csb_pad__DM[2]),
    .ENABLE_VSWITCH_H(flash_csb_pad__TIE_LO_ESD),
    .HLD_H_N(flash_csb_pad__HLD_H_N),
    .HLD_OVR(flash_csb_pad__SLOW),
    .IB_MODE_SEL(flash_csb_pad__SLOW),
    .IN(flash_csb_pad__IN),
    .IN_H(flash_csb_pad__IN_H),
    .INP_DIS(flash_csb_pad__SLOW),
    .OE_N(flash_csb_oeb_core),
    .OUT(flash_csb_core),
    .PAD(flash_csb),
    .PAD_A_ESD_0_H(flash_csb_pad__PAD_A_ESD_0_H),
    .PAD_A_ESD_1_H(flash_csb_pad__PAD_A_ESD_1_H),
    .PAD_A_NOESD_H(flash_csb_pad__PAD_A_NOESD_H),
    .SLOW(flash_csb_pad__SLOW),
    .TIE_HI_ESD(flash_csb_pad__HLD_H_N),
    .TIE_LO_ESD(flash_csb_pad__TIE_LO_ESD),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(flash_csb_pad__SLOW),
    .DM({flash_csb_pad__DM[2],
    flash_csb_pad__DM[2],
    flash_csb_pad__SLOW}));
 sky130_ef_io__com_bus_slice_10um FILLER_250 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_251 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_253 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_252 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_249 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_255 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 constant_block constant_block_2 (.one(flash_csb_pad__DM[2]),
    .vccd(vccd),
    .vssd(vssd),
    .zero(flash_csb_pad__SLOW));
 sky130_ef_io__com_bus_slice_10um FILLER_256 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_257 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_259 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_258 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_31 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_32 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_33 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_34 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_35 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped flash_clk_pad (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(flash_clk_pad__SLOW),
    .ANALOG_POL(flash_clk_pad__SLOW),
    .ANALOG_SEL(flash_clk_pad__SLOW),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(flash_clk_pad__TIE_LO_ESD),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(flash_clk_pad__DM[2]),
    .ENABLE_VSWITCH_H(flash_clk_pad__TIE_LO_ESD),
    .HLD_H_N(flash_clk_pad__HLD_H_N),
    .HLD_OVR(flash_clk_pad__SLOW),
    .IB_MODE_SEL(flash_clk_pad__SLOW),
    .IN(flash_clk_pad__IN),
    .IN_H(flash_clk_pad__IN_H),
    .INP_DIS(flash_clk_pad__SLOW),
    .OE_N(flash_clk_oeb_core),
    .OUT(flash_clk_core),
    .PAD(flash_clk),
    .PAD_A_ESD_0_H(flash_clk_pad__PAD_A_ESD_0_H),
    .PAD_A_ESD_1_H(flash_clk_pad__PAD_A_ESD_1_H),
    .PAD_A_NOESD_H(flash_clk_pad__PAD_A_NOESD_H),
    .SLOW(flash_clk_pad__SLOW),
    .TIE_HI_ESD(flash_clk_pad__HLD_H_N),
    .TIE_LO_ESD(flash_clk_pad__TIE_LO_ESD),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(flash_clk_pad__SLOW),
    .DM({flash_clk_pad__DM[2],
    flash_clk_pad__DM[2],
    flash_clk_pad__SLOW}));
 sky130_ef_io__com_bus_slice_10um FILLER_267 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_268 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_270 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_269 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_36 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_266 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 constant_block constant_block_3 (.one(flash_clk_pad__DM[2]),
    .vccd(vccd),
    .vssd(vssd),
    .zero(flash_clk_pad__SLOW));
 sky130_ef_io__com_bus_slice_20um FILLER_272 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_10um FILLER_273 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_274 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_276 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_275 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_38 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_37 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_42 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_41 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_40 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_39 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped flash_io0_pad (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(flash_io0_pad__SLOW),
    .ANALOG_POL(flash_io0_pad__SLOW),
    .ANALOG_SEL(flash_io0_pad__SLOW),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(flash_io0_pad__TIE_LO_ESD),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(constant_block_4__one),
    .ENABLE_VSWITCH_H(flash_io0_pad__TIE_LO_ESD),
    .HLD_H_N(flash_io0_pad__HLD_H_N),
    .HLD_OVR(flash_io0_pad__SLOW),
    .IB_MODE_SEL(flash_io0_pad__SLOW),
    .IN(flash_io0_di_core),
    .IN_H(flash_io0_pad__IN_H),
    .INP_DIS(flash_io0_ieb_core),
    .OE_N(flash_io0_oeb_core),
    .OUT(flash_io0_do_core),
    .PAD(flash_io0),
    .PAD_A_ESD_0_H(flash_io0_pad__PAD_A_ESD_0_H),
    .PAD_A_ESD_1_H(flash_io0_pad__PAD_A_ESD_1_H),
    .PAD_A_NOESD_H(flash_io0_pad__PAD_A_NOESD_H),
    .SLOW(flash_io0_pad__SLOW),
    .TIE_HI_ESD(flash_io0_pad__HLD_H_N),
    .TIE_LO_ESD(flash_io0_pad__TIE_LO_ESD),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(flash_io0_pad__SLOW),
    .DM({flash_io0_ieb_core,
    flash_io0_ieb_core,
    flash_io0_oeb_core}));
 sky130_ef_io__com_bus_slice_10um FILLER_284 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_285 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_287 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_286 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_283 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_289 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 constant_block constant_block_4 (.one(constant_block_4__one),
    .vccd(vccd),
    .vssd(vssd),
    .zero(flash_io0_pad__SLOW));
 sky130_ef_io__com_bus_slice_10um FILLER_290 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_291 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_293 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_292 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_45 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_44 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_43 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_48 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_47 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_46 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_300 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped flash_io1_pad (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(flash_io1_pad__SLOW),
    .ANALOG_POL(flash_io1_pad__SLOW),
    .ANALOG_SEL(flash_io1_pad__SLOW),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(flash_io1_pad__TIE_LO_ESD),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(constant_block_5__one),
    .ENABLE_VSWITCH_H(flash_io1_pad__TIE_LO_ESD),
    .HLD_H_N(flash_io1_pad__HLD_H_N),
    .HLD_OVR(flash_io1_pad__SLOW),
    .IB_MODE_SEL(flash_io1_pad__SLOW),
    .IN(flash_io1_di_core),
    .IN_H(flash_io1_pad__IN_H),
    .INP_DIS(flash_io1_ieb_core),
    .OE_N(flash_io1_oeb_core),
    .OUT(flash_io1_do_core),
    .PAD(flash_io1),
    .PAD_A_ESD_0_H(flash_io1_pad__PAD_A_ESD_0_H),
    .PAD_A_ESD_1_H(flash_io1_pad__PAD_A_ESD_1_H),
    .PAD_A_NOESD_H(flash_io1_pad__PAD_A_NOESD_H),
    .SLOW(flash_io1_pad__SLOW),
    .TIE_HI_ESD(flash_io1_pad__HLD_H_N),
    .TIE_LO_ESD(flash_io1_pad__TIE_LO_ESD),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(flash_io1_pad__SLOW),
    .DM({flash_io1_ieb_core,
    flash_io1_ieb_core,
    flash_io1_oeb_core}));
 sky130_ef_io__com_bus_slice_10um FILLER_301 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_302 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_304 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_303 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_306 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 constant_block constant_block_5 (.one(constant_block_5__one),
    .vccd(vccd),
    .vssd(vssd),
    .zero(flash_io1_pad__SLOW));
 sky130_ef_io__com_bus_slice_10um FILLER_307 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_308 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_310 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_309 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_49 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_50 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_51 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_52 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_53 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_54 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped gpio_pad (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(gpio_pad__SLOW),
    .ANALOG_POL(gpio_pad__SLOW),
    .ANALOG_SEL(gpio_pad__SLOW),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(gpio_pad__TIE_LO_ESD),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(constant_block_6__one),
    .ENABLE_VSWITCH_H(gpio_pad__TIE_LO_ESD),
    .HLD_H_N(gpio_pad__HLD_H_N),
    .HLD_OVR(gpio_pad__SLOW),
    .IB_MODE_SEL(gpio_pad__SLOW),
    .IN(gpio_in_core),
    .IN_H(gpio_pad__IN_H),
    .INP_DIS(gpio_inenb_core),
    .OE_N(gpio_outenb_core),
    .OUT(gpio_out_core),
    .PAD(gpio),
    .PAD_A_ESD_0_H(gpio_pad__PAD_A_ESD_0_H),
    .PAD_A_ESD_1_H(gpio_pad__PAD_A_ESD_1_H),
    .PAD_A_NOESD_H(gpio_pad__PAD_A_NOESD_H),
    .SLOW(gpio_pad__SLOW),
    .TIE_HI_ESD(gpio_pad__HLD_H_N),
    .TIE_LO_ESD(gpio_pad__TIE_LO_ESD),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(gpio_pad__SLOW),
    .DM({gpio_mode1_core,
    gpio_mode1_core,
    gpio_mode0_core}));
 sky130_ef_io__com_bus_slice_10um FILLER_318 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_319 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_321 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_320 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_317 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 constant_block constant_block_6 (.one(constant_block_6__one),
    .vccd(vccd),
    .vssd(vssd),
    .zero(gpio_pad__SLOW));
 sky130_ef_io__com_bus_slice_10um FILLER_324 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_325 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_327 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_326 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_55 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_323 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_57 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_56 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_60 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_59 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_58 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_334 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__vssio_hvc_clamped_pad \mgmt_vssio_hvclamp_pad[0]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSIO_PAD(vssio_pad),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_10um FILLER_335 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_336 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_338 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_337 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_10um FILLER_341 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_342 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_340 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_344 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_343 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_64 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_63 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_62 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_61 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_10um FILLER_352 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_66 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_65 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_351 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__vdda_hvc_clamped_pad mgmt_vdda_hvclamp_pad (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VDDA_PAD(vdda_pad),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_353 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_355 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_354 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_357 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_10um FILLER_358 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_359 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_360 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_361 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_67 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_68 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_69 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_70 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_71 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um bus_tie_72 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_368 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_10um FILLER_369 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_605 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__corner_pad \mgmt_corner[1]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_371 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_372 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_373 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_370 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_378 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_377 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_376 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_375 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__vccd_lvc_clamped_pad mgmt_vccd_lvclamp_pad (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VCCD_PAD(vccd_pad),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_10um FILLER_380 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_381 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_382 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_379 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_384 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_606 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_607 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_608 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_609 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_610 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_611 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__disconnect_vdda_slice_5um disconnect_vdda_1 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_SB1 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_612 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_615 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_616 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_617 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_618 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_388 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_387 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_386 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_385 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__vddio_hvc_clamped_pad \mgmt_vddio_hvclamp_pad[0]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VDDIO_PAD(vddio_pad),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_10um FILLER_390 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_391 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_392 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_389 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_394 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_619 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_620 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_621 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_624 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_625 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_626 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_622 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area1_io_pad[0]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[0]),
    .ANALOG_POL(mprj_io_analog_pol[0]),
    .ANALOG_SEL(mprj_io_analog_sel[0]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area1_io_pad[0]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[0]),
    .ENABLE_VSWITCH_H(\mprj_pads.area1_io_pad[0]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area1_io_pad[0]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[0]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[0]),
    .IN(mprj_io_in[0]),
    .IN_H(\mprj_pads.area1_io_pad[0]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[0]),
    .OE_N(mprj_io_oeb[0]),
    .OUT(mprj_io_out[0]),
    .PAD(mprj_io[0]),
    .PAD_A_ESD_0_H(\mprj_pads.area1_io_pad[0]__PAD_A_ESD_0_H ),
    .PAD_A_ESD_1_H(\mprj_pads.area1_io_pad[0]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area1_io_pad[0]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[0]),
    .TIE_HI_ESD(\mprj_pads.area1_io_pad[0]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area1_io_pad[0]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda1),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa1),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[0]),
    .DM({mprj_io_dm[2],
    mprj_io_dm[1],
    mprj_io_dm[0]}));
 sky130_ef_io__com_bus_slice_20um FILLER_395 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_396 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_397 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_398 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_399 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_10um FILLER_400 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__disconnect_vdda_slice_5um disconnect_vdda_2 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_SB2 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_401 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_402 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa),
    .VDDA(vdda),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_405 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_406 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_407 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_408 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_627 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_628 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_629 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_630 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_632 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_631 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area1_io_pad[1]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[1]),
    .ANALOG_POL(mprj_io_analog_pol[1]),
    .ANALOG_SEL(mprj_io_analog_sel[1]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area1_io_pad[1]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[1]),
    .ENABLE_VSWITCH_H(\mprj_pads.area1_io_pad[1]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area1_io_pad[1]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[1]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[1]),
    .IN(mprj_io_in[1]),
    .IN_H(\mprj_pads.area1_io_pad[1]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[1]),
    .OE_N(mprj_io_oeb[1]),
    .OUT(mprj_io_out[1]),
    .PAD(mprj_io[1]),
    .PAD_A_ESD_0_H(\mprj_pads.area1_io_pad[1]__PAD_A_ESD_0_H ),
    .PAD_A_ESD_1_H(\mprj_pads.area1_io_pad[1]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area1_io_pad[1]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[1]),
    .TIE_HI_ESD(\mprj_pads.area1_io_pad[1]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area1_io_pad[1]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda1),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa1),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[1]),
    .DM({mprj_io_dm[5],
    mprj_io_dm[4],
    mprj_io_dm[3]}));
 sky130_ef_io__com_bus_slice_20um FILLER_634 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_635 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area2_io_pad[18]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[37]),
    .ANALOG_POL(mprj_io_analog_pol[37]),
    .ANALOG_SEL(mprj_io_analog_sel[37]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area2_io_pad[18]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[37]),
    .ENABLE_VSWITCH_H(\mprj_pads.area2_io_pad[18]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area2_io_pad[18]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[37]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[37]),
    .IN(mprj_io_in[37]),
    .IN_H(\mprj_pads.area2_io_pad[18]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[37]),
    .OE_N(mprj_io_oeb[37]),
    .OUT(mprj_io_out[37]),
    .PAD(mprj_io[37]),
    .PAD_A_ESD_0_H(\mprj_pads.area2_io_pad[18]__PAD_A_ESD_0_H ),
    .PAD_A_ESD_1_H(\mprj_pads.area2_io_pad[18]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area2_io_pad[18]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[37]),
    .TIE_HI_ESD(\mprj_pads.area2_io_pad[18]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area2_io_pad[18]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda2),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa2),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[37]),
    .DM({mprj_io_dm[113],
    mprj_io_dm[112],
    mprj_io_dm[111]}));
 sky130_ef_io__com_bus_slice_10um FILLER_411 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_412 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_413 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_410 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_409 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_415 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_418 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_417 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_416 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_636 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_637 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_638 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_639 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_640 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_641 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area1_io_pad[2]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[2]),
    .ANALOG_POL(mprj_io_analog_pol[2]),
    .ANALOG_SEL(mprj_io_analog_sel[2]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area1_io_pad[2]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[2]),
    .ENABLE_VSWITCH_H(\mprj_pads.area1_io_pad[2]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area1_io_pad[2]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[2]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[2]),
    .IN(mprj_io_in[2]),
    .IN_H(\mprj_pads.area1_io_pad[2]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[2]),
    .OE_N(mprj_io_oeb[2]),
    .OUT(mprj_io_out[2]),
    .PAD(mprj_io[2]),
    .PAD_A_ESD_0_H(\mprj_pads.area1_io_pad[2]__PAD_A_ESD_0_H ),
    .PAD_A_ESD_1_H(\mprj_pads.area1_io_pad[2]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area1_io_pad[2]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[2]),
    .TIE_HI_ESD(\mprj_pads.area1_io_pad[2]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area1_io_pad[2]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda1),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa1),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[2]),
    .DM({mprj_io_dm[8],
    mprj_io_dm[7],
    mprj_io_dm[6]}));
 sky130_ef_io__com_bus_slice_20um FILLER_643 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_644 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area2_io_pad[17]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[36]),
    .ANALOG_POL(mprj_io_analog_pol[36]),
    .ANALOG_SEL(mprj_io_analog_sel[36]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area2_io_pad[17]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[36]),
    .ENABLE_VSWITCH_H(\mprj_pads.area2_io_pad[17]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area2_io_pad[17]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[36]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[36]),
    .IN(mprj_io_in[36]),
    .IN_H(\mprj_pads.area2_io_pad[17]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[36]),
    .OE_N(mprj_io_oeb[36]),
    .OUT(mprj_io_out[36]),
    .PAD(mprj_io[36]),
    .PAD_A_ESD_0_H(\mprj_pads.area2_io_pad[17]__PAD_A_ESD_0_H ),
    .PAD_A_ESD_1_H(\mprj_pads.area2_io_pad[17]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area2_io_pad[17]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[36]),
    .TIE_HI_ESD(\mprj_pads.area2_io_pad[17]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area2_io_pad[17]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda2),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa2),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[36]),
    .DM({mprj_io_dm[110],
    mprj_io_dm[109],
    mprj_io_dm[108]}));
 sky130_ef_io__com_bus_slice_10um FILLER_421 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_422 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_423 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_420 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_419 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_425 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_428 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_427 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_426 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_645 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_646 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_647 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_648 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_649 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_651 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_650 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area1_io_pad[3]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[3]),
    .ANALOG_POL(mprj_io_analog_pol[3]),
    .ANALOG_SEL(mprj_io_analog_sel[3]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area1_io_pad[3]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[3]),
    .ENABLE_VSWITCH_H(\mprj_pads.area1_io_pad[3]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area1_io_pad[3]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[3]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[3]),
    .IN(mprj_io_in[3]),
    .IN_H(\mprj_pads.area1_io_pad[3]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[3]),
    .OE_N(mprj_io_oeb[3]),
    .OUT(mprj_io_out[3]),
    .PAD(mprj_io[3]),
    .PAD_A_ESD_0_H(\mprj_pads.area1_io_pad[3]__PAD_A_ESD_0_H ),
    .PAD_A_ESD_1_H(\mprj_pads.area1_io_pad[3]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area1_io_pad[3]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[3]),
    .TIE_HI_ESD(\mprj_pads.area1_io_pad[3]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area1_io_pad[3]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda1),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa1),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[3]),
    .DM({mprj_io_dm[11],
    mprj_io_dm[10],
    mprj_io_dm[9]}));
 sky130_ef_io__com_bus_slice_20um FILLER_653 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_429 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_430 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_433 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_432 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_10um FILLER_431 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area2_io_pad[16]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[35]),
    .ANALOG_POL(mprj_io_analog_pol[35]),
    .ANALOG_SEL(mprj_io_analog_sel[35]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area2_io_pad[16]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[35]),
    .ENABLE_VSWITCH_H(\mprj_pads.area2_io_pad[16]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area2_io_pad[16]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[35]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[35]),
    .IN(mprj_io_in[35]),
    .IN_H(\mprj_pads.area2_io_pad[16]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[35]),
    .OE_N(mprj_io_oeb[35]),
    .OUT(mprj_io_out[35]),
    .PAD(mprj_io[35]),
    .PAD_A_ESD_0_H(mprj_analog_io[28]),
    .PAD_A_ESD_1_H(\mprj_pads.area2_io_pad[16]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area2_io_pad[16]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[35]),
    .TIE_HI_ESD(\mprj_pads.area2_io_pad[16]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area2_io_pad[16]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda2),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa2),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[35]),
    .DM({mprj_io_dm[107],
    mprj_io_dm[106],
    mprj_io_dm[105]}));
 sky130_ef_io__com_bus_slice_20um FILLER_435 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_436 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_437 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_654 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_655 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_656 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_657 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_658 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_659 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_660 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area1_io_pad[4]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[4]),
    .ANALOG_POL(mprj_io_analog_pol[4]),
    .ANALOG_SEL(mprj_io_analog_sel[4]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area1_io_pad[4]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[4]),
    .ENABLE_VSWITCH_H(\mprj_pads.area1_io_pad[4]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area1_io_pad[4]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[4]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[4]),
    .IN(mprj_io_in[4]),
    .IN_H(\mprj_pads.area1_io_pad[4]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[4]),
    .OE_N(mprj_io_oeb[4]),
    .OUT(mprj_io_out[4]),
    .PAD(mprj_io[4]),
    .PAD_A_ESD_0_H(\mprj_pads.area1_io_pad[4]__PAD_A_ESD_0_H ),
    .PAD_A_ESD_1_H(\mprj_pads.area1_io_pad[4]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area1_io_pad[4]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[4]),
    .TIE_HI_ESD(\mprj_pads.area1_io_pad[4]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area1_io_pad[4]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda1),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa1),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[4]),
    .DM({mprj_io_dm[14],
    mprj_io_dm[13],
    mprj_io_dm[12]}));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area2_io_pad[15]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[34]),
    .ANALOG_POL(mprj_io_analog_pol[34]),
    .ANALOG_SEL(mprj_io_analog_sel[34]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area2_io_pad[15]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[34]),
    .ENABLE_VSWITCH_H(\mprj_pads.area2_io_pad[15]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area2_io_pad[15]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[34]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[34]),
    .IN(mprj_io_in[34]),
    .IN_H(\mprj_pads.area2_io_pad[15]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[34]),
    .OE_N(mprj_io_oeb[34]),
    .OUT(mprj_io_out[34]),
    .PAD(mprj_io[34]),
    .PAD_A_ESD_0_H(mprj_analog_io[27]),
    .PAD_A_ESD_1_H(\mprj_pads.area2_io_pad[15]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area2_io_pad[15]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[34]),
    .TIE_HI_ESD(\mprj_pads.area2_io_pad[15]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area2_io_pad[15]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda2),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa2),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[34]),
    .DM({mprj_io_dm[104],
    mprj_io_dm[103],
    mprj_io_dm[102]}));
 sky130_ef_io__com_bus_slice_10um FILLER_441 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_442 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_443 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_440 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_439 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_438 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_445 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_447 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_446 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_662 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_663 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_664 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_665 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_666 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_667 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_668 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_669 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area1_io_pad[5]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[5]),
    .ANALOG_POL(mprj_io_analog_pol[5]),
    .ANALOG_SEL(mprj_io_analog_sel[5]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area1_io_pad[5]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[5]),
    .ENABLE_VSWITCH_H(\mprj_pads.area1_io_pad[5]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area1_io_pad[5]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[5]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[5]),
    .IN(mprj_io_in[5]),
    .IN_H(\mprj_pads.area1_io_pad[5]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[5]),
    .OE_N(mprj_io_oeb[5]),
    .OUT(mprj_io_out[5]),
    .PAD(mprj_io[5]),
    .PAD_A_ESD_0_H(\mprj_pads.area1_io_pad[5]__PAD_A_ESD_0_H ),
    .PAD_A_ESD_1_H(\mprj_pads.area1_io_pad[5]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area1_io_pad[5]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[5]),
    .TIE_HI_ESD(\mprj_pads.area1_io_pad[5]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area1_io_pad[5]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda1),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa1),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[5]),
    .DM({mprj_io_dm[17],
    mprj_io_dm[16],
    mprj_io_dm[15]}));
 sky130_ef_io__com_bus_slice_10um FILLER_451 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_452 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_450 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_449 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_448 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area2_io_pad[14]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[33]),
    .ANALOG_POL(mprj_io_analog_pol[33]),
    .ANALOG_SEL(mprj_io_analog_sel[33]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area2_io_pad[14]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[33]),
    .ENABLE_VSWITCH_H(\mprj_pads.area2_io_pad[14]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area2_io_pad[14]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[33]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[33]),
    .IN(mprj_io_in[33]),
    .IN_H(\mprj_pads.area2_io_pad[14]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[33]),
    .OE_N(mprj_io_oeb[33]),
    .OUT(mprj_io_out[33]),
    .PAD(mprj_io[33]),
    .PAD_A_ESD_0_H(mprj_analog_io[26]),
    .PAD_A_ESD_1_H(\mprj_pads.area2_io_pad[14]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area2_io_pad[14]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[33]),
    .TIE_HI_ESD(\mprj_pads.area2_io_pad[14]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area2_io_pad[14]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda2),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa2),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[33]),
    .DM({mprj_io_dm[101],
    mprj_io_dm[100],
    mprj_io_dm[99]}));
 sky130_ef_io__com_bus_slice_1um FILLER_453 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_457 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_456 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_455 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_674 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_673 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_672 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_671 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_678 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_677 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_676 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_675 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area1_io_pad[6]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[6]),
    .ANALOG_POL(mprj_io_analog_pol[6]),
    .ANALOG_SEL(mprj_io_analog_sel[6]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area1_io_pad[6]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[6]),
    .ENABLE_VSWITCH_H(\mprj_pads.area1_io_pad[6]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area1_io_pad[6]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[6]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[6]),
    .IN(mprj_io_in[6]),
    .IN_H(\mprj_pads.area1_io_pad[6]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[6]),
    .OE_N(mprj_io_oeb[6]),
    .OUT(mprj_io_out[6]),
    .PAD(mprj_io[6]),
    .PAD_A_ESD_0_H(\mprj_pads.area1_io_pad[6]__PAD_A_ESD_0_H ),
    .PAD_A_ESD_1_H(\mprj_pads.area1_io_pad[6]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area1_io_pad[6]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[6]),
    .TIE_HI_ESD(\mprj_pads.area1_io_pad[6]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area1_io_pad[6]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda1),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa1),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[6]),
    .DM({mprj_io_dm[20],
    mprj_io_dm[19],
    mprj_io_dm[18]}));
 sky130_ef_io__com_bus_slice_1um FILLER_679 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_10um FILLER_461 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_460 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_459 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_458 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area2_io_pad[13]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[32]),
    .ANALOG_POL(mprj_io_analog_pol[32]),
    .ANALOG_SEL(mprj_io_analog_sel[32]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area2_io_pad[13]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[32]),
    .ENABLE_VSWITCH_H(\mprj_pads.area2_io_pad[13]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area2_io_pad[13]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[32]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[32]),
    .IN(mprj_io_in[32]),
    .IN_H(\mprj_pads.area2_io_pad[13]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[32]),
    .OE_N(mprj_io_oeb[32]),
    .OUT(mprj_io_out[32]),
    .PAD(mprj_io[32]),
    .PAD_A_ESD_0_H(mprj_analog_io[25]),
    .PAD_A_ESD_1_H(\mprj_pads.area2_io_pad[13]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area2_io_pad[13]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[32]),
    .TIE_HI_ESD(\mprj_pads.area2_io_pad[13]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area2_io_pad[13]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda2),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa2),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[32]),
    .DM({mprj_io_dm[98],
    mprj_io_dm[97],
    mprj_io_dm[96]}));
 sky130_ef_io__com_bus_slice_5um FILLER_462 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_463 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_467 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_466 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_465 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_681 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_682 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_683 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_684 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_685 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_686 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_687 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_688 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__vssa_hvc_clamped_pad \user1_vssa_hvclamp_pad[1]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA_PAD(vssa1_pad2),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_10um FILLER_471 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_470 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_469 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_468 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__vssd_lvc_clamped3_pad user2_vssd_lvclamp_pad (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSD_PAD(vssd2_pad),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSSD1(vssd2),
    .VCCD1(vccd2));
 sky130_ef_io__com_bus_slice_5um FILLER_472 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_473 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_475 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_477 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_476 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_692 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_691 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_690 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_696 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_695 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_694 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_693 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__vssd_lvc_clamped3_pad user1_vssd_lvclamp_pad (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSD_PAD(vssd1_pad),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSSD1(vssd1),
    .VCCD1(vccd1));
 sky130_ef_io__com_bus_slice_5um FILLER_697 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_698 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_480 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_479 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_478 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__vdda_hvc_clamped_pad user2_vdda_hvclamp_pad (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VDDA_PAD(vdda2_pad),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_10um FILLER_481 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_482 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_483 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_487 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_486 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_485 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_700 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_701 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_702 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_703 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_704 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_705 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_706 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_707 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__vdda_hvc_clamped_pad \user1_vdda_hvclamp_pad[1]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VDDA_PAD(vdda1_pad2),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_488 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_489 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_490 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_10um FILLER_491 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_493 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_492 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area2_io_pad[12]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[31]),
    .ANALOG_POL(mprj_io_analog_pol[31]),
    .ANALOG_SEL(mprj_io_analog_sel[31]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area2_io_pad[12]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[31]),
    .ENABLE_VSWITCH_H(\mprj_pads.area2_io_pad[12]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area2_io_pad[12]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[31]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[31]),
    .IN(mprj_io_in[31]),
    .IN_H(\mprj_pads.area2_io_pad[12]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[31]),
    .OE_N(mprj_io_oeb[31]),
    .OUT(mprj_io_out[31]),
    .PAD(mprj_io[31]),
    .PAD_A_ESD_0_H(mprj_analog_io[24]),
    .PAD_A_ESD_1_H(\mprj_pads.area2_io_pad[12]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area2_io_pad[12]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[31]),
    .TIE_HI_ESD(\mprj_pads.area2_io_pad[12]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area2_io_pad[12]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda2),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa2),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[31]),
    .DM({mprj_io_dm[95],
    mprj_io_dm[94],
    mprj_io_dm[93]}));
 sky130_ef_io__com_bus_slice_20um FILLER_495 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_496 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_709 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_710 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_711 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_712 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_713 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_714 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_715 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_716 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area1_io_pad[7]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[7]),
    .ANALOG_POL(mprj_io_analog_pol[7]),
    .ANALOG_SEL(mprj_io_analog_sel[7]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area1_io_pad[7]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[7]),
    .ENABLE_VSWITCH_H(\mprj_pads.area1_io_pad[7]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area1_io_pad[7]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[7]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[7]),
    .IN(mprj_io_in[7]),
    .IN_H(\mprj_pads.area1_io_pad[7]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[7]),
    .OE_N(mprj_io_oeb[7]),
    .OUT(mprj_io_out[7]),
    .PAD(mprj_io[7]),
    .PAD_A_ESD_0_H(mprj_analog_io[0]),
    .PAD_A_ESD_1_H(\mprj_pads.area1_io_pad[7]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area1_io_pad[7]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[7]),
    .TIE_HI_ESD(\mprj_pads.area1_io_pad[7]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area1_io_pad[7]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda1),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa1),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[7]),
    .DM({mprj_io_dm[23],
    mprj_io_dm[22],
    mprj_io_dm[21]}));
 sky130_ef_io__com_bus_slice_20um FILLER_500 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_499 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_498 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_497 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area2_io_pad[11]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[30]),
    .ANALOG_POL(mprj_io_analog_pol[30]),
    .ANALOG_SEL(mprj_io_analog_sel[30]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area2_io_pad[11]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[30]),
    .ENABLE_VSWITCH_H(\mprj_pads.area2_io_pad[11]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area2_io_pad[11]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[30]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[30]),
    .IN(mprj_io_in[30]),
    .IN_H(\mprj_pads.area2_io_pad[11]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[30]),
    .OE_N(mprj_io_oeb[30]),
    .OUT(mprj_io_out[30]),
    .PAD(mprj_io[30]),
    .PAD_A_ESD_0_H(mprj_analog_io[23]),
    .PAD_A_ESD_1_H(\mprj_pads.area2_io_pad[11]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area2_io_pad[11]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[30]),
    .TIE_HI_ESD(\mprj_pads.area2_io_pad[11]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area2_io_pad[11]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda2),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa2),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[30]),
    .DM({mprj_io_dm[92],
    mprj_io_dm[91],
    mprj_io_dm[90]}));
 sky130_ef_io__com_bus_slice_10um FILLER_501 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_502 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_503 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_506 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_505 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_718 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_719 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_720 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_721 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_722 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_723 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_724 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_510 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_509 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_508 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_507 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area2_io_pad[10]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[29]),
    .ANALOG_POL(mprj_io_analog_pol[29]),
    .ANALOG_SEL(mprj_io_analog_sel[29]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area2_io_pad[10]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[29]),
    .ENABLE_VSWITCH_H(\mprj_pads.area2_io_pad[10]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area2_io_pad[10]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[29]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[29]),
    .IN(mprj_io_in[29]),
    .IN_H(\mprj_pads.area2_io_pad[10]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[29]),
    .OE_N(mprj_io_oeb[29]),
    .OUT(mprj_io_out[29]),
    .PAD(mprj_io[29]),
    .PAD_A_ESD_0_H(mprj_analog_io[22]),
    .PAD_A_ESD_1_H(\mprj_pads.area2_io_pad[10]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area2_io_pad[10]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[29]),
    .TIE_HI_ESD(\mprj_pads.area2_io_pad[10]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area2_io_pad[10]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda2),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa2),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[29]),
    .DM({mprj_io_dm[89],
    mprj_io_dm[88],
    mprj_io_dm[87]}));
 sky130_ef_io__com_bus_slice_10um FILLER_511 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_512 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_513 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_516 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_515 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_726 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_725 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area1_io_pad[8]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[8]),
    .ANALOG_POL(mprj_io_analog_pol[8]),
    .ANALOG_SEL(mprj_io_analog_sel[8]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area1_io_pad[8]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[8]),
    .ENABLE_VSWITCH_H(\mprj_pads.area1_io_pad[8]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area1_io_pad[8]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[8]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[8]),
    .IN(mprj_io_in[8]),
    .IN_H(\mprj_pads.area1_io_pad[8]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[8]),
    .OE_N(mprj_io_oeb[8]),
    .OUT(mprj_io_out[8]),
    .PAD(mprj_io[8]),
    .PAD_A_ESD_0_H(mprj_analog_io[1]),
    .PAD_A_ESD_1_H(\mprj_pads.area1_io_pad[8]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area1_io_pad[8]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[8]),
    .TIE_HI_ESD(\mprj_pads.area1_io_pad[8]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area1_io_pad[8]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda1),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa1),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[8]),
    .DM({mprj_io_dm[26],
    mprj_io_dm[25],
    mprj_io_dm[24]}));
 sky130_ef_io__com_bus_slice_20um FILLER_728 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_729 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_730 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_731 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_732 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_733 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_520 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_519 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_518 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_517 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area2_io_pad[9]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[28]),
    .ANALOG_POL(mprj_io_analog_pol[28]),
    .ANALOG_SEL(mprj_io_analog_sel[28]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area2_io_pad[9]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[28]),
    .ENABLE_VSWITCH_H(\mprj_pads.area2_io_pad[9]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area2_io_pad[9]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[28]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[28]),
    .IN(mprj_io_in[28]),
    .IN_H(\mprj_pads.area2_io_pad[9]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[28]),
    .OE_N(mprj_io_oeb[28]),
    .OUT(mprj_io_out[28]),
    .PAD(mprj_io[28]),
    .PAD_A_ESD_0_H(mprj_analog_io[21]),
    .PAD_A_ESD_1_H(\mprj_pads.area2_io_pad[9]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area2_io_pad[9]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[28]),
    .TIE_HI_ESD(\mprj_pads.area2_io_pad[9]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area2_io_pad[9]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda2),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa2),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[28]),
    .DM({mprj_io_dm[86],
    mprj_io_dm[85],
    mprj_io_dm[84]}));
 sky130_ef_io__com_bus_slice_10um FILLER_521 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_522 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_523 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_526 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_525 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_734 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_735 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area1_io_pad[9]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[9]),
    .ANALOG_POL(mprj_io_analog_pol[9]),
    .ANALOG_SEL(mprj_io_analog_sel[9]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area1_io_pad[9]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[9]),
    .ENABLE_VSWITCH_H(\mprj_pads.area1_io_pad[9]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area1_io_pad[9]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[9]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[9]),
    .IN(mprj_io_in[9]),
    .IN_H(\mprj_pads.area1_io_pad[9]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[9]),
    .OE_N(mprj_io_oeb[9]),
    .OUT(mprj_io_out[9]),
    .PAD(mprj_io[9]),
    .PAD_A_ESD_0_H(mprj_analog_io[2]),
    .PAD_A_ESD_1_H(\mprj_pads.area1_io_pad[9]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area1_io_pad[9]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[9]),
    .TIE_HI_ESD(\mprj_pads.area1_io_pad[9]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area1_io_pad[9]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda1),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa1),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[9]),
    .DM({mprj_io_dm[29],
    mprj_io_dm[28],
    mprj_io_dm[27]}));
 sky130_ef_io__com_bus_slice_20um FILLER_737 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_738 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_739 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_740 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_741 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_742 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_527 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_528 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_529 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_530 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_533 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_532 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_10um FILLER_531 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area2_io_pad[8]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[27]),
    .ANALOG_POL(mprj_io_analog_pol[27]),
    .ANALOG_SEL(mprj_io_analog_sel[27]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area2_io_pad[8]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[27]),
    .ENABLE_VSWITCH_H(\mprj_pads.area2_io_pad[8]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area2_io_pad[8]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[27]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[27]),
    .IN(mprj_io_in[27]),
    .IN_H(\mprj_pads.area2_io_pad[8]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[27]),
    .OE_N(mprj_io_oeb[27]),
    .OUT(mprj_io_out[27]),
    .PAD(mprj_io[27]),
    .PAD_A_ESD_0_H(mprj_analog_io[20]),
    .PAD_A_ESD_1_H(\mprj_pads.area2_io_pad[8]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area2_io_pad[8]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[27]),
    .TIE_HI_ESD(\mprj_pads.area2_io_pad[8]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area2_io_pad[8]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda2),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa2),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[27]),
    .DM({mprj_io_dm[83],
    mprj_io_dm[82],
    mprj_io_dm[81]}));
 sky130_ef_io__com_bus_slice_20um FILLER_535 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_743 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_745 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_744 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area1_io_pad[10]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[10]),
    .ANALOG_POL(mprj_io_analog_pol[10]),
    .ANALOG_SEL(mprj_io_analog_sel[10]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area1_io_pad[10]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[10]),
    .ENABLE_VSWITCH_H(\mprj_pads.area1_io_pad[10]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area1_io_pad[10]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[10]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[10]),
    .IN(mprj_io_in[10]),
    .IN_H(\mprj_pads.area1_io_pad[10]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[10]),
    .OE_N(mprj_io_oeb[10]),
    .OUT(mprj_io_out[10]),
    .PAD(mprj_io[10]),
    .PAD_A_ESD_0_H(mprj_analog_io[3]),
    .PAD_A_ESD_1_H(\mprj_pads.area1_io_pad[10]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area1_io_pad[10]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[10]),
    .TIE_HI_ESD(\mprj_pads.area1_io_pad[10]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area1_io_pad[10]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda1),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa1),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[10]),
    .DM({mprj_io_dm[32],
    mprj_io_dm[31],
    mprj_io_dm[30]}));
 sky130_ef_io__com_bus_slice_20um FILLER_747 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_748 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_749 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_750 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_751 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_539 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_538 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_537 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_536 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area2_io_pad[7]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[26]),
    .ANALOG_POL(mprj_io_analog_pol[26]),
    .ANALOG_SEL(mprj_io_analog_sel[26]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area2_io_pad[7]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[26]),
    .ENABLE_VSWITCH_H(\mprj_pads.area2_io_pad[7]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area2_io_pad[7]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[26]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[26]),
    .IN(mprj_io_in[26]),
    .IN_H(\mprj_pads.area2_io_pad[7]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[26]),
    .OE_N(mprj_io_oeb[26]),
    .OUT(mprj_io_out[26]),
    .PAD(mprj_io[26]),
    .PAD_A_ESD_0_H(mprj_analog_io[19]),
    .PAD_A_ESD_1_H(\mprj_pads.area2_io_pad[7]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area2_io_pad[7]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[26]),
    .TIE_HI_ESD(\mprj_pads.area2_io_pad[7]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area2_io_pad[7]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda2),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa2),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[26]),
    .DM({mprj_io_dm[80],
    mprj_io_dm[79],
    mprj_io_dm[78]}));
 sky130_ef_io__com_bus_slice_10um FILLER_541 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_542 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_543 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_540 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_545 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_752 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_753 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_756 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_757 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_758 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_759 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_754 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area1_io_pad[11]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[11]),
    .ANALOG_POL(mprj_io_analog_pol[11]),
    .ANALOG_SEL(mprj_io_analog_sel[11]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area1_io_pad[11]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[11]),
    .ENABLE_VSWITCH_H(\mprj_pads.area1_io_pad[11]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area1_io_pad[11]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[11]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[11]),
    .IN(mprj_io_in[11]),
    .IN_H(\mprj_pads.area1_io_pad[11]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[11]),
    .OE_N(mprj_io_oeb[11]),
    .OUT(mprj_io_out[11]),
    .PAD(mprj_io[11]),
    .PAD_A_ESD_0_H(mprj_analog_io[4]),
    .PAD_A_ESD_1_H(\mprj_pads.area1_io_pad[11]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area1_io_pad[11]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[11]),
    .TIE_HI_ESD(\mprj_pads.area1_io_pad[11]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area1_io_pad[11]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda1),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa1),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[11]),
    .DM({mprj_io_dm[35],
    mprj_io_dm[34],
    mprj_io_dm[33]}));
 sky130_ef_io__com_bus_slice_20um FILLER_549 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_548 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_547 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_546 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area2_io_pad[6]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[25]),
    .ANALOG_POL(mprj_io_analog_pol[25]),
    .ANALOG_SEL(mprj_io_analog_sel[25]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area2_io_pad[6]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[25]),
    .ENABLE_VSWITCH_H(\mprj_pads.area2_io_pad[6]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area2_io_pad[6]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[25]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[25]),
    .IN(mprj_io_in[25]),
    .IN_H(\mprj_pads.area2_io_pad[6]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[25]),
    .OE_N(mprj_io_oeb[25]),
    .OUT(mprj_io_out[25]),
    .PAD(mprj_io[25]),
    .PAD_A_ESD_0_H(mprj_analog_io[18]),
    .PAD_A_ESD_1_H(\mprj_pads.area2_io_pad[6]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area2_io_pad[6]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[25]),
    .TIE_HI_ESD(\mprj_pads.area2_io_pad[6]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area2_io_pad[6]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda2),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa2),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[25]),
    .DM({mprj_io_dm[77],
    mprj_io_dm[76],
    mprj_io_dm[75]}));
 sky130_ef_io__com_bus_slice_10um FILLER_551 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_552 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_553 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_550 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_555 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_760 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_761 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_762 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_763 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area1_io_pad[12]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[12]),
    .ANALOG_POL(mprj_io_analog_pol[12]),
    .ANALOG_SEL(mprj_io_analog_sel[12]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area1_io_pad[12]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[12]),
    .ENABLE_VSWITCH_H(\mprj_pads.area1_io_pad[12]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area1_io_pad[12]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[12]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[12]),
    .IN(mprj_io_in[12]),
    .IN_H(\mprj_pads.area1_io_pad[12]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[12]),
    .OE_N(mprj_io_oeb[12]),
    .OUT(mprj_io_out[12]),
    .PAD(mprj_io[12]),
    .PAD_A_ESD_0_H(mprj_analog_io[5]),
    .PAD_A_ESD_1_H(\mprj_pads.area1_io_pad[12]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area1_io_pad[12]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[12]),
    .TIE_HI_ESD(\mprj_pads.area1_io_pad[12]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area1_io_pad[12]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda1),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa1),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[12]),
    .DM({mprj_io_dm[38],
    mprj_io_dm[37],
    mprj_io_dm[36]}));
 sky130_ef_io__com_bus_slice_20um FILLER_765 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_766 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_767 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_768 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_559 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_558 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_557 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_556 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__vssa_hvc_clamped_pad user2_vssa_hvclamp_pad (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA_PAD(vssa2_pad),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_10um FILLER_561 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_562 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_563 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_560 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_565 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_769 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_770 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_771 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_775 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_776 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_777 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_773 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_772 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__vdda_hvc_clamped_pad \user1_vdda_hvclamp_pad[0]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VDDA_PAD(vdda1_pad),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_569 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_568 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_567 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_566 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__vddio_hvc_clamped_pad \mgmt_vddio_hvclamp_pad[1]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VDDIO_PAD(vddio_pad2),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_10um FILLER_571 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_572 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_573 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_570 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_575 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_778 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_779 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_780 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_781 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_784 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_785 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_782 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area1_io_pad[13]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[13]),
    .ANALOG_POL(mprj_io_analog_pol[13]),
    .ANALOG_SEL(mprj_io_analog_sel[13]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area1_io_pad[13]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[13]),
    .ENABLE_VSWITCH_H(\mprj_pads.area1_io_pad[13]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area1_io_pad[13]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[13]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[13]),
    .IN(mprj_io_in[13]),
    .IN_H(\mprj_pads.area1_io_pad[13]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[13]),
    .OE_N(mprj_io_oeb[13]),
    .OUT(mprj_io_out[13]),
    .PAD(mprj_io[13]),
    .PAD_A_ESD_0_H(mprj_analog_io[6]),
    .PAD_A_ESD_1_H(\mprj_pads.area1_io_pad[13]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area1_io_pad[13]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[13]),
    .TIE_HI_ESD(\mprj_pads.area1_io_pad[13]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area1_io_pad[13]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda1),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa1),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[13]),
    .DM({mprj_io_dm[41],
    mprj_io_dm[40],
    mprj_io_dm[39]}));
 sky130_ef_io__com_bus_slice_20um FILLER_579 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_578 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_577 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_576 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__vccd_lvc_clamped3_pad user2_vccd_lvclamp_pad (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VCCD_PAD(vccd2_pad),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VCCD1(vccd2),
    .VSSD1(vssd2));
 sky130_ef_io__com_bus_slice_10um FILLER_581 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_582 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_583 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_580 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_585 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_790 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_789 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_788 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_787 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_786 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__vccd_lvc_clamped3_pad user1_vccd_lvclamp_pad (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VCCD_PAD(vccd1_pad),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VCCD1(vccd1),
    .VSSD1(vssd1));
 sky130_ef_io__com_bus_slice_5um FILLER_791 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_792 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_795 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_794 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_589 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_588 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_587 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_586 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area2_io_pad[5]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[24]),
    .ANALOG_POL(mprj_io_analog_pol[24]),
    .ANALOG_SEL(mprj_io_analog_sel[24]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area2_io_pad[5]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[24]),
    .ENABLE_VSWITCH_H(\mprj_pads.area2_io_pad[5]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area2_io_pad[5]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[24]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[24]),
    .IN(mprj_io_in[24]),
    .IN_H(\mprj_pads.area2_io_pad[5]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[24]),
    .OE_N(mprj_io_oeb[24]),
    .OUT(mprj_io_out[24]),
    .PAD(mprj_io[24]),
    .PAD_A_ESD_0_H(mprj_analog_io[17]),
    .PAD_A_ESD_1_H(\mprj_pads.area2_io_pad[5]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area2_io_pad[5]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[24]),
    .TIE_HI_ESD(\mprj_pads.area2_io_pad[5]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area2_io_pad[5]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda2),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa2),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[24]),
    .DM({mprj_io_dm[74],
    mprj_io_dm[73],
    mprj_io_dm[72]}));
 sky130_ef_io__com_bus_slice_10um FILLER_591 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_592 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_593 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_590 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_595 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_796 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_797 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_798 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_799 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_800 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_803 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_801 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area1_io_pad[14]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[14]),
    .ANALOG_POL(mprj_io_analog_pol[14]),
    .ANALOG_SEL(mprj_io_analog_sel[14]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area1_io_pad[14]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[14]),
    .ENABLE_VSWITCH_H(\mprj_pads.area1_io_pad[14]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area1_io_pad[14]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[14]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[14]),
    .IN(mprj_io_in[14]),
    .IN_H(\mprj_pads.area1_io_pad[14]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[14]),
    .OE_N(mprj_io_oeb[14]),
    .OUT(mprj_io_out[14]),
    .PAD(mprj_io[14]),
    .PAD_A_ESD_0_H(mprj_analog_io[7]),
    .PAD_A_ESD_1_H(\mprj_pads.area1_io_pad[14]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area1_io_pad[14]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[14]),
    .TIE_HI_ESD(\mprj_pads.area1_io_pad[14]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area1_io_pad[14]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda1),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa1),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[14]),
    .DM({mprj_io_dm[44],
    mprj_io_dm[43],
    mprj_io_dm[42]}));
 sky130_ef_io__com_bus_slice_20um FILLER_600 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_599 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_598 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_597 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_596 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_10um FILLER_601 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_602 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_604 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_603 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__corner_pad user2_corner (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_5 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_9 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_8 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_7 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_6 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_10um FILLER_13 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_12 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_11 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_10 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area2_io_pad[4]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[23]),
    .ANALOG_POL(mprj_io_analog_pol[23]),
    .ANALOG_SEL(mprj_io_analog_sel[23]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area2_io_pad[4]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[23]),
    .ENABLE_VSWITCH_H(\mprj_pads.area2_io_pad[4]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area2_io_pad[4]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[23]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[23]),
    .IN(mprj_io_in[23]),
    .IN_H(\mprj_pads.area2_io_pad[4]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[23]),
    .OE_N(mprj_io_oeb[23]),
    .OUT(mprj_io_out[23]),
    .PAD(mprj_io[23]),
    .PAD_A_ESD_0_H(mprj_analog_io[16]),
    .PAD_A_ESD_1_H(\mprj_pads.area2_io_pad[4]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area2_io_pad[4]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[23]),
    .TIE_HI_ESD(\mprj_pads.area2_io_pad[4]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area2_io_pad[4]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda2),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa2),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[23]),
    .DM({mprj_io_dm[71],
    mprj_io_dm[70],
    mprj_io_dm[69]}));
 sky130_ef_io__com_bus_slice_5um FILLER_14 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_16 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_15 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_18 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_19 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_20 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_21 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_22 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_23 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_24 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_25 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_10um FILLER_26 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_27 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area2_io_pad[3]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[22]),
    .ANALOG_POL(mprj_io_analog_pol[22]),
    .ANALOG_SEL(mprj_io_analog_sel[22]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area2_io_pad[3]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[22]),
    .ENABLE_VSWITCH_H(\mprj_pads.area2_io_pad[3]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area2_io_pad[3]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[22]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[22]),
    .IN(mprj_io_in[22]),
    .IN_H(\mprj_pads.area2_io_pad[3]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[22]),
    .OE_N(mprj_io_oeb[22]),
    .OUT(mprj_io_out[22]),
    .PAD(mprj_io[22]),
    .PAD_A_ESD_0_H(mprj_analog_io[15]),
    .PAD_A_ESD_1_H(\mprj_pads.area2_io_pad[3]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area2_io_pad[3]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[22]),
    .TIE_HI_ESD(\mprj_pads.area2_io_pad[3]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area2_io_pad[3]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda2),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa2),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[22]),
    .DM({mprj_io_dm[68],
    mprj_io_dm[67],
    mprj_io_dm[66]}));
 sky130_ef_io__com_bus_slice_1um FILLER_29 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_28 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_34 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_33 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_32 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_31 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_37 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_36 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_35 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area2_io_pad[2]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[21]),
    .ANALOG_POL(mprj_io_analog_pol[21]),
    .ANALOG_SEL(mprj_io_analog_sel[21]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area2_io_pad[2]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[21]),
    .ENABLE_VSWITCH_H(\mprj_pads.area2_io_pad[2]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area2_io_pad[2]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[21]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[21]),
    .IN(mprj_io_in[21]),
    .IN_H(\mprj_pads.area2_io_pad[2]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[21]),
    .OE_N(mprj_io_oeb[21]),
    .OUT(mprj_io_out[21]),
    .PAD(mprj_io[21]),
    .PAD_A_ESD_0_H(mprj_analog_io[14]),
    .PAD_A_ESD_1_H(\mprj_pads.area2_io_pad[2]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area2_io_pad[2]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[21]),
    .TIE_HI_ESD(\mprj_pads.area2_io_pad[2]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area2_io_pad[2]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda2),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa2),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[21]),
    .DM({mprj_io_dm[65],
    mprj_io_dm[64],
    mprj_io_dm[63]}));
 sky130_ef_io__com_bus_slice_10um FILLER_39 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_40 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_42 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_41 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_38 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_45 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_44 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_47 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_46 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_10um FILLER_52 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_51 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_50 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_49 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_48 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area2_io_pad[1]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[20]),
    .ANALOG_POL(mprj_io_analog_pol[20]),
    .ANALOG_SEL(mprj_io_analog_sel[20]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area2_io_pad[1]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[20]),
    .ENABLE_VSWITCH_H(\mprj_pads.area2_io_pad[1]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area2_io_pad[1]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[20]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[20]),
    .IN(mprj_io_in[20]),
    .IN_H(\mprj_pads.area2_io_pad[1]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[20]),
    .OE_N(mprj_io_oeb[20]),
    .OUT(mprj_io_out[20]),
    .PAD(mprj_io[20]),
    .PAD_A_ESD_0_H(mprj_analog_io[13]),
    .PAD_A_ESD_1_H(\mprj_pads.area2_io_pad[1]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area2_io_pad[1]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[20]),
    .TIE_HI_ESD(\mprj_pads.area2_io_pad[1]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area2_io_pad[1]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda2),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa2),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[20]),
    .DM({mprj_io_dm[62],
    mprj_io_dm[61],
    mprj_io_dm[60]}));
 sky130_ef_io__com_bus_slice_5um FILLER_53 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_55 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_54 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_58 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_57 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_62 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_61 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_60 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_59 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area2_io_pad[0]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[19]),
    .ANALOG_POL(mprj_io_analog_pol[19]),
    .ANALOG_SEL(mprj_io_analog_sel[19]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area2_io_pad[0]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[19]),
    .ENABLE_VSWITCH_H(\mprj_pads.area2_io_pad[0]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area2_io_pad[0]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[19]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[19]),
    .IN(mprj_io_in[19]),
    .IN_H(\mprj_pads.area2_io_pad[0]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[19]),
    .OE_N(mprj_io_oeb[19]),
    .OUT(mprj_io_out[19]),
    .PAD(mprj_io[19]),
    .PAD_A_ESD_0_H(mprj_analog_io[12]),
    .PAD_A_ESD_1_H(\mprj_pads.area2_io_pad[0]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area2_io_pad[0]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[19]),
    .TIE_HI_ESD(\mprj_pads.area2_io_pad[0]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area2_io_pad[0]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda2),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa2),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[19]),
    .DM({mprj_io_dm[59],
    mprj_io_dm[58],
    mprj_io_dm[57]}));
 sky130_ef_io__com_bus_slice_10um FILLER_65 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_66 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_69 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_68 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_67 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_64 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_63 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_74 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_73 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_72 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_71 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_77 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_76 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_75 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__vssio_hvc_clamped_pad \mgmt_vssio_hvclamp_pad[1]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSIO_PAD(vssio_pad2),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_10um FILLER_79 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_80 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_82 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_81 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_78 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa2),
    .VDDA(vdda2),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__disconnect_vdda_slice_5um disconnect_vdda_0 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_SB3 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_87 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_86 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_88 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_89 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_90 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_91 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_92 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_93 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area1_io_pad[18]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[18]),
    .ANALOG_POL(mprj_io_analog_pol[18]),
    .ANALOG_SEL(mprj_io_analog_sel[18]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area1_io_pad[18]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[18]),
    .ENABLE_VSWITCH_H(\mprj_pads.area1_io_pad[18]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area1_io_pad[18]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[18]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[18]),
    .IN(mprj_io_in[18]),
    .IN_H(\mprj_pads.area1_io_pad[18]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[18]),
    .OE_N(mprj_io_oeb[18]),
    .OUT(mprj_io_out[18]),
    .PAD(mprj_io[18]),
    .PAD_A_ESD_0_H(mprj_analog_io[11]),
    .PAD_A_ESD_1_H(\mprj_pads.area1_io_pad[18]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area1_io_pad[18]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[18]),
    .TIE_HI_ESD(\mprj_pads.area1_io_pad[18]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area1_io_pad[18]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda1),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa1),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[18]),
    .DM({mprj_io_dm[56],
    mprj_io_dm[55],
    mprj_io_dm[54]}));
 sky130_ef_io__com_bus_slice_5um FILLER_94 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_96 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_95 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_101 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_100 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_99 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_98 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_103 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_102 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_104 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_105 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_106 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_107 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_108 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_109 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_110 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_111 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_112 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_113 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_114 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_115 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_118 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_119 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_120 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_121 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_122 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_116 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area1_io_pad[17]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[17]),
    .ANALOG_POL(mprj_io_analog_pol[17]),
    .ANALOG_SEL(mprj_io_analog_sel[17]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area1_io_pad[17]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[17]),
    .ENABLE_VSWITCH_H(\mprj_pads.area1_io_pad[17]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area1_io_pad[17]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[17]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[17]),
    .IN(mprj_io_in[17]),
    .IN_H(\mprj_pads.area1_io_pad[17]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[17]),
    .OE_N(mprj_io_oeb[17]),
    .OUT(mprj_io_out[17]),
    .PAD(mprj_io[17]),
    .PAD_A_ESD_0_H(mprj_analog_io[10]),
    .PAD_A_ESD_1_H(\mprj_pads.area1_io_pad[17]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area1_io_pad[17]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[17]),
    .TIE_HI_ESD(\mprj_pads.area1_io_pad[17]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area1_io_pad[17]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda1),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa1),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[17]),
    .DM({mprj_io_dm[53],
    mprj_io_dm[52],
    mprj_io_dm[51]}));
 sky130_ef_io__com_bus_slice_10um FILLER_126 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_125 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_124 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_123 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area1_io_pad[16]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[16]),
    .ANALOG_POL(mprj_io_analog_pol[16]),
    .ANALOG_SEL(mprj_io_analog_sel[16]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area1_io_pad[16]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[16]),
    .ENABLE_VSWITCH_H(\mprj_pads.area1_io_pad[16]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area1_io_pad[16]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[16]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[16]),
    .IN(mprj_io_in[16]),
    .IN_H(\mprj_pads.area1_io_pad[16]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[16]),
    .OE_N(mprj_io_oeb[16]),
    .OUT(mprj_io_out[16]),
    .PAD(mprj_io[16]),
    .PAD_A_ESD_0_H(mprj_analog_io[9]),
    .PAD_A_ESD_1_H(\mprj_pads.area1_io_pad[16]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area1_io_pad[16]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[16]),
    .TIE_HI_ESD(\mprj_pads.area1_io_pad[16]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area1_io_pad[16]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda1),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa1),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[16]),
    .DM({mprj_io_dm[50],
    mprj_io_dm[49],
    mprj_io_dm[48]}));
 sky130_ef_io__com_bus_slice_5um FILLER_127 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_129 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_128 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_133 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_132 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_131 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_136 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_135 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_134 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__vssa_hvc_clamped_pad \user1_vssa_hvclamp_pad[0]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA_PAD(vssa1_pad),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_10um FILLER_139 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_140 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_142 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_141 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_138 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_137 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_144 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_148 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_147 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_146 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_145 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_10um FILLER_152 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_151 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_150 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_149 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__gpiov2_pad_wrapped \mprj_pads.area1_io_pad[15]  (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .ANALOG_EN(mprj_io_analog_en[15]),
    .ANALOG_POL(mprj_io_analog_pol[15]),
    .ANALOG_SEL(mprj_io_analog_sel[15]),
    .ENABLE_H(porb_h),
    .ENABLE_INP_H(\mprj_pads.area1_io_pad[15]__TIE_LO_ESD ),
    .ENABLE_VDDA_H(porb_h),
    .ENABLE_VDDIO(mprj_io_one[15]),
    .ENABLE_VSWITCH_H(\mprj_pads.area1_io_pad[15]__TIE_LO_ESD ),
    .HLD_H_N(\mprj_pads.area1_io_pad[15]__HLD_H_N ),
    .HLD_OVR(mprj_io_holdover[15]),
    .IB_MODE_SEL(mprj_io_ib_mode_sel[15]),
    .IN(mprj_io_in[15]),
    .IN_H(\mprj_pads.area1_io_pad[15]__IN_H ),
    .INP_DIS(mprj_io_inp_dis[15]),
    .OE_N(mprj_io_oeb[15]),
    .OUT(mprj_io_out[15]),
    .PAD(mprj_io[15]),
    .PAD_A_ESD_0_H(mprj_analog_io[8]),
    .PAD_A_ESD_1_H(\mprj_pads.area1_io_pad[15]__PAD_A_ESD_1_H ),
    .PAD_A_NOESD_H(\mprj_pads.area1_io_pad[15]__PAD_A_NOESD_H ),
    .SLOW(mprj_io_slow_sel[15]),
    .TIE_HI_ESD(\mprj_pads.area1_io_pad[15]__HLD_H_N ),
    .TIE_LO_ESD(\mprj_pads.area1_io_pad[15]__TIE_LO_ESD ),
    .VCCD(vccd),
    .VCCHIB(vccd),
    .VDDA(vdda1),
    .VDDIO(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VSSA(vssa1),
    .VSSD(vssd),
    .VSSIO(vssio),
    .VSSIO_Q(gpio_pad__VSSIO_Q),
    .VSWITCH(vddio),
    .VTRIP_SEL(mprj_io_vtrip_sel[15]),
    .DM({mprj_io_dm[47],
    mprj_io_dm[46],
    mprj_io_dm[45]}));
 sky130_ef_io__com_bus_slice_5um FILLER_153 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_155 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_154 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_157 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_158 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_159 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_160 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_161 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_162 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_163 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_164 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_10um FILLER_165 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_808 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_807 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_806 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_805 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_804 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_810 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_811 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_20um FILLER_809 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_5um FILLER_166 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_169 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_168 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__com_bus_slice_1um FILLER_167 (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
 sky130_ef_io__corner_pad user1_corner (.AMUXBUS_A(gpio_pad__AMUXBUS_A),
    .AMUXBUS_B(gpio_pad__AMUXBUS_B),
    .VSSA(vssa1),
    .VDDA(vdda1),
    .VSWITCH(vddio),
    .VDDIO_Q(gpio_pad__VDDIO_Q),
    .VCCHIB(vccd),
    .VDDIO(vddio),
    .VCCD(vccd),
    .VSSIO(vssio),
    .VSSD(vssd),
    .VSSIO_Q(gpio_pad__VSSIO_Q));
endmodule
