*----------------------------------------------------------
* sky130_ef_io__gpiov2_pad
* Wrapper around SkyWater gpiov2 pad
*----------------------------------------------------------

.SUBCKT sky130_ef_io__gpiov2_pad
+ IN_H PAD_A_NOESD_H PAD_A_ESD_0_H PAD_A_ESD_1_H
+ PAD DM[2] DM[1] DM[0] HLD_H_N IN INP_DIS IB_MODE_SEL ENABLE_H ENABLE_VDDA_H
+ ENABLE_INP_H OE_N TIE_HI_ESD TIE_LO_ESD SLOW VTRIP_SEL HLD_OVR
+ ANALOG_EN ANALOG_SEL ENABLE_VDDIO ENABLE_VSWITCH_H ANALOG_POL OUT
+ AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD
+ VSSIO VSSD VSSIO_Q

* Instantiate original version with metal4-only power bus
Xgpiov2_base
+ AMUXBUS_A AMUXBUS_B ANALOG_EN ANALOG_POL ANALOG_SEL
+ DM[2] DM[1] DM[0]
+ ENABLE_H ENABLE_INP_H ENABLE_VDDA_H ENABLE_VDDIO ENABLE_VSWITCH_H
+ HLD_H_N HLD_OVR IB_MODE_SEL
+ IN IN_H INP_DIS OE_N OUT
+ PAD PAD_A_ESD_0_H PAD_A_ESD_1_H PAD_A_NOESD_H
+ SLOW TIE_HI_ESD TIE_LO_ESD
+ VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH
+ VTRIP_SEL
+ sky130_fd_io__top_gpiov2

.ENDS

*----------------------------------------------------------
* sky130_ef_io__gpiov2_pad_wrapped
* Wrapper around sky130_ef_io__gpiov2_pad that forces
* the core-facing pins on tracks
*----------------------------------------------------------

.SUBCKT sky130_ef_io__gpiov2_pad_wrapped
+ IN_H PAD_A_NOESD_H PAD_A_ESD_0_H PAD_A_ESD_1_H
+ PAD DM[2] DM[1] DM[0] HLD_H_N IN INP_DIS IB_MODE_SEL ENABLE_H ENABLE_VDDA_H
+ ENABLE_INP_H OE_N TIE_HI_ESD TIE_LO_ESD SLOW VTRIP_SEL HLD_OVR
+ ANALOG_EN ANALOG_SEL ENABLE_VDDIO ENABLE_VSWITCH_H ANALOG_POL OUT
+ AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD
+ VSSIO VSSD VSSIO_Q

Xgpiov2_ef
+ IN_H PAD_A_NOESD_H PAD_A_ESD_0_H PAD_A_ESD_1_H
+ PAD DM[2] DM[1] DM[0] HLD_H_N IN INP_DIS IB_MODE_SEL ENABLE_H ENABLE_VDDA_H
+ ENABLE_INP_H OE_N TIE_HI_ESD TIE_LO_ESD SLOW VTRIP_SEL HLD_OVR
+ ANALOG_EN ANALOG_SEL ENABLE_VDDIO ENABLE_VSWITCH_H ANALOG_POL OUT
+ AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD
+ VSSIO VSSD VSSIO_Q sky130_ef_io__gpiov2_pad

.ENDS

