magic
tech sky130A
magscale 1 2
timestamp 1665595734
<< viali >>
rect 3617 4641 3651 4675
rect 6469 4641 6503 4675
rect 3249 4573 3283 4607
rect 6837 4573 6871 4607
rect 2329 4097 2363 4131
rect 3617 4097 3651 4131
rect 5089 4097 5123 4131
rect 5825 4097 5859 4131
rect 1961 4029 1995 4063
rect 3341 4029 3375 4063
rect 4629 4029 4663 4063
rect 6193 4029 6227 4063
rect 1869 3553 1903 3587
rect 3801 3553 3835 3587
rect 5273 3553 5307 3587
rect 1593 3485 1627 3519
rect 3617 3485 3651 3519
rect 4905 3485 4939 3519
rect 1133 3009 1167 3043
rect 4353 3009 4387 3043
rect 6837 3009 6871 3043
rect 1501 2941 1535 2975
rect 4537 2941 4571 2975
rect 6469 2941 6503 2975
rect 1501 2465 1535 2499
rect 6285 2465 6319 2499
rect 1133 2397 1167 2431
rect 6561 2397 6595 2431
rect 765 1921 799 1955
rect 2237 1921 2271 1955
rect 5273 1921 5307 1955
rect 5825 1921 5859 1955
rect 949 1853 983 1887
rect 2513 1853 2547 1887
rect 4905 1853 4939 1887
rect 6193 1853 6227 1887
rect 1501 1309 1535 1343
rect 2145 1309 2179 1343
rect 6745 1309 6779 1343
rect 6009 1241 6043 1275
<< metal1 >>
rect 368 4922 7544 4944
rect 368 4870 1110 4922
rect 1162 4870 1174 4922
rect 1226 4870 1238 4922
rect 1290 4870 1302 4922
rect 1354 4870 1366 4922
rect 1418 4870 2903 4922
rect 2955 4870 2967 4922
rect 3019 4870 3031 4922
rect 3083 4870 3095 4922
rect 3147 4870 3159 4922
rect 3211 4870 4696 4922
rect 4748 4870 4760 4922
rect 4812 4870 4824 4922
rect 4876 4870 4888 4922
rect 4940 4870 4952 4922
rect 5004 4870 6489 4922
rect 6541 4870 6553 4922
rect 6605 4870 6617 4922
rect 6669 4870 6681 4922
rect 6733 4870 6745 4922
rect 6797 4870 7544 4922
rect 368 4848 7544 4870
rect 3234 4700 3240 4752
rect 3292 4740 3298 4752
rect 3292 4712 3648 4740
rect 3292 4700 3298 4712
rect 3620 4681 3648 4712
rect 3605 4675 3663 4681
rect 3605 4641 3617 4675
rect 3651 4641 3663 4675
rect 3605 4635 3663 4641
rect 6457 4675 6515 4681
rect 6457 4641 6469 4675
rect 6503 4672 6515 4675
rect 7466 4672 7472 4684
rect 6503 4644 7472 4672
rect 6503 4641 6515 4644
rect 6457 4635 6515 4641
rect 7466 4632 7472 4644
rect 7524 4632 7530 4684
rect 3234 4604 3240 4616
rect 3195 4576 3240 4604
rect 3234 4564 3240 4576
rect 3292 4564 3298 4616
rect 6825 4607 6883 4613
rect 6825 4573 6837 4607
rect 6871 4604 6883 4607
rect 7282 4604 7288 4616
rect 6871 4576 7288 4604
rect 6871 4573 6883 4576
rect 6825 4567 6883 4573
rect 7282 4564 7288 4576
rect 7340 4564 7346 4616
rect 368 4378 7699 4400
rect 368 4326 2006 4378
rect 2058 4326 2070 4378
rect 2122 4326 2134 4378
rect 2186 4326 2198 4378
rect 2250 4326 2262 4378
rect 2314 4326 3799 4378
rect 3851 4326 3863 4378
rect 3915 4326 3927 4378
rect 3979 4326 3991 4378
rect 4043 4326 4055 4378
rect 4107 4326 5592 4378
rect 5644 4326 5656 4378
rect 5708 4326 5720 4378
rect 5772 4326 5784 4378
rect 5836 4326 5848 4378
rect 5900 4326 7385 4378
rect 7437 4326 7449 4378
rect 7501 4326 7513 4378
rect 7565 4326 7577 4378
rect 7629 4326 7641 4378
rect 7693 4326 7699 4378
rect 368 4304 7699 4326
rect 2317 4131 2375 4137
rect 2317 4097 2329 4131
rect 2363 4128 2375 4131
rect 2682 4128 2688 4140
rect 2363 4100 2688 4128
rect 2363 4097 2375 4100
rect 2317 4091 2375 4097
rect 2682 4088 2688 4100
rect 2740 4088 2746 4140
rect 3418 4088 3424 4140
rect 3476 4128 3482 4140
rect 3605 4131 3663 4137
rect 3605 4128 3617 4131
rect 3476 4100 3617 4128
rect 3476 4088 3482 4100
rect 3605 4097 3617 4100
rect 3651 4097 3663 4131
rect 5074 4128 5080 4140
rect 5035 4100 5080 4128
rect 3605 4091 3663 4097
rect 5074 4088 5080 4100
rect 5132 4088 5138 4140
rect 5258 4088 5264 4140
rect 5316 4128 5322 4140
rect 5813 4131 5871 4137
rect 5813 4128 5825 4131
rect 5316 4100 5825 4128
rect 5316 4088 5322 4100
rect 5813 4097 5825 4100
rect 5859 4097 5871 4131
rect 5813 4091 5871 4097
rect 1949 4063 2007 4069
rect 1949 4029 1961 4063
rect 1995 4060 2007 4063
rect 2590 4060 2596 4072
rect 1995 4032 2596 4060
rect 1995 4029 2007 4032
rect 1949 4023 2007 4029
rect 2590 4020 2596 4032
rect 2648 4020 2654 4072
rect 3326 4060 3332 4072
rect 3287 4032 3332 4060
rect 3326 4020 3332 4032
rect 3384 4020 3390 4072
rect 4614 4060 4620 4072
rect 4575 4032 4620 4060
rect 4614 4020 4620 4032
rect 4672 4020 4678 4072
rect 5534 4020 5540 4072
rect 5592 4060 5598 4072
rect 6181 4063 6239 4069
rect 6181 4060 6193 4063
rect 5592 4032 6193 4060
rect 5592 4020 5598 4032
rect 6181 4029 6193 4032
rect 6227 4029 6239 4063
rect 6181 4023 6239 4029
rect 368 3834 7544 3856
rect 368 3782 1110 3834
rect 1162 3782 1174 3834
rect 1226 3782 1238 3834
rect 1290 3782 1302 3834
rect 1354 3782 1366 3834
rect 1418 3782 2903 3834
rect 2955 3782 2967 3834
rect 3019 3782 3031 3834
rect 3083 3782 3095 3834
rect 3147 3782 3159 3834
rect 3211 3782 4696 3834
rect 4748 3782 4760 3834
rect 4812 3782 4824 3834
rect 4876 3782 4888 3834
rect 4940 3782 4952 3834
rect 5004 3782 6489 3834
rect 6541 3782 6553 3834
rect 6605 3782 6617 3834
rect 6669 3782 6681 3834
rect 6733 3782 6745 3834
rect 6797 3782 7544 3834
rect 368 3760 7544 3782
rect 3694 3612 3700 3664
rect 3752 3652 3758 3664
rect 3752 3624 3832 3652
rect 3752 3612 3758 3624
rect 1854 3584 1860 3596
rect 1815 3556 1860 3584
rect 1854 3544 1860 3556
rect 1912 3544 1918 3596
rect 3804 3593 3832 3624
rect 4154 3612 4160 3664
rect 4212 3652 4218 3664
rect 4212 3624 5304 3652
rect 4212 3612 4218 3624
rect 5276 3593 5304 3624
rect 3789 3587 3847 3593
rect 3789 3553 3801 3587
rect 3835 3553 3847 3587
rect 3789 3547 3847 3553
rect 5261 3587 5319 3593
rect 5261 3553 5273 3587
rect 5307 3553 5319 3587
rect 5261 3547 5319 3553
rect 1581 3519 1639 3525
rect 1581 3485 1593 3519
rect 1627 3485 1639 3519
rect 1581 3479 1639 3485
rect 3605 3519 3663 3525
rect 3605 3485 3617 3519
rect 3651 3516 3663 3519
rect 3694 3516 3700 3528
rect 3651 3488 3700 3516
rect 3651 3485 3663 3488
rect 3605 3479 3663 3485
rect 1596 3448 1624 3479
rect 3694 3476 3700 3488
rect 3752 3476 3758 3528
rect 4154 3476 4160 3528
rect 4212 3516 4218 3528
rect 4893 3519 4951 3525
rect 4893 3516 4905 3519
rect 4212 3488 4905 3516
rect 4212 3476 4218 3488
rect 4893 3485 4905 3488
rect 4939 3485 4951 3519
rect 4893 3479 4951 3485
rect 1854 3448 1860 3460
rect 1596 3420 1860 3448
rect 1854 3408 1860 3420
rect 1912 3408 1918 3460
rect 368 3290 7699 3312
rect 368 3238 2006 3290
rect 2058 3238 2070 3290
rect 2122 3238 2134 3290
rect 2186 3238 2198 3290
rect 2250 3238 2262 3290
rect 2314 3238 3799 3290
rect 3851 3238 3863 3290
rect 3915 3238 3927 3290
rect 3979 3238 3991 3290
rect 4043 3238 4055 3290
rect 4107 3238 5592 3290
rect 5644 3238 5656 3290
rect 5708 3238 5720 3290
rect 5772 3238 5784 3290
rect 5836 3238 5848 3290
rect 5900 3238 7385 3290
rect 7437 3238 7449 3290
rect 7501 3238 7513 3290
rect 7565 3238 7577 3290
rect 7629 3238 7641 3290
rect 7693 3238 7699 3290
rect 368 3216 7699 3238
rect 1026 3000 1032 3052
rect 1084 3040 1090 3052
rect 1121 3043 1179 3049
rect 1121 3040 1133 3043
rect 1084 3012 1133 3040
rect 1084 3000 1090 3012
rect 1121 3009 1133 3012
rect 1167 3009 1179 3043
rect 1121 3003 1179 3009
rect 4341 3043 4399 3049
rect 4341 3009 4353 3043
rect 4387 3040 4399 3043
rect 4430 3040 4436 3052
rect 4387 3012 4436 3040
rect 4387 3009 4399 3012
rect 4341 3003 4399 3009
rect 4430 3000 4436 3012
rect 4488 3000 4494 3052
rect 6825 3043 6883 3049
rect 6825 3009 6837 3043
rect 6871 3040 6883 3043
rect 7098 3040 7104 3052
rect 6871 3012 7104 3040
rect 6871 3009 6883 3012
rect 6825 3003 6883 3009
rect 7098 3000 7104 3012
rect 7156 3000 7162 3052
rect 1394 2932 1400 2984
rect 1452 2972 1458 2984
rect 1489 2975 1547 2981
rect 1489 2972 1501 2975
rect 1452 2944 1501 2972
rect 1452 2932 1458 2944
rect 1489 2941 1501 2944
rect 1535 2941 1547 2975
rect 4522 2972 4528 2984
rect 4483 2944 4528 2972
rect 1489 2935 1547 2941
rect 4522 2932 4528 2944
rect 4580 2932 4586 2984
rect 6457 2975 6515 2981
rect 6457 2941 6469 2975
rect 6503 2972 6515 2975
rect 7006 2972 7012 2984
rect 6503 2944 7012 2972
rect 6503 2941 6515 2944
rect 6457 2935 6515 2941
rect 7006 2932 7012 2944
rect 7064 2932 7070 2984
rect 368 2746 7544 2768
rect 368 2694 1110 2746
rect 1162 2694 1174 2746
rect 1226 2694 1238 2746
rect 1290 2694 1302 2746
rect 1354 2694 1366 2746
rect 1418 2694 2903 2746
rect 2955 2694 2967 2746
rect 3019 2694 3031 2746
rect 3083 2694 3095 2746
rect 3147 2694 3159 2746
rect 3211 2694 4696 2746
rect 4748 2694 4760 2746
rect 4812 2694 4824 2746
rect 4876 2694 4888 2746
rect 4940 2694 4952 2746
rect 5004 2694 6489 2746
rect 6541 2694 6553 2746
rect 6605 2694 6617 2746
rect 6669 2694 6681 2746
rect 6733 2694 6745 2746
rect 6797 2694 7544 2746
rect 368 2672 7544 2694
rect 474 2524 480 2576
rect 532 2564 538 2576
rect 6362 2564 6368 2576
rect 532 2536 1532 2564
rect 532 2524 538 2536
rect 1504 2505 1532 2536
rect 6288 2536 6368 2564
rect 6288 2505 6316 2536
rect 6362 2524 6368 2536
rect 6420 2524 6426 2576
rect 1489 2499 1547 2505
rect 1489 2465 1501 2499
rect 1535 2465 1547 2499
rect 1489 2459 1547 2465
rect 6273 2499 6331 2505
rect 6273 2465 6285 2499
rect 6319 2465 6331 2499
rect 6273 2459 6331 2465
rect 474 2388 480 2440
rect 532 2428 538 2440
rect 1121 2431 1179 2437
rect 1121 2428 1133 2431
rect 532 2400 1133 2428
rect 532 2388 538 2400
rect 1121 2397 1133 2400
rect 1167 2397 1179 2431
rect 1121 2391 1179 2397
rect 6362 2388 6368 2440
rect 6420 2428 6426 2440
rect 6549 2431 6607 2437
rect 6549 2428 6561 2431
rect 6420 2400 6561 2428
rect 6420 2388 6426 2400
rect 6549 2397 6561 2400
rect 6595 2397 6607 2431
rect 6549 2391 6607 2397
rect 368 2202 7699 2224
rect 368 2150 2006 2202
rect 2058 2150 2070 2202
rect 2122 2150 2134 2202
rect 2186 2150 2198 2202
rect 2250 2150 2262 2202
rect 2314 2150 3799 2202
rect 3851 2150 3863 2202
rect 3915 2150 3927 2202
rect 3979 2150 3991 2202
rect 4043 2150 4055 2202
rect 4107 2150 5592 2202
rect 5644 2150 5656 2202
rect 5708 2150 5720 2202
rect 5772 2150 5784 2202
rect 5836 2150 5848 2202
rect 5900 2150 7385 2202
rect 7437 2150 7449 2202
rect 7501 2150 7513 2202
rect 7565 2150 7577 2202
rect 7629 2150 7641 2202
rect 7693 2150 7699 2202
rect 368 2128 7699 2150
rect 753 1955 811 1961
rect 753 1921 765 1955
rect 799 1952 811 1955
rect 842 1952 848 1964
rect 799 1924 848 1952
rect 799 1921 811 1924
rect 753 1915 811 1921
rect 842 1912 848 1924
rect 900 1912 906 1964
rect 2225 1955 2283 1961
rect 2225 1921 2237 1955
rect 2271 1952 2283 1955
rect 2406 1952 2412 1964
rect 2271 1924 2412 1952
rect 2271 1921 2283 1924
rect 2225 1915 2283 1921
rect 2406 1912 2412 1924
rect 2464 1912 2470 1964
rect 5261 1955 5319 1961
rect 5261 1921 5273 1955
rect 5307 1921 5319 1955
rect 5261 1915 5319 1921
rect 934 1884 940 1896
rect 895 1856 940 1884
rect 934 1844 940 1856
rect 992 1844 998 1896
rect 2498 1884 2504 1896
rect 2459 1856 2504 1884
rect 2498 1844 2504 1856
rect 2556 1844 2562 1896
rect 4893 1887 4951 1893
rect 4893 1853 4905 1887
rect 4939 1853 4951 1887
rect 5276 1884 5304 1915
rect 5534 1912 5540 1964
rect 5592 1952 5598 1964
rect 5813 1955 5871 1961
rect 5813 1952 5825 1955
rect 5592 1924 5825 1952
rect 5592 1912 5598 1924
rect 5813 1921 5825 1924
rect 5859 1921 5871 1955
rect 5813 1915 5871 1921
rect 6086 1884 6092 1896
rect 5276 1856 6092 1884
rect 4893 1847 4951 1853
rect 4908 1816 4936 1847
rect 6086 1844 6092 1856
rect 6144 1844 6150 1896
rect 6178 1844 6184 1896
rect 6236 1884 6242 1896
rect 6236 1856 6281 1884
rect 6236 1844 6242 1856
rect 6270 1816 6276 1828
rect 4908 1788 6276 1816
rect 6270 1776 6276 1788
rect 6328 1776 6334 1828
rect 368 1658 7544 1680
rect 368 1606 1110 1658
rect 1162 1606 1174 1658
rect 1226 1606 1238 1658
rect 1290 1606 1302 1658
rect 1354 1606 1366 1658
rect 1418 1606 2903 1658
rect 2955 1606 2967 1658
rect 3019 1606 3031 1658
rect 3083 1606 3095 1658
rect 3147 1606 3159 1658
rect 3211 1606 4696 1658
rect 4748 1606 4760 1658
rect 4812 1606 4824 1658
rect 4876 1606 4888 1658
rect 4940 1606 4952 1658
rect 5004 1606 6489 1658
rect 6541 1606 6553 1658
rect 6605 1606 6617 1658
rect 6669 1606 6681 1658
rect 6733 1606 6745 1658
rect 6797 1606 7544 1658
rect 368 1584 7544 1606
rect 1489 1343 1547 1349
rect 1489 1309 1501 1343
rect 1535 1340 1547 1343
rect 1578 1340 1584 1352
rect 1535 1312 1584 1340
rect 1535 1309 1547 1312
rect 1489 1303 1547 1309
rect 1578 1300 1584 1312
rect 1636 1300 1642 1352
rect 1670 1300 1676 1352
rect 1728 1340 1734 1352
rect 2133 1343 2191 1349
rect 2133 1340 2145 1343
rect 1728 1312 2145 1340
rect 1728 1300 1734 1312
rect 2133 1309 2145 1312
rect 2179 1309 2191 1343
rect 6730 1340 6736 1352
rect 6691 1312 6736 1340
rect 2133 1303 2191 1309
rect 6730 1300 6736 1312
rect 6788 1300 6794 1352
rect 5997 1275 6055 1281
rect 5997 1241 6009 1275
rect 6043 1272 6055 1275
rect 6822 1272 6828 1284
rect 6043 1244 6828 1272
rect 6043 1241 6055 1244
rect 5997 1235 6055 1241
rect 6822 1232 6828 1244
rect 6880 1232 6886 1284
rect 368 1114 7699 1136
rect 368 1062 2006 1114
rect 2058 1062 2070 1114
rect 2122 1062 2134 1114
rect 2186 1062 2198 1114
rect 2250 1062 2262 1114
rect 2314 1062 3799 1114
rect 3851 1062 3863 1114
rect 3915 1062 3927 1114
rect 3979 1062 3991 1114
rect 4043 1062 4055 1114
rect 4107 1062 5592 1114
rect 5644 1062 5656 1114
rect 5708 1062 5720 1114
rect 5772 1062 5784 1114
rect 5836 1062 5848 1114
rect 5900 1062 7385 1114
rect 7437 1062 7449 1114
rect 7501 1062 7513 1114
rect 7565 1062 7577 1114
rect 7629 1062 7641 1114
rect 7693 1062 7699 1114
rect 368 1040 7699 1062
<< via1 >>
rect 1110 4870 1162 4922
rect 1174 4870 1226 4922
rect 1238 4870 1290 4922
rect 1302 4870 1354 4922
rect 1366 4870 1418 4922
rect 2903 4870 2955 4922
rect 2967 4870 3019 4922
rect 3031 4870 3083 4922
rect 3095 4870 3147 4922
rect 3159 4870 3211 4922
rect 4696 4870 4748 4922
rect 4760 4870 4812 4922
rect 4824 4870 4876 4922
rect 4888 4870 4940 4922
rect 4952 4870 5004 4922
rect 6489 4870 6541 4922
rect 6553 4870 6605 4922
rect 6617 4870 6669 4922
rect 6681 4870 6733 4922
rect 6745 4870 6797 4922
rect 3240 4700 3292 4752
rect 7472 4632 7524 4684
rect 3240 4607 3292 4616
rect 3240 4573 3249 4607
rect 3249 4573 3283 4607
rect 3283 4573 3292 4607
rect 3240 4564 3292 4573
rect 7288 4564 7340 4616
rect 2006 4326 2058 4378
rect 2070 4326 2122 4378
rect 2134 4326 2186 4378
rect 2198 4326 2250 4378
rect 2262 4326 2314 4378
rect 3799 4326 3851 4378
rect 3863 4326 3915 4378
rect 3927 4326 3979 4378
rect 3991 4326 4043 4378
rect 4055 4326 4107 4378
rect 5592 4326 5644 4378
rect 5656 4326 5708 4378
rect 5720 4326 5772 4378
rect 5784 4326 5836 4378
rect 5848 4326 5900 4378
rect 7385 4326 7437 4378
rect 7449 4326 7501 4378
rect 7513 4326 7565 4378
rect 7577 4326 7629 4378
rect 7641 4326 7693 4378
rect 2688 4088 2740 4140
rect 3424 4088 3476 4140
rect 5080 4131 5132 4140
rect 5080 4097 5089 4131
rect 5089 4097 5123 4131
rect 5123 4097 5132 4131
rect 5080 4088 5132 4097
rect 5264 4088 5316 4140
rect 2596 4020 2648 4072
rect 3332 4063 3384 4072
rect 3332 4029 3341 4063
rect 3341 4029 3375 4063
rect 3375 4029 3384 4063
rect 3332 4020 3384 4029
rect 4620 4063 4672 4072
rect 4620 4029 4629 4063
rect 4629 4029 4663 4063
rect 4663 4029 4672 4063
rect 4620 4020 4672 4029
rect 5540 4020 5592 4072
rect 1110 3782 1162 3834
rect 1174 3782 1226 3834
rect 1238 3782 1290 3834
rect 1302 3782 1354 3834
rect 1366 3782 1418 3834
rect 2903 3782 2955 3834
rect 2967 3782 3019 3834
rect 3031 3782 3083 3834
rect 3095 3782 3147 3834
rect 3159 3782 3211 3834
rect 4696 3782 4748 3834
rect 4760 3782 4812 3834
rect 4824 3782 4876 3834
rect 4888 3782 4940 3834
rect 4952 3782 5004 3834
rect 6489 3782 6541 3834
rect 6553 3782 6605 3834
rect 6617 3782 6669 3834
rect 6681 3782 6733 3834
rect 6745 3782 6797 3834
rect 3700 3612 3752 3664
rect 1860 3587 1912 3596
rect 1860 3553 1869 3587
rect 1869 3553 1903 3587
rect 1903 3553 1912 3587
rect 1860 3544 1912 3553
rect 4160 3612 4212 3664
rect 3700 3476 3752 3528
rect 4160 3476 4212 3528
rect 1860 3408 1912 3460
rect 2006 3238 2058 3290
rect 2070 3238 2122 3290
rect 2134 3238 2186 3290
rect 2198 3238 2250 3290
rect 2262 3238 2314 3290
rect 3799 3238 3851 3290
rect 3863 3238 3915 3290
rect 3927 3238 3979 3290
rect 3991 3238 4043 3290
rect 4055 3238 4107 3290
rect 5592 3238 5644 3290
rect 5656 3238 5708 3290
rect 5720 3238 5772 3290
rect 5784 3238 5836 3290
rect 5848 3238 5900 3290
rect 7385 3238 7437 3290
rect 7449 3238 7501 3290
rect 7513 3238 7565 3290
rect 7577 3238 7629 3290
rect 7641 3238 7693 3290
rect 1032 3000 1084 3052
rect 4436 3000 4488 3052
rect 7104 3000 7156 3052
rect 1400 2932 1452 2984
rect 4528 2975 4580 2984
rect 4528 2941 4537 2975
rect 4537 2941 4571 2975
rect 4571 2941 4580 2975
rect 4528 2932 4580 2941
rect 7012 2932 7064 2984
rect 1110 2694 1162 2746
rect 1174 2694 1226 2746
rect 1238 2694 1290 2746
rect 1302 2694 1354 2746
rect 1366 2694 1418 2746
rect 2903 2694 2955 2746
rect 2967 2694 3019 2746
rect 3031 2694 3083 2746
rect 3095 2694 3147 2746
rect 3159 2694 3211 2746
rect 4696 2694 4748 2746
rect 4760 2694 4812 2746
rect 4824 2694 4876 2746
rect 4888 2694 4940 2746
rect 4952 2694 5004 2746
rect 6489 2694 6541 2746
rect 6553 2694 6605 2746
rect 6617 2694 6669 2746
rect 6681 2694 6733 2746
rect 6745 2694 6797 2746
rect 480 2524 532 2576
rect 6368 2524 6420 2576
rect 480 2388 532 2440
rect 6368 2388 6420 2440
rect 2006 2150 2058 2202
rect 2070 2150 2122 2202
rect 2134 2150 2186 2202
rect 2198 2150 2250 2202
rect 2262 2150 2314 2202
rect 3799 2150 3851 2202
rect 3863 2150 3915 2202
rect 3927 2150 3979 2202
rect 3991 2150 4043 2202
rect 4055 2150 4107 2202
rect 5592 2150 5644 2202
rect 5656 2150 5708 2202
rect 5720 2150 5772 2202
rect 5784 2150 5836 2202
rect 5848 2150 5900 2202
rect 7385 2150 7437 2202
rect 7449 2150 7501 2202
rect 7513 2150 7565 2202
rect 7577 2150 7629 2202
rect 7641 2150 7693 2202
rect 848 1912 900 1964
rect 2412 1912 2464 1964
rect 940 1887 992 1896
rect 940 1853 949 1887
rect 949 1853 983 1887
rect 983 1853 992 1887
rect 940 1844 992 1853
rect 2504 1887 2556 1896
rect 2504 1853 2513 1887
rect 2513 1853 2547 1887
rect 2547 1853 2556 1887
rect 2504 1844 2556 1853
rect 5540 1912 5592 1964
rect 6092 1844 6144 1896
rect 6184 1887 6236 1896
rect 6184 1853 6193 1887
rect 6193 1853 6227 1887
rect 6227 1853 6236 1887
rect 6184 1844 6236 1853
rect 6276 1776 6328 1828
rect 1110 1606 1162 1658
rect 1174 1606 1226 1658
rect 1238 1606 1290 1658
rect 1302 1606 1354 1658
rect 1366 1606 1418 1658
rect 2903 1606 2955 1658
rect 2967 1606 3019 1658
rect 3031 1606 3083 1658
rect 3095 1606 3147 1658
rect 3159 1606 3211 1658
rect 4696 1606 4748 1658
rect 4760 1606 4812 1658
rect 4824 1606 4876 1658
rect 4888 1606 4940 1658
rect 4952 1606 5004 1658
rect 6489 1606 6541 1658
rect 6553 1606 6605 1658
rect 6617 1606 6669 1658
rect 6681 1606 6733 1658
rect 6745 1606 6797 1658
rect 1584 1300 1636 1352
rect 1676 1300 1728 1352
rect 6736 1343 6788 1352
rect 6736 1309 6745 1343
rect 6745 1309 6779 1343
rect 6779 1309 6788 1343
rect 6736 1300 6788 1309
rect 6828 1232 6880 1284
rect 2006 1062 2058 1114
rect 2070 1062 2122 1114
rect 2134 1062 2186 1114
rect 2198 1062 2250 1114
rect 2262 1062 2314 1114
rect 3799 1062 3851 1114
rect 3863 1062 3915 1114
rect 3927 1062 3979 1114
rect 3991 1062 4043 1114
rect 4055 1062 4107 1114
rect 5592 1062 5644 1114
rect 5656 1062 5708 1114
rect 5720 1062 5772 1114
rect 5784 1062 5836 1114
rect 5848 1062 5900 1114
rect 7385 1062 7437 1114
rect 7449 1062 7501 1114
rect 7513 1062 7565 1114
rect 7577 1062 7629 1114
rect 7641 1062 7693 1114
<< metal2 >>
rect 478 5200 534 6000
rect 846 5200 902 6000
rect 1214 5200 1270 6000
rect 1582 5200 1638 6000
rect 1950 5200 2006 6000
rect 2318 5200 2374 6000
rect 2686 5200 2742 6000
rect 3054 5200 3110 6000
rect 3422 5200 3478 6000
rect 3790 5200 3846 6000
rect 4158 5200 4214 6000
rect 4526 5200 4582 6000
rect 4632 5222 4844 5250
rect 492 2582 520 5200
rect 860 3618 888 5200
rect 1228 5114 1256 5200
rect 1044 5086 1256 5114
rect 860 3590 980 3618
rect 480 2576 532 2582
rect 480 2518 532 2524
rect 480 2440 532 2446
rect 480 2382 532 2388
rect 492 800 520 2382
rect 848 1964 900 1970
rect 848 1906 900 1912
rect 860 800 888 1906
rect 952 1902 980 3590
rect 1044 3210 1072 5086
rect 1110 4924 1418 4933
rect 1110 4922 1116 4924
rect 1172 4922 1196 4924
rect 1252 4922 1276 4924
rect 1332 4922 1356 4924
rect 1412 4922 1418 4924
rect 1172 4870 1174 4922
rect 1354 4870 1356 4922
rect 1110 4868 1116 4870
rect 1172 4868 1196 4870
rect 1252 4868 1276 4870
rect 1332 4868 1356 4870
rect 1412 4868 1418 4870
rect 1110 4859 1418 4868
rect 1110 3836 1418 3845
rect 1110 3834 1116 3836
rect 1172 3834 1196 3836
rect 1252 3834 1276 3836
rect 1332 3834 1356 3836
rect 1412 3834 1418 3836
rect 1172 3782 1174 3834
rect 1354 3782 1356 3834
rect 1110 3780 1116 3782
rect 1172 3780 1196 3782
rect 1252 3780 1276 3782
rect 1332 3780 1356 3782
rect 1412 3780 1418 3782
rect 1110 3771 1418 3780
rect 1044 3182 1440 3210
rect 1032 3052 1084 3058
rect 1032 2994 1084 3000
rect 940 1896 992 1902
rect 940 1838 992 1844
rect 1044 1442 1072 2994
rect 1412 2990 1440 3182
rect 1400 2984 1452 2990
rect 1400 2926 1452 2932
rect 1110 2748 1418 2757
rect 1110 2746 1116 2748
rect 1172 2746 1196 2748
rect 1252 2746 1276 2748
rect 1332 2746 1356 2748
rect 1412 2746 1418 2748
rect 1172 2694 1174 2746
rect 1354 2694 1356 2746
rect 1110 2692 1116 2694
rect 1172 2692 1196 2694
rect 1252 2692 1276 2694
rect 1332 2692 1356 2694
rect 1412 2692 1418 2694
rect 1110 2683 1418 2692
rect 1596 2666 1624 5200
rect 1964 4570 1992 5200
rect 1872 4542 1992 4570
rect 2332 4570 2360 5200
rect 2332 4542 2544 4570
rect 1872 3602 1900 4542
rect 2006 4380 2314 4389
rect 2006 4378 2012 4380
rect 2068 4378 2092 4380
rect 2148 4378 2172 4380
rect 2228 4378 2252 4380
rect 2308 4378 2314 4380
rect 2068 4326 2070 4378
rect 2250 4326 2252 4378
rect 2006 4324 2012 4326
rect 2068 4324 2092 4326
rect 2148 4324 2172 4326
rect 2228 4324 2252 4326
rect 2308 4324 2314 4326
rect 2006 4315 2314 4324
rect 1860 3596 1912 3602
rect 1860 3538 1912 3544
rect 1860 3460 1912 3466
rect 1860 3402 1912 3408
rect 1596 2638 1716 2666
rect 1110 1660 1418 1669
rect 1110 1658 1116 1660
rect 1172 1658 1196 1660
rect 1252 1658 1276 1660
rect 1332 1658 1356 1660
rect 1412 1658 1418 1660
rect 1172 1606 1174 1658
rect 1354 1606 1356 1658
rect 1110 1604 1116 1606
rect 1172 1604 1196 1606
rect 1252 1604 1276 1606
rect 1332 1604 1356 1606
rect 1412 1604 1418 1606
rect 1110 1595 1418 1604
rect 1044 1414 1256 1442
rect 1228 800 1256 1414
rect 1688 1358 1716 2638
rect 1584 1352 1636 1358
rect 1584 1294 1636 1300
rect 1676 1352 1728 1358
rect 1676 1294 1728 1300
rect 1596 800 1624 1294
rect 1872 898 1900 3402
rect 2006 3292 2314 3301
rect 2006 3290 2012 3292
rect 2068 3290 2092 3292
rect 2148 3290 2172 3292
rect 2228 3290 2252 3292
rect 2308 3290 2314 3292
rect 2068 3238 2070 3290
rect 2250 3238 2252 3290
rect 2006 3236 2012 3238
rect 2068 3236 2092 3238
rect 2148 3236 2172 3238
rect 2228 3236 2252 3238
rect 2308 3236 2314 3238
rect 2006 3227 2314 3236
rect 2006 2204 2314 2213
rect 2006 2202 2012 2204
rect 2068 2202 2092 2204
rect 2148 2202 2172 2204
rect 2228 2202 2252 2204
rect 2308 2202 2314 2204
rect 2068 2150 2070 2202
rect 2250 2150 2252 2202
rect 2006 2148 2012 2150
rect 2068 2148 2092 2150
rect 2148 2148 2172 2150
rect 2228 2148 2252 2150
rect 2308 2148 2314 2150
rect 2006 2139 2314 2148
rect 2412 1964 2464 1970
rect 2412 1906 2464 1912
rect 2006 1116 2314 1125
rect 2006 1114 2012 1116
rect 2068 1114 2092 1116
rect 2148 1114 2172 1116
rect 2228 1114 2252 1116
rect 2308 1114 2314 1116
rect 2068 1062 2070 1114
rect 2250 1062 2252 1114
rect 2006 1060 2012 1062
rect 2068 1060 2092 1062
rect 2148 1060 2172 1062
rect 2228 1060 2252 1062
rect 2308 1060 2314 1062
rect 2006 1051 2314 1060
rect 2424 898 2452 1906
rect 2516 1902 2544 4542
rect 2700 4298 2728 5200
rect 3068 5114 3096 5200
rect 3068 5086 3280 5114
rect 2903 4924 3211 4933
rect 2903 4922 2909 4924
rect 2965 4922 2989 4924
rect 3045 4922 3069 4924
rect 3125 4922 3149 4924
rect 3205 4922 3211 4924
rect 2965 4870 2967 4922
rect 3147 4870 3149 4922
rect 2903 4868 2909 4870
rect 2965 4868 2989 4870
rect 3045 4868 3069 4870
rect 3125 4868 3149 4870
rect 3205 4868 3211 4870
rect 2903 4859 3211 4868
rect 3252 4758 3280 5086
rect 3240 4752 3292 4758
rect 3436 4706 3464 5200
rect 3240 4694 3292 4700
rect 3344 4678 3464 4706
rect 3240 4616 3292 4622
rect 3240 4558 3292 4564
rect 2608 4270 2728 4298
rect 2608 4078 2636 4270
rect 2688 4140 2740 4146
rect 2688 4082 2740 4088
rect 2596 4072 2648 4078
rect 2596 4014 2648 4020
rect 2504 1896 2556 1902
rect 2504 1838 2556 1844
rect 1872 870 1992 898
rect 1964 800 1992 870
rect 2332 870 2452 898
rect 2332 800 2360 870
rect 2700 800 2728 4082
rect 2903 3836 3211 3845
rect 2903 3834 2909 3836
rect 2965 3834 2989 3836
rect 3045 3834 3069 3836
rect 3125 3834 3149 3836
rect 3205 3834 3211 3836
rect 2965 3782 2967 3834
rect 3147 3782 3149 3834
rect 2903 3780 2909 3782
rect 2965 3780 2989 3782
rect 3045 3780 3069 3782
rect 3125 3780 3149 3782
rect 3205 3780 3211 3782
rect 2903 3771 3211 3780
rect 2903 2748 3211 2757
rect 2903 2746 2909 2748
rect 2965 2746 2989 2748
rect 3045 2746 3069 2748
rect 3125 2746 3149 2748
rect 3205 2746 3211 2748
rect 2965 2694 2967 2746
rect 3147 2694 3149 2746
rect 2903 2692 2909 2694
rect 2965 2692 2989 2694
rect 3045 2692 3069 2694
rect 3125 2692 3149 2694
rect 3205 2692 3211 2694
rect 2903 2683 3211 2692
rect 2903 1660 3211 1669
rect 2903 1658 2909 1660
rect 2965 1658 2989 1660
rect 3045 1658 3069 1660
rect 3125 1658 3149 1660
rect 3205 1658 3211 1660
rect 2965 1606 2967 1658
rect 3147 1606 3149 1658
rect 2903 1604 2909 1606
rect 2965 1604 2989 1606
rect 3045 1604 3069 1606
rect 3125 1604 3149 1606
rect 3205 1604 3211 1606
rect 2903 1595 3211 1604
rect 3252 1442 3280 4558
rect 3344 4078 3372 4678
rect 3804 4570 3832 5200
rect 3712 4542 3832 4570
rect 3424 4140 3476 4146
rect 3424 4082 3476 4088
rect 3332 4072 3384 4078
rect 3332 4014 3384 4020
rect 3068 1414 3280 1442
rect 3068 800 3096 1414
rect 3436 800 3464 4082
rect 3712 3670 3740 4542
rect 3799 4380 4107 4389
rect 3799 4378 3805 4380
rect 3861 4378 3885 4380
rect 3941 4378 3965 4380
rect 4021 4378 4045 4380
rect 4101 4378 4107 4380
rect 3861 4326 3863 4378
rect 4043 4326 4045 4378
rect 3799 4324 3805 4326
rect 3861 4324 3885 4326
rect 3941 4324 3965 4326
rect 4021 4324 4045 4326
rect 4101 4324 4107 4326
rect 3799 4315 4107 4324
rect 4172 3670 4200 5200
rect 3700 3664 3752 3670
rect 3700 3606 3752 3612
rect 4160 3664 4212 3670
rect 4160 3606 4212 3612
rect 3700 3528 3752 3534
rect 3700 3470 3752 3476
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 3712 898 3740 3470
rect 3799 3292 4107 3301
rect 3799 3290 3805 3292
rect 3861 3290 3885 3292
rect 3941 3290 3965 3292
rect 4021 3290 4045 3292
rect 4101 3290 4107 3292
rect 3861 3238 3863 3290
rect 4043 3238 4045 3290
rect 3799 3236 3805 3238
rect 3861 3236 3885 3238
rect 3941 3236 3965 3238
rect 4021 3236 4045 3238
rect 4101 3236 4107 3238
rect 3799 3227 4107 3236
rect 3799 2204 4107 2213
rect 3799 2202 3805 2204
rect 3861 2202 3885 2204
rect 3941 2202 3965 2204
rect 4021 2202 4045 2204
rect 4101 2202 4107 2204
rect 3861 2150 3863 2202
rect 4043 2150 4045 2202
rect 3799 2148 3805 2150
rect 3861 2148 3885 2150
rect 3941 2148 3965 2150
rect 4021 2148 4045 2150
rect 4101 2148 4107 2150
rect 3799 2139 4107 2148
rect 3799 1116 4107 1125
rect 3799 1114 3805 1116
rect 3861 1114 3885 1116
rect 3941 1114 3965 1116
rect 4021 1114 4045 1116
rect 4101 1114 4107 1116
rect 3861 1062 3863 1114
rect 4043 1062 4045 1114
rect 3799 1060 3805 1062
rect 3861 1060 3885 1062
rect 3941 1060 3965 1062
rect 4021 1060 4045 1062
rect 4101 1060 4107 1062
rect 3799 1051 4107 1060
rect 3712 870 3832 898
rect 3804 800 3832 870
rect 4172 800 4200 3470
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 4448 2802 4476 2994
rect 4540 2990 4568 5200
rect 4632 4078 4660 5222
rect 4816 5114 4844 5222
rect 4894 5200 4950 6000
rect 5262 5200 5318 6000
rect 5630 5200 5686 6000
rect 5736 5222 5948 5250
rect 4908 5114 4936 5200
rect 4816 5086 4936 5114
rect 4696 4924 5004 4933
rect 4696 4922 4702 4924
rect 4758 4922 4782 4924
rect 4838 4922 4862 4924
rect 4918 4922 4942 4924
rect 4998 4922 5004 4924
rect 4758 4870 4760 4922
rect 4940 4870 4942 4922
rect 4696 4868 4702 4870
rect 4758 4868 4782 4870
rect 4838 4868 4862 4870
rect 4918 4868 4942 4870
rect 4998 4868 5004 4870
rect 4696 4859 5004 4868
rect 5276 4298 5304 5200
rect 5644 5114 5672 5200
rect 5736 5114 5764 5222
rect 5644 5086 5764 5114
rect 5920 4570 5948 5222
rect 5998 5200 6054 6000
rect 6104 5222 6316 5250
rect 6012 5114 6040 5200
rect 6104 5114 6132 5222
rect 6012 5086 6132 5114
rect 5920 4542 6224 4570
rect 5592 4380 5900 4389
rect 5592 4378 5598 4380
rect 5654 4378 5678 4380
rect 5734 4378 5758 4380
rect 5814 4378 5838 4380
rect 5894 4378 5900 4380
rect 5654 4326 5656 4378
rect 5836 4326 5838 4378
rect 5592 4324 5598 4326
rect 5654 4324 5678 4326
rect 5734 4324 5758 4326
rect 5814 4324 5838 4326
rect 5894 4324 5900 4326
rect 5592 4315 5900 4324
rect 5276 4270 5488 4298
rect 5080 4140 5132 4146
rect 5080 4082 5132 4088
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 4620 4072 4672 4078
rect 4620 4014 4672 4020
rect 4696 3836 5004 3845
rect 4696 3834 4702 3836
rect 4758 3834 4782 3836
rect 4838 3834 4862 3836
rect 4918 3834 4942 3836
rect 4998 3834 5004 3836
rect 4758 3782 4760 3834
rect 4940 3782 4942 3834
rect 4696 3780 4702 3782
rect 4758 3780 4782 3782
rect 4838 3780 4862 3782
rect 4918 3780 4942 3782
rect 4998 3780 5004 3782
rect 4696 3771 5004 3780
rect 4528 2984 4580 2990
rect 4528 2926 4580 2932
rect 4448 2774 4568 2802
rect 4540 800 4568 2774
rect 4696 2748 5004 2757
rect 4696 2746 4702 2748
rect 4758 2746 4782 2748
rect 4838 2746 4862 2748
rect 4918 2746 4942 2748
rect 4998 2746 5004 2748
rect 4758 2694 4760 2746
rect 4940 2694 4942 2746
rect 4696 2692 4702 2694
rect 4758 2692 4782 2694
rect 4838 2692 4862 2694
rect 4918 2692 4942 2694
rect 4998 2692 5004 2694
rect 4696 2683 5004 2692
rect 4696 1660 5004 1669
rect 4696 1658 4702 1660
rect 4758 1658 4782 1660
rect 4838 1658 4862 1660
rect 4918 1658 4942 1660
rect 4998 1658 5004 1660
rect 4758 1606 4760 1658
rect 4940 1606 4942 1658
rect 4696 1604 4702 1606
rect 4758 1604 4782 1606
rect 4838 1604 4862 1606
rect 4918 1604 4942 1606
rect 4998 1604 5004 1606
rect 4696 1595 5004 1604
rect 5092 1442 5120 4082
rect 4908 1414 5120 1442
rect 4908 800 4936 1414
rect 5276 800 5304 4082
rect 5460 4026 5488 4270
rect 5540 4072 5592 4078
rect 5460 4020 5540 4026
rect 5460 4014 5592 4020
rect 5460 3998 5580 4014
rect 5592 3292 5900 3301
rect 5592 3290 5598 3292
rect 5654 3290 5678 3292
rect 5734 3290 5758 3292
rect 5814 3290 5838 3292
rect 5894 3290 5900 3292
rect 5654 3238 5656 3290
rect 5836 3238 5838 3290
rect 5592 3236 5598 3238
rect 5654 3236 5678 3238
rect 5734 3236 5758 3238
rect 5814 3236 5838 3238
rect 5894 3236 5900 3238
rect 5592 3227 5900 3236
rect 5592 2204 5900 2213
rect 5592 2202 5598 2204
rect 5654 2202 5678 2204
rect 5734 2202 5758 2204
rect 5814 2202 5838 2204
rect 5894 2202 5900 2204
rect 5654 2150 5656 2202
rect 5836 2150 5838 2202
rect 5592 2148 5598 2150
rect 5654 2148 5678 2150
rect 5734 2148 5758 2150
rect 5814 2148 5838 2150
rect 5894 2148 5900 2150
rect 5592 2139 5900 2148
rect 5540 1964 5592 1970
rect 5540 1906 5592 1912
rect 5552 1306 5580 1906
rect 6196 1902 6224 4542
rect 6092 1896 6144 1902
rect 6092 1838 6144 1844
rect 6184 1896 6236 1902
rect 6184 1838 6236 1844
rect 5460 1278 5580 1306
rect 5460 898 5488 1278
rect 5592 1116 5900 1125
rect 5592 1114 5598 1116
rect 5654 1114 5678 1116
rect 5734 1114 5758 1116
rect 5814 1114 5838 1116
rect 5894 1114 5900 1116
rect 5654 1062 5656 1114
rect 5836 1062 5838 1114
rect 5592 1060 5598 1062
rect 5654 1060 5678 1062
rect 5734 1060 5758 1062
rect 5814 1060 5838 1062
rect 5894 1060 5900 1062
rect 5592 1051 5900 1060
rect 6104 898 6132 1838
rect 6288 1834 6316 5222
rect 6366 5200 6422 6000
rect 6734 5200 6790 6000
rect 7102 5200 7158 6000
rect 7470 5200 7526 6000
rect 6380 2582 6408 5200
rect 6748 5114 6776 5200
rect 6748 5086 6868 5114
rect 6489 4924 6797 4933
rect 6489 4922 6495 4924
rect 6551 4922 6575 4924
rect 6631 4922 6655 4924
rect 6711 4922 6735 4924
rect 6791 4922 6797 4924
rect 6551 4870 6553 4922
rect 6733 4870 6735 4922
rect 6489 4868 6495 4870
rect 6551 4868 6575 4870
rect 6631 4868 6655 4870
rect 6711 4868 6735 4870
rect 6791 4868 6797 4870
rect 6489 4859 6797 4868
rect 6489 3836 6797 3845
rect 6489 3834 6495 3836
rect 6551 3834 6575 3836
rect 6631 3834 6655 3836
rect 6711 3834 6735 3836
rect 6791 3834 6797 3836
rect 6551 3782 6553 3834
rect 6733 3782 6735 3834
rect 6489 3780 6495 3782
rect 6551 3780 6575 3782
rect 6631 3780 6655 3782
rect 6711 3780 6735 3782
rect 6791 3780 6797 3782
rect 6489 3771 6797 3780
rect 6489 2748 6797 2757
rect 6489 2746 6495 2748
rect 6551 2746 6575 2748
rect 6631 2746 6655 2748
rect 6711 2746 6735 2748
rect 6791 2746 6797 2748
rect 6551 2694 6553 2746
rect 6733 2694 6735 2746
rect 6489 2692 6495 2694
rect 6551 2692 6575 2694
rect 6631 2692 6655 2694
rect 6711 2692 6735 2694
rect 6791 2692 6797 2694
rect 6489 2683 6797 2692
rect 6368 2576 6420 2582
rect 6368 2518 6420 2524
rect 6368 2440 6420 2446
rect 6368 2382 6420 2388
rect 6276 1828 6328 1834
rect 6276 1770 6328 1776
rect 5460 870 5672 898
rect 5644 800 5672 870
rect 6012 870 6132 898
rect 6012 800 6040 870
rect 6380 800 6408 2382
rect 6489 1660 6797 1669
rect 6489 1658 6495 1660
rect 6551 1658 6575 1660
rect 6631 1658 6655 1660
rect 6711 1658 6735 1660
rect 6791 1658 6797 1660
rect 6551 1606 6553 1658
rect 6733 1606 6735 1658
rect 6489 1604 6495 1606
rect 6551 1604 6575 1606
rect 6631 1604 6655 1606
rect 6711 1604 6735 1606
rect 6791 1604 6797 1606
rect 6489 1595 6797 1604
rect 6736 1352 6788 1358
rect 6736 1294 6788 1300
rect 6748 800 6776 1294
rect 6840 1290 6868 5086
rect 7116 3210 7144 5200
rect 7484 4690 7512 5200
rect 7472 4684 7524 4690
rect 7472 4626 7524 4632
rect 7288 4616 7340 4622
rect 7288 4558 7340 4564
rect 7024 3182 7144 3210
rect 7024 2990 7052 3182
rect 7104 3052 7156 3058
rect 7104 2994 7156 3000
rect 7012 2984 7064 2990
rect 7012 2926 7064 2932
rect 6828 1284 6880 1290
rect 6828 1226 6880 1232
rect 7116 800 7144 2994
rect 7300 898 7328 4558
rect 7385 4380 7693 4389
rect 7385 4378 7391 4380
rect 7447 4378 7471 4380
rect 7527 4378 7551 4380
rect 7607 4378 7631 4380
rect 7687 4378 7693 4380
rect 7447 4326 7449 4378
rect 7629 4326 7631 4378
rect 7385 4324 7391 4326
rect 7447 4324 7471 4326
rect 7527 4324 7551 4326
rect 7607 4324 7631 4326
rect 7687 4324 7693 4326
rect 7385 4315 7693 4324
rect 7385 3292 7693 3301
rect 7385 3290 7391 3292
rect 7447 3290 7471 3292
rect 7527 3290 7551 3292
rect 7607 3290 7631 3292
rect 7687 3290 7693 3292
rect 7447 3238 7449 3290
rect 7629 3238 7631 3290
rect 7385 3236 7391 3238
rect 7447 3236 7471 3238
rect 7527 3236 7551 3238
rect 7607 3236 7631 3238
rect 7687 3236 7693 3238
rect 7385 3227 7693 3236
rect 7385 2204 7693 2213
rect 7385 2202 7391 2204
rect 7447 2202 7471 2204
rect 7527 2202 7551 2204
rect 7607 2202 7631 2204
rect 7687 2202 7693 2204
rect 7447 2150 7449 2202
rect 7629 2150 7631 2202
rect 7385 2148 7391 2150
rect 7447 2148 7471 2150
rect 7527 2148 7551 2150
rect 7607 2148 7631 2150
rect 7687 2148 7693 2150
rect 7385 2139 7693 2148
rect 7385 1116 7693 1125
rect 7385 1114 7391 1116
rect 7447 1114 7471 1116
rect 7527 1114 7551 1116
rect 7607 1114 7631 1116
rect 7687 1114 7693 1116
rect 7447 1062 7449 1114
rect 7629 1062 7631 1114
rect 7385 1060 7391 1062
rect 7447 1060 7471 1062
rect 7527 1060 7551 1062
rect 7607 1060 7631 1062
rect 7687 1060 7693 1062
rect 7385 1051 7693 1060
rect 7300 870 7512 898
rect 7484 800 7512 870
rect 478 0 534 800
rect 846 0 902 800
rect 1214 0 1270 800
rect 1582 0 1638 800
rect 1950 0 2006 800
rect 2318 0 2374 800
rect 2686 0 2742 800
rect 3054 0 3110 800
rect 3422 0 3478 800
rect 3790 0 3846 800
rect 4158 0 4214 800
rect 4526 0 4582 800
rect 4894 0 4950 800
rect 5262 0 5318 800
rect 5630 0 5686 800
rect 5998 0 6054 800
rect 6366 0 6422 800
rect 6734 0 6790 800
rect 7102 0 7158 800
rect 7470 0 7526 800
<< via2 >>
rect 1116 4922 1172 4924
rect 1196 4922 1252 4924
rect 1276 4922 1332 4924
rect 1356 4922 1412 4924
rect 1116 4870 1162 4922
rect 1162 4870 1172 4922
rect 1196 4870 1226 4922
rect 1226 4870 1238 4922
rect 1238 4870 1252 4922
rect 1276 4870 1290 4922
rect 1290 4870 1302 4922
rect 1302 4870 1332 4922
rect 1356 4870 1366 4922
rect 1366 4870 1412 4922
rect 1116 4868 1172 4870
rect 1196 4868 1252 4870
rect 1276 4868 1332 4870
rect 1356 4868 1412 4870
rect 1116 3834 1172 3836
rect 1196 3834 1252 3836
rect 1276 3834 1332 3836
rect 1356 3834 1412 3836
rect 1116 3782 1162 3834
rect 1162 3782 1172 3834
rect 1196 3782 1226 3834
rect 1226 3782 1238 3834
rect 1238 3782 1252 3834
rect 1276 3782 1290 3834
rect 1290 3782 1302 3834
rect 1302 3782 1332 3834
rect 1356 3782 1366 3834
rect 1366 3782 1412 3834
rect 1116 3780 1172 3782
rect 1196 3780 1252 3782
rect 1276 3780 1332 3782
rect 1356 3780 1412 3782
rect 1116 2746 1172 2748
rect 1196 2746 1252 2748
rect 1276 2746 1332 2748
rect 1356 2746 1412 2748
rect 1116 2694 1162 2746
rect 1162 2694 1172 2746
rect 1196 2694 1226 2746
rect 1226 2694 1238 2746
rect 1238 2694 1252 2746
rect 1276 2694 1290 2746
rect 1290 2694 1302 2746
rect 1302 2694 1332 2746
rect 1356 2694 1366 2746
rect 1366 2694 1412 2746
rect 1116 2692 1172 2694
rect 1196 2692 1252 2694
rect 1276 2692 1332 2694
rect 1356 2692 1412 2694
rect 2012 4378 2068 4380
rect 2092 4378 2148 4380
rect 2172 4378 2228 4380
rect 2252 4378 2308 4380
rect 2012 4326 2058 4378
rect 2058 4326 2068 4378
rect 2092 4326 2122 4378
rect 2122 4326 2134 4378
rect 2134 4326 2148 4378
rect 2172 4326 2186 4378
rect 2186 4326 2198 4378
rect 2198 4326 2228 4378
rect 2252 4326 2262 4378
rect 2262 4326 2308 4378
rect 2012 4324 2068 4326
rect 2092 4324 2148 4326
rect 2172 4324 2228 4326
rect 2252 4324 2308 4326
rect 1116 1658 1172 1660
rect 1196 1658 1252 1660
rect 1276 1658 1332 1660
rect 1356 1658 1412 1660
rect 1116 1606 1162 1658
rect 1162 1606 1172 1658
rect 1196 1606 1226 1658
rect 1226 1606 1238 1658
rect 1238 1606 1252 1658
rect 1276 1606 1290 1658
rect 1290 1606 1302 1658
rect 1302 1606 1332 1658
rect 1356 1606 1366 1658
rect 1366 1606 1412 1658
rect 1116 1604 1172 1606
rect 1196 1604 1252 1606
rect 1276 1604 1332 1606
rect 1356 1604 1412 1606
rect 2012 3290 2068 3292
rect 2092 3290 2148 3292
rect 2172 3290 2228 3292
rect 2252 3290 2308 3292
rect 2012 3238 2058 3290
rect 2058 3238 2068 3290
rect 2092 3238 2122 3290
rect 2122 3238 2134 3290
rect 2134 3238 2148 3290
rect 2172 3238 2186 3290
rect 2186 3238 2198 3290
rect 2198 3238 2228 3290
rect 2252 3238 2262 3290
rect 2262 3238 2308 3290
rect 2012 3236 2068 3238
rect 2092 3236 2148 3238
rect 2172 3236 2228 3238
rect 2252 3236 2308 3238
rect 2012 2202 2068 2204
rect 2092 2202 2148 2204
rect 2172 2202 2228 2204
rect 2252 2202 2308 2204
rect 2012 2150 2058 2202
rect 2058 2150 2068 2202
rect 2092 2150 2122 2202
rect 2122 2150 2134 2202
rect 2134 2150 2148 2202
rect 2172 2150 2186 2202
rect 2186 2150 2198 2202
rect 2198 2150 2228 2202
rect 2252 2150 2262 2202
rect 2262 2150 2308 2202
rect 2012 2148 2068 2150
rect 2092 2148 2148 2150
rect 2172 2148 2228 2150
rect 2252 2148 2308 2150
rect 2012 1114 2068 1116
rect 2092 1114 2148 1116
rect 2172 1114 2228 1116
rect 2252 1114 2308 1116
rect 2012 1062 2058 1114
rect 2058 1062 2068 1114
rect 2092 1062 2122 1114
rect 2122 1062 2134 1114
rect 2134 1062 2148 1114
rect 2172 1062 2186 1114
rect 2186 1062 2198 1114
rect 2198 1062 2228 1114
rect 2252 1062 2262 1114
rect 2262 1062 2308 1114
rect 2012 1060 2068 1062
rect 2092 1060 2148 1062
rect 2172 1060 2228 1062
rect 2252 1060 2308 1062
rect 2909 4922 2965 4924
rect 2989 4922 3045 4924
rect 3069 4922 3125 4924
rect 3149 4922 3205 4924
rect 2909 4870 2955 4922
rect 2955 4870 2965 4922
rect 2989 4870 3019 4922
rect 3019 4870 3031 4922
rect 3031 4870 3045 4922
rect 3069 4870 3083 4922
rect 3083 4870 3095 4922
rect 3095 4870 3125 4922
rect 3149 4870 3159 4922
rect 3159 4870 3205 4922
rect 2909 4868 2965 4870
rect 2989 4868 3045 4870
rect 3069 4868 3125 4870
rect 3149 4868 3205 4870
rect 2909 3834 2965 3836
rect 2989 3834 3045 3836
rect 3069 3834 3125 3836
rect 3149 3834 3205 3836
rect 2909 3782 2955 3834
rect 2955 3782 2965 3834
rect 2989 3782 3019 3834
rect 3019 3782 3031 3834
rect 3031 3782 3045 3834
rect 3069 3782 3083 3834
rect 3083 3782 3095 3834
rect 3095 3782 3125 3834
rect 3149 3782 3159 3834
rect 3159 3782 3205 3834
rect 2909 3780 2965 3782
rect 2989 3780 3045 3782
rect 3069 3780 3125 3782
rect 3149 3780 3205 3782
rect 2909 2746 2965 2748
rect 2989 2746 3045 2748
rect 3069 2746 3125 2748
rect 3149 2746 3205 2748
rect 2909 2694 2955 2746
rect 2955 2694 2965 2746
rect 2989 2694 3019 2746
rect 3019 2694 3031 2746
rect 3031 2694 3045 2746
rect 3069 2694 3083 2746
rect 3083 2694 3095 2746
rect 3095 2694 3125 2746
rect 3149 2694 3159 2746
rect 3159 2694 3205 2746
rect 2909 2692 2965 2694
rect 2989 2692 3045 2694
rect 3069 2692 3125 2694
rect 3149 2692 3205 2694
rect 2909 1658 2965 1660
rect 2989 1658 3045 1660
rect 3069 1658 3125 1660
rect 3149 1658 3205 1660
rect 2909 1606 2955 1658
rect 2955 1606 2965 1658
rect 2989 1606 3019 1658
rect 3019 1606 3031 1658
rect 3031 1606 3045 1658
rect 3069 1606 3083 1658
rect 3083 1606 3095 1658
rect 3095 1606 3125 1658
rect 3149 1606 3159 1658
rect 3159 1606 3205 1658
rect 2909 1604 2965 1606
rect 2989 1604 3045 1606
rect 3069 1604 3125 1606
rect 3149 1604 3205 1606
rect 3805 4378 3861 4380
rect 3885 4378 3941 4380
rect 3965 4378 4021 4380
rect 4045 4378 4101 4380
rect 3805 4326 3851 4378
rect 3851 4326 3861 4378
rect 3885 4326 3915 4378
rect 3915 4326 3927 4378
rect 3927 4326 3941 4378
rect 3965 4326 3979 4378
rect 3979 4326 3991 4378
rect 3991 4326 4021 4378
rect 4045 4326 4055 4378
rect 4055 4326 4101 4378
rect 3805 4324 3861 4326
rect 3885 4324 3941 4326
rect 3965 4324 4021 4326
rect 4045 4324 4101 4326
rect 3805 3290 3861 3292
rect 3885 3290 3941 3292
rect 3965 3290 4021 3292
rect 4045 3290 4101 3292
rect 3805 3238 3851 3290
rect 3851 3238 3861 3290
rect 3885 3238 3915 3290
rect 3915 3238 3927 3290
rect 3927 3238 3941 3290
rect 3965 3238 3979 3290
rect 3979 3238 3991 3290
rect 3991 3238 4021 3290
rect 4045 3238 4055 3290
rect 4055 3238 4101 3290
rect 3805 3236 3861 3238
rect 3885 3236 3941 3238
rect 3965 3236 4021 3238
rect 4045 3236 4101 3238
rect 3805 2202 3861 2204
rect 3885 2202 3941 2204
rect 3965 2202 4021 2204
rect 4045 2202 4101 2204
rect 3805 2150 3851 2202
rect 3851 2150 3861 2202
rect 3885 2150 3915 2202
rect 3915 2150 3927 2202
rect 3927 2150 3941 2202
rect 3965 2150 3979 2202
rect 3979 2150 3991 2202
rect 3991 2150 4021 2202
rect 4045 2150 4055 2202
rect 4055 2150 4101 2202
rect 3805 2148 3861 2150
rect 3885 2148 3941 2150
rect 3965 2148 4021 2150
rect 4045 2148 4101 2150
rect 3805 1114 3861 1116
rect 3885 1114 3941 1116
rect 3965 1114 4021 1116
rect 4045 1114 4101 1116
rect 3805 1062 3851 1114
rect 3851 1062 3861 1114
rect 3885 1062 3915 1114
rect 3915 1062 3927 1114
rect 3927 1062 3941 1114
rect 3965 1062 3979 1114
rect 3979 1062 3991 1114
rect 3991 1062 4021 1114
rect 4045 1062 4055 1114
rect 4055 1062 4101 1114
rect 3805 1060 3861 1062
rect 3885 1060 3941 1062
rect 3965 1060 4021 1062
rect 4045 1060 4101 1062
rect 4702 4922 4758 4924
rect 4782 4922 4838 4924
rect 4862 4922 4918 4924
rect 4942 4922 4998 4924
rect 4702 4870 4748 4922
rect 4748 4870 4758 4922
rect 4782 4870 4812 4922
rect 4812 4870 4824 4922
rect 4824 4870 4838 4922
rect 4862 4870 4876 4922
rect 4876 4870 4888 4922
rect 4888 4870 4918 4922
rect 4942 4870 4952 4922
rect 4952 4870 4998 4922
rect 4702 4868 4758 4870
rect 4782 4868 4838 4870
rect 4862 4868 4918 4870
rect 4942 4868 4998 4870
rect 5598 4378 5654 4380
rect 5678 4378 5734 4380
rect 5758 4378 5814 4380
rect 5838 4378 5894 4380
rect 5598 4326 5644 4378
rect 5644 4326 5654 4378
rect 5678 4326 5708 4378
rect 5708 4326 5720 4378
rect 5720 4326 5734 4378
rect 5758 4326 5772 4378
rect 5772 4326 5784 4378
rect 5784 4326 5814 4378
rect 5838 4326 5848 4378
rect 5848 4326 5894 4378
rect 5598 4324 5654 4326
rect 5678 4324 5734 4326
rect 5758 4324 5814 4326
rect 5838 4324 5894 4326
rect 4702 3834 4758 3836
rect 4782 3834 4838 3836
rect 4862 3834 4918 3836
rect 4942 3834 4998 3836
rect 4702 3782 4748 3834
rect 4748 3782 4758 3834
rect 4782 3782 4812 3834
rect 4812 3782 4824 3834
rect 4824 3782 4838 3834
rect 4862 3782 4876 3834
rect 4876 3782 4888 3834
rect 4888 3782 4918 3834
rect 4942 3782 4952 3834
rect 4952 3782 4998 3834
rect 4702 3780 4758 3782
rect 4782 3780 4838 3782
rect 4862 3780 4918 3782
rect 4942 3780 4998 3782
rect 4702 2746 4758 2748
rect 4782 2746 4838 2748
rect 4862 2746 4918 2748
rect 4942 2746 4998 2748
rect 4702 2694 4748 2746
rect 4748 2694 4758 2746
rect 4782 2694 4812 2746
rect 4812 2694 4824 2746
rect 4824 2694 4838 2746
rect 4862 2694 4876 2746
rect 4876 2694 4888 2746
rect 4888 2694 4918 2746
rect 4942 2694 4952 2746
rect 4952 2694 4998 2746
rect 4702 2692 4758 2694
rect 4782 2692 4838 2694
rect 4862 2692 4918 2694
rect 4942 2692 4998 2694
rect 4702 1658 4758 1660
rect 4782 1658 4838 1660
rect 4862 1658 4918 1660
rect 4942 1658 4998 1660
rect 4702 1606 4748 1658
rect 4748 1606 4758 1658
rect 4782 1606 4812 1658
rect 4812 1606 4824 1658
rect 4824 1606 4838 1658
rect 4862 1606 4876 1658
rect 4876 1606 4888 1658
rect 4888 1606 4918 1658
rect 4942 1606 4952 1658
rect 4952 1606 4998 1658
rect 4702 1604 4758 1606
rect 4782 1604 4838 1606
rect 4862 1604 4918 1606
rect 4942 1604 4998 1606
rect 5598 3290 5654 3292
rect 5678 3290 5734 3292
rect 5758 3290 5814 3292
rect 5838 3290 5894 3292
rect 5598 3238 5644 3290
rect 5644 3238 5654 3290
rect 5678 3238 5708 3290
rect 5708 3238 5720 3290
rect 5720 3238 5734 3290
rect 5758 3238 5772 3290
rect 5772 3238 5784 3290
rect 5784 3238 5814 3290
rect 5838 3238 5848 3290
rect 5848 3238 5894 3290
rect 5598 3236 5654 3238
rect 5678 3236 5734 3238
rect 5758 3236 5814 3238
rect 5838 3236 5894 3238
rect 5598 2202 5654 2204
rect 5678 2202 5734 2204
rect 5758 2202 5814 2204
rect 5838 2202 5894 2204
rect 5598 2150 5644 2202
rect 5644 2150 5654 2202
rect 5678 2150 5708 2202
rect 5708 2150 5720 2202
rect 5720 2150 5734 2202
rect 5758 2150 5772 2202
rect 5772 2150 5784 2202
rect 5784 2150 5814 2202
rect 5838 2150 5848 2202
rect 5848 2150 5894 2202
rect 5598 2148 5654 2150
rect 5678 2148 5734 2150
rect 5758 2148 5814 2150
rect 5838 2148 5894 2150
rect 5598 1114 5654 1116
rect 5678 1114 5734 1116
rect 5758 1114 5814 1116
rect 5838 1114 5894 1116
rect 5598 1062 5644 1114
rect 5644 1062 5654 1114
rect 5678 1062 5708 1114
rect 5708 1062 5720 1114
rect 5720 1062 5734 1114
rect 5758 1062 5772 1114
rect 5772 1062 5784 1114
rect 5784 1062 5814 1114
rect 5838 1062 5848 1114
rect 5848 1062 5894 1114
rect 5598 1060 5654 1062
rect 5678 1060 5734 1062
rect 5758 1060 5814 1062
rect 5838 1060 5894 1062
rect 6495 4922 6551 4924
rect 6575 4922 6631 4924
rect 6655 4922 6711 4924
rect 6735 4922 6791 4924
rect 6495 4870 6541 4922
rect 6541 4870 6551 4922
rect 6575 4870 6605 4922
rect 6605 4870 6617 4922
rect 6617 4870 6631 4922
rect 6655 4870 6669 4922
rect 6669 4870 6681 4922
rect 6681 4870 6711 4922
rect 6735 4870 6745 4922
rect 6745 4870 6791 4922
rect 6495 4868 6551 4870
rect 6575 4868 6631 4870
rect 6655 4868 6711 4870
rect 6735 4868 6791 4870
rect 6495 3834 6551 3836
rect 6575 3834 6631 3836
rect 6655 3834 6711 3836
rect 6735 3834 6791 3836
rect 6495 3782 6541 3834
rect 6541 3782 6551 3834
rect 6575 3782 6605 3834
rect 6605 3782 6617 3834
rect 6617 3782 6631 3834
rect 6655 3782 6669 3834
rect 6669 3782 6681 3834
rect 6681 3782 6711 3834
rect 6735 3782 6745 3834
rect 6745 3782 6791 3834
rect 6495 3780 6551 3782
rect 6575 3780 6631 3782
rect 6655 3780 6711 3782
rect 6735 3780 6791 3782
rect 6495 2746 6551 2748
rect 6575 2746 6631 2748
rect 6655 2746 6711 2748
rect 6735 2746 6791 2748
rect 6495 2694 6541 2746
rect 6541 2694 6551 2746
rect 6575 2694 6605 2746
rect 6605 2694 6617 2746
rect 6617 2694 6631 2746
rect 6655 2694 6669 2746
rect 6669 2694 6681 2746
rect 6681 2694 6711 2746
rect 6735 2694 6745 2746
rect 6745 2694 6791 2746
rect 6495 2692 6551 2694
rect 6575 2692 6631 2694
rect 6655 2692 6711 2694
rect 6735 2692 6791 2694
rect 6495 1658 6551 1660
rect 6575 1658 6631 1660
rect 6655 1658 6711 1660
rect 6735 1658 6791 1660
rect 6495 1606 6541 1658
rect 6541 1606 6551 1658
rect 6575 1606 6605 1658
rect 6605 1606 6617 1658
rect 6617 1606 6631 1658
rect 6655 1606 6669 1658
rect 6669 1606 6681 1658
rect 6681 1606 6711 1658
rect 6735 1606 6745 1658
rect 6745 1606 6791 1658
rect 6495 1604 6551 1606
rect 6575 1604 6631 1606
rect 6655 1604 6711 1606
rect 6735 1604 6791 1606
rect 7391 4378 7447 4380
rect 7471 4378 7527 4380
rect 7551 4378 7607 4380
rect 7631 4378 7687 4380
rect 7391 4326 7437 4378
rect 7437 4326 7447 4378
rect 7471 4326 7501 4378
rect 7501 4326 7513 4378
rect 7513 4326 7527 4378
rect 7551 4326 7565 4378
rect 7565 4326 7577 4378
rect 7577 4326 7607 4378
rect 7631 4326 7641 4378
rect 7641 4326 7687 4378
rect 7391 4324 7447 4326
rect 7471 4324 7527 4326
rect 7551 4324 7607 4326
rect 7631 4324 7687 4326
rect 7391 3290 7447 3292
rect 7471 3290 7527 3292
rect 7551 3290 7607 3292
rect 7631 3290 7687 3292
rect 7391 3238 7437 3290
rect 7437 3238 7447 3290
rect 7471 3238 7501 3290
rect 7501 3238 7513 3290
rect 7513 3238 7527 3290
rect 7551 3238 7565 3290
rect 7565 3238 7577 3290
rect 7577 3238 7607 3290
rect 7631 3238 7641 3290
rect 7641 3238 7687 3290
rect 7391 3236 7447 3238
rect 7471 3236 7527 3238
rect 7551 3236 7607 3238
rect 7631 3236 7687 3238
rect 7391 2202 7447 2204
rect 7471 2202 7527 2204
rect 7551 2202 7607 2204
rect 7631 2202 7687 2204
rect 7391 2150 7437 2202
rect 7437 2150 7447 2202
rect 7471 2150 7501 2202
rect 7501 2150 7513 2202
rect 7513 2150 7527 2202
rect 7551 2150 7565 2202
rect 7565 2150 7577 2202
rect 7577 2150 7607 2202
rect 7631 2150 7641 2202
rect 7641 2150 7687 2202
rect 7391 2148 7447 2150
rect 7471 2148 7527 2150
rect 7551 2148 7607 2150
rect 7631 2148 7687 2150
rect 7391 1114 7447 1116
rect 7471 1114 7527 1116
rect 7551 1114 7607 1116
rect 7631 1114 7687 1116
rect 7391 1062 7437 1114
rect 7437 1062 7447 1114
rect 7471 1062 7501 1114
rect 7501 1062 7513 1114
rect 7513 1062 7527 1114
rect 7551 1062 7565 1114
rect 7565 1062 7577 1114
rect 7577 1062 7607 1114
rect 7631 1062 7641 1114
rect 7641 1062 7687 1114
rect 7391 1060 7447 1062
rect 7471 1060 7527 1062
rect 7551 1060 7607 1062
rect 7631 1060 7687 1062
<< metal3 >>
rect 1106 4928 1422 4929
rect 1106 4864 1112 4928
rect 1176 4864 1192 4928
rect 1256 4864 1272 4928
rect 1336 4864 1352 4928
rect 1416 4864 1422 4928
rect 1106 4863 1422 4864
rect 2899 4928 3215 4929
rect 2899 4864 2905 4928
rect 2969 4864 2985 4928
rect 3049 4864 3065 4928
rect 3129 4864 3145 4928
rect 3209 4864 3215 4928
rect 2899 4863 3215 4864
rect 4692 4928 5008 4929
rect 4692 4864 4698 4928
rect 4762 4864 4778 4928
rect 4842 4864 4858 4928
rect 4922 4864 4938 4928
rect 5002 4864 5008 4928
rect 4692 4863 5008 4864
rect 6485 4928 6801 4929
rect 6485 4864 6491 4928
rect 6555 4864 6571 4928
rect 6635 4864 6651 4928
rect 6715 4864 6731 4928
rect 6795 4864 6801 4928
rect 6485 4863 6801 4864
rect 2002 4384 2318 4385
rect 2002 4320 2008 4384
rect 2072 4320 2088 4384
rect 2152 4320 2168 4384
rect 2232 4320 2248 4384
rect 2312 4320 2318 4384
rect 2002 4319 2318 4320
rect 3795 4384 4111 4385
rect 3795 4320 3801 4384
rect 3865 4320 3881 4384
rect 3945 4320 3961 4384
rect 4025 4320 4041 4384
rect 4105 4320 4111 4384
rect 3795 4319 4111 4320
rect 5588 4384 5904 4385
rect 5588 4320 5594 4384
rect 5658 4320 5674 4384
rect 5738 4320 5754 4384
rect 5818 4320 5834 4384
rect 5898 4320 5904 4384
rect 5588 4319 5904 4320
rect 7381 4384 7697 4385
rect 7381 4320 7387 4384
rect 7451 4320 7467 4384
rect 7531 4320 7547 4384
rect 7611 4320 7627 4384
rect 7691 4320 7697 4384
rect 7381 4319 7697 4320
rect 1106 3840 1422 3841
rect 1106 3776 1112 3840
rect 1176 3776 1192 3840
rect 1256 3776 1272 3840
rect 1336 3776 1352 3840
rect 1416 3776 1422 3840
rect 1106 3775 1422 3776
rect 2899 3840 3215 3841
rect 2899 3776 2905 3840
rect 2969 3776 2985 3840
rect 3049 3776 3065 3840
rect 3129 3776 3145 3840
rect 3209 3776 3215 3840
rect 2899 3775 3215 3776
rect 4692 3840 5008 3841
rect 4692 3776 4698 3840
rect 4762 3776 4778 3840
rect 4842 3776 4858 3840
rect 4922 3776 4938 3840
rect 5002 3776 5008 3840
rect 4692 3775 5008 3776
rect 6485 3840 6801 3841
rect 6485 3776 6491 3840
rect 6555 3776 6571 3840
rect 6635 3776 6651 3840
rect 6715 3776 6731 3840
rect 6795 3776 6801 3840
rect 6485 3775 6801 3776
rect 2002 3296 2318 3297
rect 2002 3232 2008 3296
rect 2072 3232 2088 3296
rect 2152 3232 2168 3296
rect 2232 3232 2248 3296
rect 2312 3232 2318 3296
rect 2002 3231 2318 3232
rect 3795 3296 4111 3297
rect 3795 3232 3801 3296
rect 3865 3232 3881 3296
rect 3945 3232 3961 3296
rect 4025 3232 4041 3296
rect 4105 3232 4111 3296
rect 3795 3231 4111 3232
rect 5588 3296 5904 3297
rect 5588 3232 5594 3296
rect 5658 3232 5674 3296
rect 5738 3232 5754 3296
rect 5818 3232 5834 3296
rect 5898 3232 5904 3296
rect 5588 3231 5904 3232
rect 7381 3296 7697 3297
rect 7381 3232 7387 3296
rect 7451 3232 7467 3296
rect 7531 3232 7547 3296
rect 7611 3232 7627 3296
rect 7691 3232 7697 3296
rect 7381 3231 7697 3232
rect 1106 2752 1422 2753
rect 1106 2688 1112 2752
rect 1176 2688 1192 2752
rect 1256 2688 1272 2752
rect 1336 2688 1352 2752
rect 1416 2688 1422 2752
rect 1106 2687 1422 2688
rect 2899 2752 3215 2753
rect 2899 2688 2905 2752
rect 2969 2688 2985 2752
rect 3049 2688 3065 2752
rect 3129 2688 3145 2752
rect 3209 2688 3215 2752
rect 2899 2687 3215 2688
rect 4692 2752 5008 2753
rect 4692 2688 4698 2752
rect 4762 2688 4778 2752
rect 4842 2688 4858 2752
rect 4922 2688 4938 2752
rect 5002 2688 5008 2752
rect 4692 2687 5008 2688
rect 6485 2752 6801 2753
rect 6485 2688 6491 2752
rect 6555 2688 6571 2752
rect 6635 2688 6651 2752
rect 6715 2688 6731 2752
rect 6795 2688 6801 2752
rect 6485 2687 6801 2688
rect 2002 2208 2318 2209
rect 2002 2144 2008 2208
rect 2072 2144 2088 2208
rect 2152 2144 2168 2208
rect 2232 2144 2248 2208
rect 2312 2144 2318 2208
rect 2002 2143 2318 2144
rect 3795 2208 4111 2209
rect 3795 2144 3801 2208
rect 3865 2144 3881 2208
rect 3945 2144 3961 2208
rect 4025 2144 4041 2208
rect 4105 2144 4111 2208
rect 3795 2143 4111 2144
rect 5588 2208 5904 2209
rect 5588 2144 5594 2208
rect 5658 2144 5674 2208
rect 5738 2144 5754 2208
rect 5818 2144 5834 2208
rect 5898 2144 5904 2208
rect 5588 2143 5904 2144
rect 7381 2208 7697 2209
rect 7381 2144 7387 2208
rect 7451 2144 7467 2208
rect 7531 2144 7547 2208
rect 7611 2144 7627 2208
rect 7691 2144 7697 2208
rect 7381 2143 7697 2144
rect 1106 1664 1422 1665
rect 1106 1600 1112 1664
rect 1176 1600 1192 1664
rect 1256 1600 1272 1664
rect 1336 1600 1352 1664
rect 1416 1600 1422 1664
rect 1106 1599 1422 1600
rect 2899 1664 3215 1665
rect 2899 1600 2905 1664
rect 2969 1600 2985 1664
rect 3049 1600 3065 1664
rect 3129 1600 3145 1664
rect 3209 1600 3215 1664
rect 2899 1599 3215 1600
rect 4692 1664 5008 1665
rect 4692 1600 4698 1664
rect 4762 1600 4778 1664
rect 4842 1600 4858 1664
rect 4922 1600 4938 1664
rect 5002 1600 5008 1664
rect 4692 1599 5008 1600
rect 6485 1664 6801 1665
rect 6485 1600 6491 1664
rect 6555 1600 6571 1664
rect 6635 1600 6651 1664
rect 6715 1600 6731 1664
rect 6795 1600 6801 1664
rect 6485 1599 6801 1600
rect 2002 1120 2318 1121
rect 2002 1056 2008 1120
rect 2072 1056 2088 1120
rect 2152 1056 2168 1120
rect 2232 1056 2248 1120
rect 2312 1056 2318 1120
rect 2002 1055 2318 1056
rect 3795 1120 4111 1121
rect 3795 1056 3801 1120
rect 3865 1056 3881 1120
rect 3945 1056 3961 1120
rect 4025 1056 4041 1120
rect 4105 1056 4111 1120
rect 3795 1055 4111 1056
rect 5588 1120 5904 1121
rect 5588 1056 5594 1120
rect 5658 1056 5674 1120
rect 5738 1056 5754 1120
rect 5818 1056 5834 1120
rect 5898 1056 5904 1120
rect 5588 1055 5904 1056
rect 7381 1120 7697 1121
rect 7381 1056 7387 1120
rect 7451 1056 7467 1120
rect 7531 1056 7547 1120
rect 7611 1056 7627 1120
rect 7691 1056 7697 1120
rect 7381 1055 7697 1056
<< via3 >>
rect 1112 4924 1176 4928
rect 1112 4868 1116 4924
rect 1116 4868 1172 4924
rect 1172 4868 1176 4924
rect 1112 4864 1176 4868
rect 1192 4924 1256 4928
rect 1192 4868 1196 4924
rect 1196 4868 1252 4924
rect 1252 4868 1256 4924
rect 1192 4864 1256 4868
rect 1272 4924 1336 4928
rect 1272 4868 1276 4924
rect 1276 4868 1332 4924
rect 1332 4868 1336 4924
rect 1272 4864 1336 4868
rect 1352 4924 1416 4928
rect 1352 4868 1356 4924
rect 1356 4868 1412 4924
rect 1412 4868 1416 4924
rect 1352 4864 1416 4868
rect 2905 4924 2969 4928
rect 2905 4868 2909 4924
rect 2909 4868 2965 4924
rect 2965 4868 2969 4924
rect 2905 4864 2969 4868
rect 2985 4924 3049 4928
rect 2985 4868 2989 4924
rect 2989 4868 3045 4924
rect 3045 4868 3049 4924
rect 2985 4864 3049 4868
rect 3065 4924 3129 4928
rect 3065 4868 3069 4924
rect 3069 4868 3125 4924
rect 3125 4868 3129 4924
rect 3065 4864 3129 4868
rect 3145 4924 3209 4928
rect 3145 4868 3149 4924
rect 3149 4868 3205 4924
rect 3205 4868 3209 4924
rect 3145 4864 3209 4868
rect 4698 4924 4762 4928
rect 4698 4868 4702 4924
rect 4702 4868 4758 4924
rect 4758 4868 4762 4924
rect 4698 4864 4762 4868
rect 4778 4924 4842 4928
rect 4778 4868 4782 4924
rect 4782 4868 4838 4924
rect 4838 4868 4842 4924
rect 4778 4864 4842 4868
rect 4858 4924 4922 4928
rect 4858 4868 4862 4924
rect 4862 4868 4918 4924
rect 4918 4868 4922 4924
rect 4858 4864 4922 4868
rect 4938 4924 5002 4928
rect 4938 4868 4942 4924
rect 4942 4868 4998 4924
rect 4998 4868 5002 4924
rect 4938 4864 5002 4868
rect 6491 4924 6555 4928
rect 6491 4868 6495 4924
rect 6495 4868 6551 4924
rect 6551 4868 6555 4924
rect 6491 4864 6555 4868
rect 6571 4924 6635 4928
rect 6571 4868 6575 4924
rect 6575 4868 6631 4924
rect 6631 4868 6635 4924
rect 6571 4864 6635 4868
rect 6651 4924 6715 4928
rect 6651 4868 6655 4924
rect 6655 4868 6711 4924
rect 6711 4868 6715 4924
rect 6651 4864 6715 4868
rect 6731 4924 6795 4928
rect 6731 4868 6735 4924
rect 6735 4868 6791 4924
rect 6791 4868 6795 4924
rect 6731 4864 6795 4868
rect 2008 4380 2072 4384
rect 2008 4324 2012 4380
rect 2012 4324 2068 4380
rect 2068 4324 2072 4380
rect 2008 4320 2072 4324
rect 2088 4380 2152 4384
rect 2088 4324 2092 4380
rect 2092 4324 2148 4380
rect 2148 4324 2152 4380
rect 2088 4320 2152 4324
rect 2168 4380 2232 4384
rect 2168 4324 2172 4380
rect 2172 4324 2228 4380
rect 2228 4324 2232 4380
rect 2168 4320 2232 4324
rect 2248 4380 2312 4384
rect 2248 4324 2252 4380
rect 2252 4324 2308 4380
rect 2308 4324 2312 4380
rect 2248 4320 2312 4324
rect 3801 4380 3865 4384
rect 3801 4324 3805 4380
rect 3805 4324 3861 4380
rect 3861 4324 3865 4380
rect 3801 4320 3865 4324
rect 3881 4380 3945 4384
rect 3881 4324 3885 4380
rect 3885 4324 3941 4380
rect 3941 4324 3945 4380
rect 3881 4320 3945 4324
rect 3961 4380 4025 4384
rect 3961 4324 3965 4380
rect 3965 4324 4021 4380
rect 4021 4324 4025 4380
rect 3961 4320 4025 4324
rect 4041 4380 4105 4384
rect 4041 4324 4045 4380
rect 4045 4324 4101 4380
rect 4101 4324 4105 4380
rect 4041 4320 4105 4324
rect 5594 4380 5658 4384
rect 5594 4324 5598 4380
rect 5598 4324 5654 4380
rect 5654 4324 5658 4380
rect 5594 4320 5658 4324
rect 5674 4380 5738 4384
rect 5674 4324 5678 4380
rect 5678 4324 5734 4380
rect 5734 4324 5738 4380
rect 5674 4320 5738 4324
rect 5754 4380 5818 4384
rect 5754 4324 5758 4380
rect 5758 4324 5814 4380
rect 5814 4324 5818 4380
rect 5754 4320 5818 4324
rect 5834 4380 5898 4384
rect 5834 4324 5838 4380
rect 5838 4324 5894 4380
rect 5894 4324 5898 4380
rect 5834 4320 5898 4324
rect 7387 4380 7451 4384
rect 7387 4324 7391 4380
rect 7391 4324 7447 4380
rect 7447 4324 7451 4380
rect 7387 4320 7451 4324
rect 7467 4380 7531 4384
rect 7467 4324 7471 4380
rect 7471 4324 7527 4380
rect 7527 4324 7531 4380
rect 7467 4320 7531 4324
rect 7547 4380 7611 4384
rect 7547 4324 7551 4380
rect 7551 4324 7607 4380
rect 7607 4324 7611 4380
rect 7547 4320 7611 4324
rect 7627 4380 7691 4384
rect 7627 4324 7631 4380
rect 7631 4324 7687 4380
rect 7687 4324 7691 4380
rect 7627 4320 7691 4324
rect 1112 3836 1176 3840
rect 1112 3780 1116 3836
rect 1116 3780 1172 3836
rect 1172 3780 1176 3836
rect 1112 3776 1176 3780
rect 1192 3836 1256 3840
rect 1192 3780 1196 3836
rect 1196 3780 1252 3836
rect 1252 3780 1256 3836
rect 1192 3776 1256 3780
rect 1272 3836 1336 3840
rect 1272 3780 1276 3836
rect 1276 3780 1332 3836
rect 1332 3780 1336 3836
rect 1272 3776 1336 3780
rect 1352 3836 1416 3840
rect 1352 3780 1356 3836
rect 1356 3780 1412 3836
rect 1412 3780 1416 3836
rect 1352 3776 1416 3780
rect 2905 3836 2969 3840
rect 2905 3780 2909 3836
rect 2909 3780 2965 3836
rect 2965 3780 2969 3836
rect 2905 3776 2969 3780
rect 2985 3836 3049 3840
rect 2985 3780 2989 3836
rect 2989 3780 3045 3836
rect 3045 3780 3049 3836
rect 2985 3776 3049 3780
rect 3065 3836 3129 3840
rect 3065 3780 3069 3836
rect 3069 3780 3125 3836
rect 3125 3780 3129 3836
rect 3065 3776 3129 3780
rect 3145 3836 3209 3840
rect 3145 3780 3149 3836
rect 3149 3780 3205 3836
rect 3205 3780 3209 3836
rect 3145 3776 3209 3780
rect 4698 3836 4762 3840
rect 4698 3780 4702 3836
rect 4702 3780 4758 3836
rect 4758 3780 4762 3836
rect 4698 3776 4762 3780
rect 4778 3836 4842 3840
rect 4778 3780 4782 3836
rect 4782 3780 4838 3836
rect 4838 3780 4842 3836
rect 4778 3776 4842 3780
rect 4858 3836 4922 3840
rect 4858 3780 4862 3836
rect 4862 3780 4918 3836
rect 4918 3780 4922 3836
rect 4858 3776 4922 3780
rect 4938 3836 5002 3840
rect 4938 3780 4942 3836
rect 4942 3780 4998 3836
rect 4998 3780 5002 3836
rect 4938 3776 5002 3780
rect 6491 3836 6555 3840
rect 6491 3780 6495 3836
rect 6495 3780 6551 3836
rect 6551 3780 6555 3836
rect 6491 3776 6555 3780
rect 6571 3836 6635 3840
rect 6571 3780 6575 3836
rect 6575 3780 6631 3836
rect 6631 3780 6635 3836
rect 6571 3776 6635 3780
rect 6651 3836 6715 3840
rect 6651 3780 6655 3836
rect 6655 3780 6711 3836
rect 6711 3780 6715 3836
rect 6651 3776 6715 3780
rect 6731 3836 6795 3840
rect 6731 3780 6735 3836
rect 6735 3780 6791 3836
rect 6791 3780 6795 3836
rect 6731 3776 6795 3780
rect 2008 3292 2072 3296
rect 2008 3236 2012 3292
rect 2012 3236 2068 3292
rect 2068 3236 2072 3292
rect 2008 3232 2072 3236
rect 2088 3292 2152 3296
rect 2088 3236 2092 3292
rect 2092 3236 2148 3292
rect 2148 3236 2152 3292
rect 2088 3232 2152 3236
rect 2168 3292 2232 3296
rect 2168 3236 2172 3292
rect 2172 3236 2228 3292
rect 2228 3236 2232 3292
rect 2168 3232 2232 3236
rect 2248 3292 2312 3296
rect 2248 3236 2252 3292
rect 2252 3236 2308 3292
rect 2308 3236 2312 3292
rect 2248 3232 2312 3236
rect 3801 3292 3865 3296
rect 3801 3236 3805 3292
rect 3805 3236 3861 3292
rect 3861 3236 3865 3292
rect 3801 3232 3865 3236
rect 3881 3292 3945 3296
rect 3881 3236 3885 3292
rect 3885 3236 3941 3292
rect 3941 3236 3945 3292
rect 3881 3232 3945 3236
rect 3961 3292 4025 3296
rect 3961 3236 3965 3292
rect 3965 3236 4021 3292
rect 4021 3236 4025 3292
rect 3961 3232 4025 3236
rect 4041 3292 4105 3296
rect 4041 3236 4045 3292
rect 4045 3236 4101 3292
rect 4101 3236 4105 3292
rect 4041 3232 4105 3236
rect 5594 3292 5658 3296
rect 5594 3236 5598 3292
rect 5598 3236 5654 3292
rect 5654 3236 5658 3292
rect 5594 3232 5658 3236
rect 5674 3292 5738 3296
rect 5674 3236 5678 3292
rect 5678 3236 5734 3292
rect 5734 3236 5738 3292
rect 5674 3232 5738 3236
rect 5754 3292 5818 3296
rect 5754 3236 5758 3292
rect 5758 3236 5814 3292
rect 5814 3236 5818 3292
rect 5754 3232 5818 3236
rect 5834 3292 5898 3296
rect 5834 3236 5838 3292
rect 5838 3236 5894 3292
rect 5894 3236 5898 3292
rect 5834 3232 5898 3236
rect 7387 3292 7451 3296
rect 7387 3236 7391 3292
rect 7391 3236 7447 3292
rect 7447 3236 7451 3292
rect 7387 3232 7451 3236
rect 7467 3292 7531 3296
rect 7467 3236 7471 3292
rect 7471 3236 7527 3292
rect 7527 3236 7531 3292
rect 7467 3232 7531 3236
rect 7547 3292 7611 3296
rect 7547 3236 7551 3292
rect 7551 3236 7607 3292
rect 7607 3236 7611 3292
rect 7547 3232 7611 3236
rect 7627 3292 7691 3296
rect 7627 3236 7631 3292
rect 7631 3236 7687 3292
rect 7687 3236 7691 3292
rect 7627 3232 7691 3236
rect 1112 2748 1176 2752
rect 1112 2692 1116 2748
rect 1116 2692 1172 2748
rect 1172 2692 1176 2748
rect 1112 2688 1176 2692
rect 1192 2748 1256 2752
rect 1192 2692 1196 2748
rect 1196 2692 1252 2748
rect 1252 2692 1256 2748
rect 1192 2688 1256 2692
rect 1272 2748 1336 2752
rect 1272 2692 1276 2748
rect 1276 2692 1332 2748
rect 1332 2692 1336 2748
rect 1272 2688 1336 2692
rect 1352 2748 1416 2752
rect 1352 2692 1356 2748
rect 1356 2692 1412 2748
rect 1412 2692 1416 2748
rect 1352 2688 1416 2692
rect 2905 2748 2969 2752
rect 2905 2692 2909 2748
rect 2909 2692 2965 2748
rect 2965 2692 2969 2748
rect 2905 2688 2969 2692
rect 2985 2748 3049 2752
rect 2985 2692 2989 2748
rect 2989 2692 3045 2748
rect 3045 2692 3049 2748
rect 2985 2688 3049 2692
rect 3065 2748 3129 2752
rect 3065 2692 3069 2748
rect 3069 2692 3125 2748
rect 3125 2692 3129 2748
rect 3065 2688 3129 2692
rect 3145 2748 3209 2752
rect 3145 2692 3149 2748
rect 3149 2692 3205 2748
rect 3205 2692 3209 2748
rect 3145 2688 3209 2692
rect 4698 2748 4762 2752
rect 4698 2692 4702 2748
rect 4702 2692 4758 2748
rect 4758 2692 4762 2748
rect 4698 2688 4762 2692
rect 4778 2748 4842 2752
rect 4778 2692 4782 2748
rect 4782 2692 4838 2748
rect 4838 2692 4842 2748
rect 4778 2688 4842 2692
rect 4858 2748 4922 2752
rect 4858 2692 4862 2748
rect 4862 2692 4918 2748
rect 4918 2692 4922 2748
rect 4858 2688 4922 2692
rect 4938 2748 5002 2752
rect 4938 2692 4942 2748
rect 4942 2692 4998 2748
rect 4998 2692 5002 2748
rect 4938 2688 5002 2692
rect 6491 2748 6555 2752
rect 6491 2692 6495 2748
rect 6495 2692 6551 2748
rect 6551 2692 6555 2748
rect 6491 2688 6555 2692
rect 6571 2748 6635 2752
rect 6571 2692 6575 2748
rect 6575 2692 6631 2748
rect 6631 2692 6635 2748
rect 6571 2688 6635 2692
rect 6651 2748 6715 2752
rect 6651 2692 6655 2748
rect 6655 2692 6711 2748
rect 6711 2692 6715 2748
rect 6651 2688 6715 2692
rect 6731 2748 6795 2752
rect 6731 2692 6735 2748
rect 6735 2692 6791 2748
rect 6791 2692 6795 2748
rect 6731 2688 6795 2692
rect 2008 2204 2072 2208
rect 2008 2148 2012 2204
rect 2012 2148 2068 2204
rect 2068 2148 2072 2204
rect 2008 2144 2072 2148
rect 2088 2204 2152 2208
rect 2088 2148 2092 2204
rect 2092 2148 2148 2204
rect 2148 2148 2152 2204
rect 2088 2144 2152 2148
rect 2168 2204 2232 2208
rect 2168 2148 2172 2204
rect 2172 2148 2228 2204
rect 2228 2148 2232 2204
rect 2168 2144 2232 2148
rect 2248 2204 2312 2208
rect 2248 2148 2252 2204
rect 2252 2148 2308 2204
rect 2308 2148 2312 2204
rect 2248 2144 2312 2148
rect 3801 2204 3865 2208
rect 3801 2148 3805 2204
rect 3805 2148 3861 2204
rect 3861 2148 3865 2204
rect 3801 2144 3865 2148
rect 3881 2204 3945 2208
rect 3881 2148 3885 2204
rect 3885 2148 3941 2204
rect 3941 2148 3945 2204
rect 3881 2144 3945 2148
rect 3961 2204 4025 2208
rect 3961 2148 3965 2204
rect 3965 2148 4021 2204
rect 4021 2148 4025 2204
rect 3961 2144 4025 2148
rect 4041 2204 4105 2208
rect 4041 2148 4045 2204
rect 4045 2148 4101 2204
rect 4101 2148 4105 2204
rect 4041 2144 4105 2148
rect 5594 2204 5658 2208
rect 5594 2148 5598 2204
rect 5598 2148 5654 2204
rect 5654 2148 5658 2204
rect 5594 2144 5658 2148
rect 5674 2204 5738 2208
rect 5674 2148 5678 2204
rect 5678 2148 5734 2204
rect 5734 2148 5738 2204
rect 5674 2144 5738 2148
rect 5754 2204 5818 2208
rect 5754 2148 5758 2204
rect 5758 2148 5814 2204
rect 5814 2148 5818 2204
rect 5754 2144 5818 2148
rect 5834 2204 5898 2208
rect 5834 2148 5838 2204
rect 5838 2148 5894 2204
rect 5894 2148 5898 2204
rect 5834 2144 5898 2148
rect 7387 2204 7451 2208
rect 7387 2148 7391 2204
rect 7391 2148 7447 2204
rect 7447 2148 7451 2204
rect 7387 2144 7451 2148
rect 7467 2204 7531 2208
rect 7467 2148 7471 2204
rect 7471 2148 7527 2204
rect 7527 2148 7531 2204
rect 7467 2144 7531 2148
rect 7547 2204 7611 2208
rect 7547 2148 7551 2204
rect 7551 2148 7607 2204
rect 7607 2148 7611 2204
rect 7547 2144 7611 2148
rect 7627 2204 7691 2208
rect 7627 2148 7631 2204
rect 7631 2148 7687 2204
rect 7687 2148 7691 2204
rect 7627 2144 7691 2148
rect 1112 1660 1176 1664
rect 1112 1604 1116 1660
rect 1116 1604 1172 1660
rect 1172 1604 1176 1660
rect 1112 1600 1176 1604
rect 1192 1660 1256 1664
rect 1192 1604 1196 1660
rect 1196 1604 1252 1660
rect 1252 1604 1256 1660
rect 1192 1600 1256 1604
rect 1272 1660 1336 1664
rect 1272 1604 1276 1660
rect 1276 1604 1332 1660
rect 1332 1604 1336 1660
rect 1272 1600 1336 1604
rect 1352 1660 1416 1664
rect 1352 1604 1356 1660
rect 1356 1604 1412 1660
rect 1412 1604 1416 1660
rect 1352 1600 1416 1604
rect 2905 1660 2969 1664
rect 2905 1604 2909 1660
rect 2909 1604 2965 1660
rect 2965 1604 2969 1660
rect 2905 1600 2969 1604
rect 2985 1660 3049 1664
rect 2985 1604 2989 1660
rect 2989 1604 3045 1660
rect 3045 1604 3049 1660
rect 2985 1600 3049 1604
rect 3065 1660 3129 1664
rect 3065 1604 3069 1660
rect 3069 1604 3125 1660
rect 3125 1604 3129 1660
rect 3065 1600 3129 1604
rect 3145 1660 3209 1664
rect 3145 1604 3149 1660
rect 3149 1604 3205 1660
rect 3205 1604 3209 1660
rect 3145 1600 3209 1604
rect 4698 1660 4762 1664
rect 4698 1604 4702 1660
rect 4702 1604 4758 1660
rect 4758 1604 4762 1660
rect 4698 1600 4762 1604
rect 4778 1660 4842 1664
rect 4778 1604 4782 1660
rect 4782 1604 4838 1660
rect 4838 1604 4842 1660
rect 4778 1600 4842 1604
rect 4858 1660 4922 1664
rect 4858 1604 4862 1660
rect 4862 1604 4918 1660
rect 4918 1604 4922 1660
rect 4858 1600 4922 1604
rect 4938 1660 5002 1664
rect 4938 1604 4942 1660
rect 4942 1604 4998 1660
rect 4998 1604 5002 1660
rect 4938 1600 5002 1604
rect 6491 1660 6555 1664
rect 6491 1604 6495 1660
rect 6495 1604 6551 1660
rect 6551 1604 6555 1660
rect 6491 1600 6555 1604
rect 6571 1660 6635 1664
rect 6571 1604 6575 1660
rect 6575 1604 6631 1660
rect 6631 1604 6635 1660
rect 6571 1600 6635 1604
rect 6651 1660 6715 1664
rect 6651 1604 6655 1660
rect 6655 1604 6711 1660
rect 6711 1604 6715 1660
rect 6651 1600 6715 1604
rect 6731 1660 6795 1664
rect 6731 1604 6735 1660
rect 6735 1604 6791 1660
rect 6791 1604 6795 1660
rect 6731 1600 6795 1604
rect 2008 1116 2072 1120
rect 2008 1060 2012 1116
rect 2012 1060 2068 1116
rect 2068 1060 2072 1116
rect 2008 1056 2072 1060
rect 2088 1116 2152 1120
rect 2088 1060 2092 1116
rect 2092 1060 2148 1116
rect 2148 1060 2152 1116
rect 2088 1056 2152 1060
rect 2168 1116 2232 1120
rect 2168 1060 2172 1116
rect 2172 1060 2228 1116
rect 2228 1060 2232 1116
rect 2168 1056 2232 1060
rect 2248 1116 2312 1120
rect 2248 1060 2252 1116
rect 2252 1060 2308 1116
rect 2308 1060 2312 1116
rect 2248 1056 2312 1060
rect 3801 1116 3865 1120
rect 3801 1060 3805 1116
rect 3805 1060 3861 1116
rect 3861 1060 3865 1116
rect 3801 1056 3865 1060
rect 3881 1116 3945 1120
rect 3881 1060 3885 1116
rect 3885 1060 3941 1116
rect 3941 1060 3945 1116
rect 3881 1056 3945 1060
rect 3961 1116 4025 1120
rect 3961 1060 3965 1116
rect 3965 1060 4021 1116
rect 4021 1060 4025 1116
rect 3961 1056 4025 1060
rect 4041 1116 4105 1120
rect 4041 1060 4045 1116
rect 4045 1060 4101 1116
rect 4101 1060 4105 1116
rect 4041 1056 4105 1060
rect 5594 1116 5658 1120
rect 5594 1060 5598 1116
rect 5598 1060 5654 1116
rect 5654 1060 5658 1116
rect 5594 1056 5658 1060
rect 5674 1116 5738 1120
rect 5674 1060 5678 1116
rect 5678 1060 5734 1116
rect 5734 1060 5738 1116
rect 5674 1056 5738 1060
rect 5754 1116 5818 1120
rect 5754 1060 5758 1116
rect 5758 1060 5814 1116
rect 5814 1060 5818 1116
rect 5754 1056 5818 1060
rect 5834 1116 5898 1120
rect 5834 1060 5838 1116
rect 5838 1060 5894 1116
rect 5894 1060 5898 1116
rect 5834 1056 5898 1060
rect 7387 1116 7451 1120
rect 7387 1060 7391 1116
rect 7391 1060 7447 1116
rect 7447 1060 7451 1116
rect 7387 1056 7451 1060
rect 7467 1116 7531 1120
rect 7467 1060 7471 1116
rect 7471 1060 7527 1116
rect 7527 1060 7531 1116
rect 7467 1056 7531 1060
rect 7547 1116 7611 1120
rect 7547 1060 7551 1116
rect 7551 1060 7607 1116
rect 7607 1060 7611 1116
rect 7547 1056 7611 1060
rect 7627 1116 7691 1120
rect 7627 1060 7631 1116
rect 7631 1060 7687 1116
rect 7687 1060 7691 1116
rect 7627 1056 7691 1060
<< metal4 >>
rect 1104 4928 1424 4944
rect 1104 4864 1112 4928
rect 1176 4864 1192 4928
rect 1256 4864 1272 4928
rect 1336 4864 1352 4928
rect 1416 4864 1424 4928
rect 1104 3840 1424 4864
rect 1104 3776 1112 3840
rect 1176 3776 1192 3840
rect 1256 3776 1272 3840
rect 1336 3776 1352 3840
rect 1416 3776 1424 3840
rect 1104 2752 1424 3776
rect 1104 2688 1112 2752
rect 1176 2688 1192 2752
rect 1256 2688 1272 2752
rect 1336 2688 1352 2752
rect 1416 2688 1424 2752
rect 1104 1664 1424 2688
rect 1104 1600 1112 1664
rect 1176 1600 1192 1664
rect 1256 1600 1272 1664
rect 1336 1600 1352 1664
rect 1416 1600 1424 1664
rect 1104 1040 1424 1600
rect 2000 4384 2320 4944
rect 2000 4320 2008 4384
rect 2072 4320 2088 4384
rect 2152 4320 2168 4384
rect 2232 4320 2248 4384
rect 2312 4320 2320 4384
rect 2000 3296 2320 4320
rect 2000 3232 2008 3296
rect 2072 3232 2088 3296
rect 2152 3232 2168 3296
rect 2232 3232 2248 3296
rect 2312 3232 2320 3296
rect 2000 2208 2320 3232
rect 2000 2144 2008 2208
rect 2072 2144 2088 2208
rect 2152 2144 2168 2208
rect 2232 2144 2248 2208
rect 2312 2144 2320 2208
rect 2000 1120 2320 2144
rect 2000 1056 2008 1120
rect 2072 1056 2088 1120
rect 2152 1056 2168 1120
rect 2232 1056 2248 1120
rect 2312 1056 2320 1120
rect 2000 1040 2320 1056
rect 2897 4928 3217 4944
rect 2897 4864 2905 4928
rect 2969 4864 2985 4928
rect 3049 4864 3065 4928
rect 3129 4864 3145 4928
rect 3209 4864 3217 4928
rect 2897 3840 3217 4864
rect 2897 3776 2905 3840
rect 2969 3776 2985 3840
rect 3049 3776 3065 3840
rect 3129 3776 3145 3840
rect 3209 3776 3217 3840
rect 2897 2752 3217 3776
rect 2897 2688 2905 2752
rect 2969 2688 2985 2752
rect 3049 2688 3065 2752
rect 3129 2688 3145 2752
rect 3209 2688 3217 2752
rect 2897 1664 3217 2688
rect 2897 1600 2905 1664
rect 2969 1600 2985 1664
rect 3049 1600 3065 1664
rect 3129 1600 3145 1664
rect 3209 1600 3217 1664
rect 2897 1040 3217 1600
rect 3793 4384 4113 4944
rect 3793 4320 3801 4384
rect 3865 4320 3881 4384
rect 3945 4320 3961 4384
rect 4025 4320 4041 4384
rect 4105 4320 4113 4384
rect 3793 3296 4113 4320
rect 3793 3232 3801 3296
rect 3865 3232 3881 3296
rect 3945 3232 3961 3296
rect 4025 3232 4041 3296
rect 4105 3232 4113 3296
rect 3793 2208 4113 3232
rect 3793 2144 3801 2208
rect 3865 2144 3881 2208
rect 3945 2144 3961 2208
rect 4025 2144 4041 2208
rect 4105 2144 4113 2208
rect 3793 1120 4113 2144
rect 3793 1056 3801 1120
rect 3865 1056 3881 1120
rect 3945 1056 3961 1120
rect 4025 1056 4041 1120
rect 4105 1056 4113 1120
rect 3793 1040 4113 1056
rect 4690 4928 5010 4944
rect 4690 4864 4698 4928
rect 4762 4864 4778 4928
rect 4842 4864 4858 4928
rect 4922 4864 4938 4928
rect 5002 4864 5010 4928
rect 4690 3840 5010 4864
rect 4690 3776 4698 3840
rect 4762 3776 4778 3840
rect 4842 3776 4858 3840
rect 4922 3776 4938 3840
rect 5002 3776 5010 3840
rect 4690 2752 5010 3776
rect 4690 2688 4698 2752
rect 4762 2688 4778 2752
rect 4842 2688 4858 2752
rect 4922 2688 4938 2752
rect 5002 2688 5010 2752
rect 4690 1664 5010 2688
rect 4690 1600 4698 1664
rect 4762 1600 4778 1664
rect 4842 1600 4858 1664
rect 4922 1600 4938 1664
rect 5002 1600 5010 1664
rect 4690 1040 5010 1600
rect 5586 4384 5906 4944
rect 5586 4320 5594 4384
rect 5658 4320 5674 4384
rect 5738 4320 5754 4384
rect 5818 4320 5834 4384
rect 5898 4320 5906 4384
rect 5586 3296 5906 4320
rect 5586 3232 5594 3296
rect 5658 3232 5674 3296
rect 5738 3232 5754 3296
rect 5818 3232 5834 3296
rect 5898 3232 5906 3296
rect 5586 2208 5906 3232
rect 5586 2144 5594 2208
rect 5658 2144 5674 2208
rect 5738 2144 5754 2208
rect 5818 2144 5834 2208
rect 5898 2144 5906 2208
rect 5586 1120 5906 2144
rect 5586 1056 5594 1120
rect 5658 1056 5674 1120
rect 5738 1056 5754 1120
rect 5818 1056 5834 1120
rect 5898 1056 5906 1120
rect 5586 1040 5906 1056
rect 6483 4928 6803 4944
rect 6483 4864 6491 4928
rect 6555 4864 6571 4928
rect 6635 4864 6651 4928
rect 6715 4864 6731 4928
rect 6795 4864 6803 4928
rect 6483 3840 6803 4864
rect 6483 3776 6491 3840
rect 6555 3776 6571 3840
rect 6635 3776 6651 3840
rect 6715 3776 6731 3840
rect 6795 3776 6803 3840
rect 6483 2752 6803 3776
rect 6483 2688 6491 2752
rect 6555 2688 6571 2752
rect 6635 2688 6651 2752
rect 6715 2688 6731 2752
rect 6795 2688 6803 2752
rect 6483 1664 6803 2688
rect 6483 1600 6491 1664
rect 6555 1600 6571 1664
rect 6635 1600 6651 1664
rect 6715 1600 6731 1664
rect 6795 1600 6803 1664
rect 6483 1040 6803 1600
rect 7379 4384 7699 4944
rect 7379 4320 7387 4384
rect 7451 4320 7467 4384
rect 7531 4320 7547 4384
rect 7611 4320 7627 4384
rect 7691 4320 7699 4384
rect 7379 3296 7699 4320
rect 7379 3232 7387 3296
rect 7451 3232 7467 3296
rect 7531 3232 7547 3296
rect 7611 3232 7627 3296
rect 7691 3232 7699 3296
rect 7379 2208 7699 3232
rect 7379 2144 7387 2208
rect 7451 2144 7467 2208
rect 7531 2144 7547 2208
rect 7611 2144 7627 2208
rect 7691 2144 7699 2208
rect 7379 1120 7699 2144
rect 7379 1056 7387 1120
rect 7451 1056 7467 1120
rect 7531 1056 7547 1120
rect 7611 1056 7627 1120
rect 7691 1056 7699 1120
rect 7379 1040 7699 1056
use sky130_fd_sc_hd__buf_8  BUF\[0\] OL_LATEST/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 1104 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  BUF\[1\]
timestamp 1665323087
transform 1 0 552 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  BUF\[2\]
timestamp 1665323087
transform 1 0 1104 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  BUF\[3\]
timestamp 1665323087
transform 1 0 1288 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  BUF\[4\]
timestamp 1665323087
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  BUF\[5\]
timestamp 1665323087
transform 1 0 2024 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  BUF\[6\]
timestamp 1665323087
transform -1 0 2392 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  BUF\[7\]
timestamp 1665323087
transform 1 0 3220 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  BUF\[8\]
timestamp 1665323087
transform -1 0 3864 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  BUF\[9\]
timestamp 1665323087
transform 1 0 3404 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  BUF\[10\]
timestamp 1665323087
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  BUF\[11\]
timestamp 1665323087
transform 1 0 4140 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  BUF\[12\]
timestamp 1665323087
transform -1 0 5336 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  BUF\[13\]
timestamp 1665323087
transform 1 0 5796 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  BUF\[14\]
timestamp 1665323087
transform 1 0 5796 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  BUF\[15\]
timestamp 1665323087
transform -1 0 5336 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  BUF\[16\]
timestamp 1665323087
transform -1 0 6808 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  BUF\[17\]
timestamp 1665323087
transform -1 0 6900 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  BUF\[18\]
timestamp 1665323087
transform -1 0 6900 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  BUF\[19\]
timestamp 1665323087
transform -1 0 6900 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0 OL_LATEST/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 368 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8 OL_LATEST/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 1104 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22 OL_LATEST/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 2392 0 1 1088
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29 OL_LATEST/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 3036 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1665323087
transform 1 0 4140 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 OL_LATEST/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 5244 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1665323087
transform 1 0 5612 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71
timestamp 1665323087
transform 1 0 6900 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77 OL_LATEST/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 7452 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_0
timestamp 1665323087
transform 1 0 368 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_14 OL_LATEST/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 1656 0 -1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_30
timestamp 1665323087
transform 1 0 3128 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1665323087
transform 1 0 5336 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1665323087
transform 1 0 5612 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_71
timestamp 1665323087
transform 1 0 6900 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_77
timestamp 1665323087
transform 1 0 7452 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_0
timestamp 1665323087
transform 1 0 368 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20
timestamp 1665323087
transform 1 0 2208 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1665323087
transform 1 0 3036 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1665323087
transform 1 0 4140 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_53
timestamp 1665323087
transform 1 0 5244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_57
timestamp 1665323087
transform 1 0 5612 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_70
timestamp 1665323087
transform 1 0 6808 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_0
timestamp 1665323087
transform 1 0 368 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_20
timestamp 1665323087
transform 1 0 2208 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_32
timestamp 1665323087
transform 1 0 3312 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_40
timestamp 1665323087
transform 1 0 4048 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_53
timestamp 1665323087
transform 1 0 5244 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1665323087
transform 1 0 5612 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_71
timestamp 1665323087
transform 1 0 6900 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_77
timestamp 1665323087
transform 1 0 7452 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_0
timestamp 1665323087
transform 1 0 368 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_8
timestamp 1665323087
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_23
timestamp 1665323087
transform 1 0 2484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1665323087
transform 1 0 2852 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_29
timestamp 1665323087
transform 1 0 3036 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_45
timestamp 1665323087
transform 1 0 4508 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_61
timestamp 1665323087
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_73
timestamp 1665323087
transform 1 0 7084 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_77
timestamp 1665323087
transform 1 0 7452 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_0
timestamp 1665323087
transform 1 0 368 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_8
timestamp 1665323087
transform 1 0 1104 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_22
timestamp 1665323087
transform 1 0 2392 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_38
timestamp 1665323087
transform 1 0 3864 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1665323087
transform 1 0 5336 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1665323087
transform 1 0 5612 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_71
timestamp 1665323087
transform 1 0 6900 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_77
timestamp 1665323087
transform 1 0 7452 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_0
timestamp 1665323087
transform 1 0 368 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_12
timestamp 1665323087
transform 1 0 1472 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1665323087
transform 1 0 2576 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1665323087
transform 1 0 3036 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_43
timestamp 1665323087
transform 1 0 4324 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_55
timestamp 1665323087
transform 1 0 5428 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_57
timestamp 1665323087
transform 1 0 5612 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_71
timestamp 1665323087
transform 1 0 6900 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_77
timestamp 1665323087
transform 1 0 7452 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_0 OL_LATEST/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 2944 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1
timestamp 1665323087
transform 1 0 5520 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2
timestamp 1665323087
transform 1 0 5520 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3
timestamp 1665323087
transform 1 0 2944 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_4
timestamp 1665323087
transform 1 0 5520 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_5
timestamp 1665323087
transform 1 0 2944 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_6
timestamp 1665323087
transform 1 0 5520 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_7
timestamp 1665323087
transform 1 0 2944 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_8
timestamp 1665323087
transform 1 0 5520 0 1 4352
box -38 -48 130 592
<< labels >>
flabel metal4 s 2000 1040 2320 4944 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 3793 1040 4113 4944 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 5586 1040 5906 4944 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 7379 1040 7699 4944 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 1104 1040 1424 4944 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 2897 1040 3217 4944 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 4690 1040 5010 4944 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 6483 1040 6803 4944 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 478 0 534 800 0 FreeSans 224 90 0 0 in[0]
port 2 nsew signal input
flabel metal2 s 4158 0 4214 800 0 FreeSans 224 90 0 0 in[10]
port 3 nsew signal input
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 in[11]
port 4 nsew signal input
flabel metal2 s 4894 0 4950 800 0 FreeSans 224 90 0 0 in[12]
port 5 nsew signal input
flabel metal2 s 5262 0 5318 800 0 FreeSans 224 90 0 0 in[13]
port 6 nsew signal input
flabel metal2 s 5630 0 5686 800 0 FreeSans 224 90 0 0 in[14]
port 7 nsew signal input
flabel metal2 s 5998 0 6054 800 0 FreeSans 224 90 0 0 in[15]
port 8 nsew signal input
flabel metal2 s 6366 0 6422 800 0 FreeSans 224 90 0 0 in[16]
port 9 nsew signal input
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 in[17]
port 10 nsew signal input
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 in[18]
port 11 nsew signal input
flabel metal2 s 7470 0 7526 800 0 FreeSans 224 90 0 0 in[19]
port 12 nsew signal input
flabel metal2 s 846 0 902 800 0 FreeSans 224 90 0 0 in[1]
port 13 nsew signal input
flabel metal2 s 1214 0 1270 800 0 FreeSans 224 90 0 0 in[2]
port 14 nsew signal input
flabel metal2 s 1582 0 1638 800 0 FreeSans 224 90 0 0 in[3]
port 15 nsew signal input
flabel metal2 s 1950 0 2006 800 0 FreeSans 224 90 0 0 in[4]
port 16 nsew signal input
flabel metal2 s 2318 0 2374 800 0 FreeSans 224 90 0 0 in[5]
port 17 nsew signal input
flabel metal2 s 2686 0 2742 800 0 FreeSans 224 90 0 0 in[6]
port 18 nsew signal input
flabel metal2 s 3054 0 3110 800 0 FreeSans 224 90 0 0 in[7]
port 19 nsew signal input
flabel metal2 s 3422 0 3478 800 0 FreeSans 224 90 0 0 in[8]
port 20 nsew signal input
flabel metal2 s 3790 0 3846 800 0 FreeSans 224 90 0 0 in[9]
port 21 nsew signal input
flabel metal2 s 478 5200 534 6000 0 FreeSans 224 90 0 0 out[0]
port 22 nsew signal tristate
flabel metal2 s 4158 5200 4214 6000 0 FreeSans 224 90 0 0 out[10]
port 23 nsew signal tristate
flabel metal2 s 4526 5200 4582 6000 0 FreeSans 224 90 0 0 out[11]
port 24 nsew signal tristate
flabel metal2 s 4894 5200 4950 6000 0 FreeSans 224 90 0 0 out[12]
port 25 nsew signal tristate
flabel metal2 s 5262 5200 5318 6000 0 FreeSans 224 90 0 0 out[13]
port 26 nsew signal tristate
flabel metal2 s 5630 5200 5686 6000 0 FreeSans 224 90 0 0 out[14]
port 27 nsew signal tristate
flabel metal2 s 5998 5200 6054 6000 0 FreeSans 224 90 0 0 out[15]
port 28 nsew signal tristate
flabel metal2 s 6366 5200 6422 6000 0 FreeSans 224 90 0 0 out[16]
port 29 nsew signal tristate
flabel metal2 s 6734 5200 6790 6000 0 FreeSans 224 90 0 0 out[17]
port 30 nsew signal tristate
flabel metal2 s 7102 5200 7158 6000 0 FreeSans 224 90 0 0 out[18]
port 31 nsew signal tristate
flabel metal2 s 7470 5200 7526 6000 0 FreeSans 224 90 0 0 out[19]
port 32 nsew signal tristate
flabel metal2 s 846 5200 902 6000 0 FreeSans 224 90 0 0 out[1]
port 33 nsew signal tristate
flabel metal2 s 1214 5200 1270 6000 0 FreeSans 224 90 0 0 out[2]
port 34 nsew signal tristate
flabel metal2 s 1582 5200 1638 6000 0 FreeSans 224 90 0 0 out[3]
port 35 nsew signal tristate
flabel metal2 s 1950 5200 2006 6000 0 FreeSans 224 90 0 0 out[4]
port 36 nsew signal tristate
flabel metal2 s 2318 5200 2374 6000 0 FreeSans 224 90 0 0 out[5]
port 37 nsew signal tristate
flabel metal2 s 2686 5200 2742 6000 0 FreeSans 224 90 0 0 out[6]
port 38 nsew signal tristate
flabel metal2 s 3054 5200 3110 6000 0 FreeSans 224 90 0 0 out[7]
port 39 nsew signal tristate
flabel metal2 s 3422 5200 3478 6000 0 FreeSans 224 90 0 0 out[8]
port 40 nsew signal tristate
flabel metal2 s 3790 5200 3846 6000 0 FreeSans 224 90 0 0 out[9]
port 41 nsew signal tristate
rlabel via1 4033 4352 4033 4352 0 VGND
rlabel metal1 3956 4896 3956 4896 0 VPWR
rlabel metal2 506 1588 506 1588 0 in[0]
rlabel metal2 4186 2132 4186 2132 0 in[10]
rlabel metal1 4416 3026 4416 3026 0 in[11]
rlabel metal2 4922 1095 4922 1095 0 in[12]
rlabel metal2 5290 2438 5290 2438 0 in[13]
rlabel metal2 5658 823 5658 823 0 in[14]
rlabel metal1 5290 1904 5290 1904 0 in[15]
rlabel metal2 6394 1588 6394 1588 0 in[16]
rlabel metal2 6762 1044 6762 1044 0 in[17]
rlabel metal1 6992 3026 6992 3026 0 in[18]
rlabel metal1 7084 4590 7084 4590 0 in[19]
rlabel metal1 828 1938 828 1938 0 in[1]
rlabel metal2 1242 1095 1242 1095 0 in[2]
rlabel metal1 1564 1326 1564 1326 0 in[3]
rlabel metal1 1610 3468 1610 3468 0 in[4]
rlabel metal1 2346 1938 2346 1938 0 in[5]
rlabel metal1 2530 4114 2530 4114 0 in[6]
rlabel metal2 3082 1095 3082 1095 0 in[7]
rlabel metal2 3450 2438 3450 2438 0 in[8]
rlabel metal1 3680 3502 3680 3502 0 in[9]
rlabel metal1 1518 2516 1518 2516 0 out[0]
rlabel metal1 5290 3604 5290 3604 0 out[10]
rlabel metal2 4554 4090 4554 4090 0 out[11]
rlabel metal2 4646 4641 4646 4641 0 out[12]
rlabel metal1 5888 4046 5888 4046 0 out[13]
rlabel metal2 6210 3213 6210 3213 0 out[14]
rlabel metal1 4922 1836 4922 1836 0 out[15]
rlabel metal1 6302 2516 6302 2516 0 out[16]
rlabel metal1 6440 1258 6440 1258 0 out[17]
rlabel metal1 6762 2958 6762 2958 0 out[18]
rlabel metal1 6992 4658 6992 4658 0 out[19]
rlabel metal2 966 2737 966 2737 0 out[1]
rlabel metal1 1472 2958 1472 2958 0 out[2]
rlabel metal1 1932 1326 1932 1326 0 out[3]
rlabel metal2 1886 4063 1886 4063 0 out[4]
rlabel metal2 2530 3213 2530 3213 0 out[5]
rlabel metal1 2300 4046 2300 4046 0 out[6]
rlabel metal1 3634 4692 3634 4692 0 out[7]
rlabel metal2 3358 4369 3358 4369 0 out[8]
rlabel metal1 3818 3604 3818 3604 0 out[9]
<< properties >>
string FIXED_BBOX 0 0 8000 6000
<< end >>
