magic
tech sky130A
magscale 1 2
timestamp 1636370565
<< obsli1 >>
rect 1104 493 14139 13617
<< obsm1 >>
rect 934 484 14246 13648
<< metal2 >>
rect 754 14200 810 15000
rect 2226 14200 2282 15000
rect 3698 14200 3754 15000
rect 5170 14200 5226 15000
rect 6734 14200 6790 15000
rect 8206 14200 8262 15000
rect 9678 14200 9734 15000
rect 11242 14200 11298 15000
rect 12714 14200 12770 15000
rect 14186 14200 14242 15000
rect 938 0 994 800
rect 2778 0 2834 800
rect 4618 0 4674 800
rect 6550 0 6606 800
rect 8390 0 8446 800
rect 10230 0 10286 800
rect 12162 0 12218 800
rect 14002 0 14058 800
<< obsm2 >>
rect 866 14144 2170 14521
rect 2338 14144 3642 14521
rect 3810 14144 5114 14521
rect 5282 14144 6678 14521
rect 6846 14144 8150 14521
rect 8318 14144 9622 14521
rect 9790 14144 11186 14521
rect 11354 14144 12658 14521
rect 12826 14144 14130 14521
rect 754 856 14240 14144
rect 754 439 882 856
rect 1050 439 2722 856
rect 2890 439 4562 856
rect 4730 439 6494 856
rect 6662 439 8334 856
rect 8502 439 10174 856
rect 10342 439 12106 856
rect 12274 439 13946 856
rect 14114 439 14240 856
<< metal3 >>
rect 14200 14424 15000 14544
rect 14200 13608 15000 13728
rect 14200 12656 15000 12776
rect 14200 11840 15000 11960
rect 0 11160 800 11280
rect 14200 10888 15000 11008
rect 14200 10072 15000 10192
rect 14200 9120 15000 9240
rect 14200 8304 15000 8424
rect 14200 7352 15000 7472
rect 14200 6536 15000 6656
rect 14200 5584 15000 5704
rect 14200 4768 15000 4888
rect 0 3680 800 3800
rect 14200 3816 15000 3936
rect 14200 3000 15000 3120
rect 14200 2048 15000 2168
rect 14200 1232 15000 1352
rect 14200 416 15000 536
<< obsm3 >>
rect 749 14344 14120 14517
rect 749 13808 14200 14344
rect 749 13528 14120 13808
rect 749 12856 14200 13528
rect 749 12576 14120 12856
rect 749 12040 14200 12576
rect 749 11760 14120 12040
rect 749 11360 14200 11760
rect 880 11088 14200 11360
rect 880 11080 14120 11088
rect 749 10808 14120 11080
rect 749 10272 14200 10808
rect 749 9992 14120 10272
rect 749 9320 14200 9992
rect 749 9040 14120 9320
rect 749 8504 14200 9040
rect 749 8224 14120 8504
rect 749 7552 14200 8224
rect 749 7272 14120 7552
rect 749 6736 14200 7272
rect 749 6456 14120 6736
rect 749 5784 14200 6456
rect 749 5504 14120 5784
rect 749 4968 14200 5504
rect 749 4688 14120 4968
rect 749 4016 14200 4688
rect 749 3880 14120 4016
rect 880 3736 14120 3880
rect 880 3600 14200 3736
rect 749 3200 14200 3600
rect 749 2920 14120 3200
rect 749 2248 14200 2920
rect 749 1968 14120 2248
rect 749 1432 14200 1968
rect 749 1152 14120 1432
rect 749 616 14200 1152
rect 749 443 14120 616
<< metal4 >>
rect 4208 1040 4528 13648
rect 8208 1040 8528 13648
rect 12208 1040 12528 13648
<< obsm4 >>
rect 9075 4251 9877 6085
<< metal5 >>
rect 1104 12210 13892 12530
rect 1104 8210 13892 8530
rect 1104 4210 13892 4530
<< labels >>
rlabel metal5 s 1104 8210 13892 8530 6 VGND
port 1 nsew ground input
rlabel metal4 s 8208 1040 8528 13648 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 4210 13892 4530 6 VPWR
port 2 nsew power input
rlabel metal5 s 1104 12210 13892 12530 6 VPWR
port 2 nsew power input
rlabel metal4 s 4208 1040 4528 13648 6 VPWR
port 2 nsew power input
rlabel metal4 s 12208 1040 12528 13648 6 VPWR
port 2 nsew power input
rlabel metal3 s 0 3680 800 3800 6 clockp[0]
port 3 nsew signal output
rlabel metal3 s 0 11160 800 11280 6 clockp[1]
port 4 nsew signal output
rlabel metal3 s 14200 14424 15000 14544 6 dco
port 5 nsew signal input
rlabel metal3 s 14200 10072 15000 10192 6 div[0]
port 6 nsew signal input
rlabel metal3 s 14200 10888 15000 11008 6 div[1]
port 7 nsew signal input
rlabel metal3 s 14200 11840 15000 11960 6 div[2]
port 8 nsew signal input
rlabel metal3 s 14200 12656 15000 12776 6 div[3]
port 9 nsew signal input
rlabel metal3 s 14200 13608 15000 13728 6 div[4]
port 10 nsew signal input
rlabel metal3 s 14200 9120 15000 9240 6 enable
port 11 nsew signal input
rlabel metal2 s 754 14200 810 15000 6 ext_trim[0]
port 12 nsew signal input
rlabel metal3 s 14200 416 15000 536 6 ext_trim[10]
port 13 nsew signal input
rlabel metal3 s 14200 1232 15000 1352 6 ext_trim[11]
port 14 nsew signal input
rlabel metal3 s 14200 2048 15000 2168 6 ext_trim[12]
port 15 nsew signal input
rlabel metal3 s 14200 3000 15000 3120 6 ext_trim[13]
port 16 nsew signal input
rlabel metal3 s 14200 3816 15000 3936 6 ext_trim[14]
port 17 nsew signal input
rlabel metal3 s 14200 4768 15000 4888 6 ext_trim[15]
port 18 nsew signal input
rlabel metal3 s 14200 5584 15000 5704 6 ext_trim[16]
port 19 nsew signal input
rlabel metal3 s 14200 6536 15000 6656 6 ext_trim[17]
port 20 nsew signal input
rlabel metal3 s 14200 7352 15000 7472 6 ext_trim[18]
port 21 nsew signal input
rlabel metal3 s 14200 8304 15000 8424 6 ext_trim[19]
port 22 nsew signal input
rlabel metal2 s 2226 14200 2282 15000 6 ext_trim[1]
port 23 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 ext_trim[20]
port 24 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 ext_trim[21]
port 25 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 ext_trim[22]
port 26 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 ext_trim[23]
port 27 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 ext_trim[24]
port 28 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 ext_trim[25]
port 29 nsew signal input
rlabel metal2 s 3698 14200 3754 15000 6 ext_trim[2]
port 30 nsew signal input
rlabel metal2 s 5170 14200 5226 15000 6 ext_trim[3]
port 31 nsew signal input
rlabel metal2 s 6734 14200 6790 15000 6 ext_trim[4]
port 32 nsew signal input
rlabel metal2 s 8206 14200 8262 15000 6 ext_trim[5]
port 33 nsew signal input
rlabel metal2 s 9678 14200 9734 15000 6 ext_trim[6]
port 34 nsew signal input
rlabel metal2 s 11242 14200 11298 15000 6 ext_trim[7]
port 35 nsew signal input
rlabel metal2 s 12714 14200 12770 15000 6 ext_trim[8]
port 36 nsew signal input
rlabel metal2 s 14186 14200 14242 15000 6 ext_trim[9]
port 37 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 osc
port 38 nsew signal input
rlabel metal2 s 938 0 994 800 6 resetb
port 39 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 15000 15000
string LEFview TRUE
string GDS_FILE /project/openlane/digital_pll/runs/digital_pll/results/magic/digital_pll.gds
string GDS_END 1101688
string GDS_START 333802
<< end >>

